module picorv32(clk, resetn, trap, mem_valid, mem_instr, mem_ready, mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, irq, eoi, trace_valid, trace_data);
wire _00000_;
wire _00001_;
wire _00002_;
wire _00003_;
wire _00004_;
wire [31:0] _00005_;
wire [4:0] _00006_;
wire [4:0] _00007_;
wire [4:0] _00008_;
wire _00009_;
wire _00010_;
wire _00011_;
wire _00012_;
wire _00013_;
wire _00014_;
wire _00015_;
wire _00016_;
wire _00017_;
wire _00018_;
wire _00019_;
wire _00020_;
wire _00021_;
wire _00022_;
wire _00023_;
wire _00024_;
wire _00025_;
wire _00026_;
wire _00027_;
wire _00028_;
wire _00029_;
wire _00030_;
wire _00031_;
wire _00032_;
wire _00033_;
wire _00034_;
wire _00035_;
wire _00036_;
wire _00037_;
wire _00038_;
wire _00039_;
wire _00040_;
wire _00041_;
wire _00042_;
wire _00043_;
wire _00044_;
wire _00045_;
wire _00046_;
wire _00047_;
wire _00048_;
wire _00049_;
wire _00050_;
wire _00051_;
wire _00052_;
wire _00053_;
wire _00054_;
wire _00055_;
wire _00056_;
wire _00057_;
wire _00058_;
wire _00059_;
wire _00060_;
wire _00061_;
wire _00062_;
wire _00063_;
wire _00064_;
wire _00065_;
wire _00066_;
wire _00067_;
wire _00068_;
wire _00069_;
wire _00070_;
wire _00071_;
wire _00072_;
wire _00073_;
wire _00074_;
wire _00075_;
wire _00076_;
wire _00077_;
wire _00078_;
wire _00079_;
wire _00080_;
wire _00081_;
wire _00082_;
wire _00083_;
wire _00084_;
wire _00085_;
wire _00086_;
wire _00087_;
wire _00088_;
wire _00089_;
wire _00090_;
wire _00091_;
wire _00092_;
wire _00093_;
wire _00094_;
wire _00095_;
wire _00096_;
wire _00097_;
wire _00098_;
wire _00099_;
wire _00100_;
wire _00101_;
wire _00102_;
wire _00103_;
wire _00104_;
wire _00105_;
wire _00106_;
wire _00107_;
wire _00108_;
wire _00109_;
wire _00110_;
wire _00111_;
wire _00112_;
wire _00113_;
wire _00114_;
wire _00115_;
wire _00116_;
wire _00117_;
wire _00118_;
wire _00119_;
wire _00120_;
wire _00121_;
wire _00122_;
wire _00123_;
wire _00124_;
wire _00125_;
wire _00126_;
wire _00127_;
wire _00128_;
wire _00129_;
wire _00130_;
wire _00131_;
wire _00132_;
wire _00133_;
wire _00134_;
wire _00135_;
wire _00136_;
wire _00137_;
wire _00138_;
wire _00139_;
wire _00140_;
wire _00141_;
wire _00142_;
wire _00143_;
wire _00144_;
wire _00145_;
wire _00146_;
wire _00147_;
wire _00148_;
wire _00149_;
wire _00150_;
wire _00151_;
wire _00152_;
wire _00153_;
wire _00154_;
wire _00155_;
wire _00156_;
wire _00157_;
wire _00158_;
wire _00159_;
wire _00160_;
wire _00161_;
wire _00162_;
wire _00163_;
wire _00164_;
wire _00165_;
wire _00166_;
wire _00167_;
wire _00168_;
wire _00169_;
wire _00170_;
wire _00171_;
wire _00172_;
wire _00173_;
wire _00174_;
wire _00175_;
wire _00176_;
wire _00177_;
wire _00178_;
wire _00179_;
wire _00180_;
wire _00181_;
wire _00182_;
wire _00183_;
wire _00184_;
wire _00185_;
wire _00186_;
wire _00187_;
wire _00188_;
wire _00189_;
wire _00190_;
wire _00191_;
wire _00192_;
wire _00193_;
wire _00194_;
wire _00195_;
wire _00196_;
wire _00197_;
wire _00198_;
wire _00199_;
wire _00200_;
wire _00201_;
wire _00202_;
wire _00203_;
wire _00204_;
wire _00205_;
wire _00206_;
wire _00207_;
wire _00208_;
wire _00209_;
wire _00210_;
wire _00211_;
wire _00212_;
wire _00213_;
wire _00214_;
wire _00215_;
wire _00216_;
wire _00217_;
wire _00218_;
wire _00219_;
wire _00220_;
wire _00221_;
wire _00222_;
wire _00223_;
wire _00224_;
wire _00225_;
wire _00226_;
wire _00227_;
wire _00228_;
wire _00229_;
wire _00230_;
wire _00231_;
wire _00232_;
wire _00233_;
wire _00234_;
wire _00235_;
wire _00236_;
wire _00237_;
wire _00238_;
wire _00239_;
wire _00240_;
wire _00241_;
wire _00242_;
wire _00243_;
wire _00244_;
wire _00245_;
wire _00246_;
wire _00247_;
wire _00248_;
wire _00249_;
wire _00250_;
wire _00251_;
wire _00252_;
wire _00253_;
wire _00254_;
wire _00255_;
wire _00256_;
wire _00257_;
wire _00258_;
wire _00259_;
wire _00260_;
wire _00261_;
wire _00262_;
wire _00263_;
wire _00264_;
wire _00265_;
wire _00266_;
wire _00267_;
wire _00268_;
wire _00269_;
wire _00270_;
wire _00271_;
wire _00272_;
wire _00273_;
wire _00274_;
wire _00275_;
wire _00276_;
wire _00277_;
wire _00278_;
wire _00279_;
wire _00280_;
wire _00281_;
wire _00282_;
wire _00283_;
wire _00284_;
wire _00285_;
wire _00286_;
wire _00287_;
wire _00288_;
wire _00289_;
wire _00290_;
wire _00291_;
wire _00292_;
wire _00293_;
wire _00294_;
wire _00295_;
wire _00296_;
wire _00297_;
wire _00298_;
wire _00299_;
wire _00300_;
wire _00301_;
wire _00302_;
wire _00303_;
wire _00304_;
wire _00305_;
wire _00306_;
wire _00307_;
wire _00308_;
wire _00309_;
wire _00310_;
wire _00311_;
wire _00312_;
wire _00313_;
wire _00314_;
wire _00315_;
wire _00316_;
wire _00317_;
wire _00318_;
wire _00319_;
wire _00320_;
wire _00321_;
wire _00322_;
wire _00323_;
wire _00324_;
wire _00325_;
wire _00326_;
wire _00327_;
wire _00328_;
wire _00329_;
wire _00330_;
wire _00331_;
wire _00332_;
wire _00333_;
wire _00334_;
wire _00335_;
wire _00336_;
wire _00337_;
wire _00338_;
wire _00339_;
wire _00340_;
wire _00341_;
wire _00342_;
wire _00343_;
wire _00344_;
wire _00345_;
wire _00346_;
wire _00347_;
wire _00348_;
wire _00349_;
wire _00350_;
wire _00351_;
wire _00352_;
wire _00353_;
wire _00354_;
wire _00355_;
wire _00356_;
wire _00357_;
wire _00358_;
wire _00359_;
wire _00360_;
wire _00361_;
wire _00362_;
wire _00363_;
wire _00364_;
wire _00365_;
wire _00366_;
wire _00367_;
wire _00368_;
wire _00369_;
wire _00370_;
wire _00371_;
wire _00372_;
wire _00373_;
wire _00374_;
wire _00375_;
wire _00376_;
wire _00377_;
wire _00378_;
wire _00379_;
wire _00380_;
wire _00381_;
wire _00382_;
wire _00383_;
wire _00384_;
wire _00385_;
wire _00386_;
wire _00387_;
wire _00388_;
wire _00389_;
wire _00390_;
wire _00391_;
wire _00392_;
wire _00393_;
wire _00394_;
wire _00395_;
wire _00396_;
wire _00397_;
wire _00398_;
wire _00399_;
wire _00400_;
wire _00401_;
wire _00402_;
wire _00403_;
wire _00404_;
wire _00405_;
wire _00406_;
wire _00407_;
wire _00408_;
wire _00409_;
wire _00410_;
wire _00411_;
wire _00412_;
wire _00413_;
wire _00414_;
wire _00415_;
wire _00416_;
wire _00417_;
wire _00418_;
wire _00419_;
wire _00420_;
wire _00421_;
wire _00422_;
wire _00423_;
wire _00424_;
wire _00425_;
wire _00426_;
wire _00427_;
wire _00428_;
wire _00429_;
wire _00430_;
wire _00431_;
wire _00432_;
wire _00433_;
wire _00434_;
wire _00435_;
wire _00436_;
wire _00437_;
wire _00438_;
wire _00439_;
wire _00440_;
wire _00441_;
wire _00442_;
wire _00443_;
wire _00444_;
wire _00445_;
wire _00446_;
wire _00447_;
wire _00448_;
wire _00449_;
wire _00450_;
wire _00451_;
wire _00452_;
wire _00453_;
wire _00454_;
wire _00455_;
wire _00456_;
wire _00457_;
wire _00458_;
wire _00459_;
wire _00460_;
wire _00461_;
wire _00462_;
wire _00463_;
wire _00464_;
wire _00465_;
wire _00466_;
wire _00467_;
wire _00468_;
wire _00469_;
wire _00470_;
wire _00471_;
wire _00472_;
wire _00473_;
wire _00474_;
wire _00475_;
wire _00476_;
wire _00477_;
wire _00478_;
wire _00479_;
wire _00480_;
wire _00481_;
wire _00482_;
wire _00483_;
wire _00484_;
wire _00485_;
wire _00486_;
wire _00487_;
wire _00488_;
wire _00489_;
wire _00490_;
wire _00491_;
wire _00492_;
wire _00493_;
wire _00494_;
wire _00495_;
wire _00496_;
wire _00497_;
wire _00498_;
wire _00499_;
wire _00500_;
wire _00501_;
wire _00502_;
wire _00503_;
wire _00504_;
wire _00505_;
wire _00506_;
wire _00507_;
wire _00508_;
wire _00509_;
wire _00510_;
wire _00511_;
wire _00512_;
wire _00513_;
wire _00514_;
wire _00515_;
wire _00516_;
wire _00517_;
wire _00518_;
wire _00519_;
wire _00520_;
wire _00521_;
wire _00522_;
wire _00523_;
wire _00524_;
wire _00525_;
wire _00526_;
wire _00527_;
wire _00528_;
wire _00529_;
wire _00530_;
wire _00531_;
wire _00532_;
wire _00533_;
wire _00534_;
wire _00535_;
wire _00536_;
wire _00537_;
wire _00538_;
wire _00539_;
wire _00540_;
wire _00541_;
wire _00542_;
wire _00543_;
wire _00544_;
wire _00545_;
wire _00546_;
wire _00547_;
wire _00548_;
wire _00549_;
wire _00550_;
wire _00551_;
wire _00552_;
wire _00553_;
wire _00554_;
wire _00555_;
wire _00556_;
wire _00557_;
wire _00558_;
wire _00559_;
wire _00560_;
wire _00561_;
wire _00562_;
wire _00563_;
wire _00564_;
wire _00565_;
wire _00566_;
wire _00567_;
wire _00568_;
wire _00569_;
wire _00570_;
wire _00571_;
wire _00572_;
wire _00573_;
wire _00574_;
wire _00575_;
wire _00576_;
wire _00577_;
wire _00578_;
wire _00579_;
wire _00580_;
wire _00581_;
wire _00582_;
wire _00583_;
wire _00584_;
wire _00585_;
wire _00586_;
wire _00587_;
wire _00588_;
wire _00589_;
wire _00590_;
wire _00591_;
wire _00592_;
wire _00593_;
wire _00594_;
wire _00595_;
wire _00596_;
wire _00597_;
wire _00598_;
wire _00599_;
wire _00600_;
wire _00601_;
wire _00602_;
wire _00603_;
wire _00604_;
wire _00605_;
wire _00606_;
wire _00607_;
wire _00608_;
wire _00609_;
wire _00610_;
wire _00611_;
wire _00612_;
wire _00613_;
wire _00614_;
wire _00615_;
wire _00616_;
wire _00617_;
wire _00618_;
wire _00619_;
wire _00620_;
wire _00621_;
wire _00622_;
wire _00623_;
wire _00624_;
wire _00625_;
wire _00626_;
wire _00627_;
wire _00628_;
wire _00629_;
wire _00630_;
wire _00631_;
wire _00632_;
wire _00633_;
wire _00634_;
wire _00635_;
wire _00636_;
wire _00637_;
wire _00638_;
wire _00639_;
wire _00640_;
wire _00641_;
wire _00642_;
wire _00643_;
wire _00644_;
wire _00645_;
wire _00646_;
wire _00647_;
wire _00648_;
wire _00649_;
wire _00650_;
wire _00651_;
wire _00652_;
wire _00653_;
wire _00654_;
wire _00655_;
wire _00656_;
wire _00657_;
wire _00658_;
wire _00659_;
wire _00660_;
wire _00661_;
wire _00662_;
wire _00663_;
wire _00664_;
wire _00665_;
wire _00666_;
wire _00667_;
wire _00668_;
wire _00669_;
wire _00670_;
wire _00671_;
wire _00672_;
wire _00673_;
wire _00674_;
wire _00675_;
wire _00676_;
wire _00677_;
wire _00678_;
wire _00679_;
wire _00680_;
wire _00681_;
wire _00682_;
wire _00683_;
wire _00684_;
wire _00685_;
wire _00686_;
wire _00687_;
wire _00688_;
wire _00689_;
wire _00690_;
wire _00691_;
wire _00692_;
wire _00693_;
wire _00694_;
wire _00695_;
wire _00696_;
wire _00697_;
wire _00698_;
wire _00699_;
wire _00700_;
wire _00701_;
wire _00702_;
wire _00703_;
wire _00704_;
wire _00705_;
wire _00706_;
wire _00707_;
wire _00708_;
wire _00709_;
wire _00710_;
wire _00711_;
wire _00712_;
wire _00713_;
wire _00714_;
wire _00715_;
wire _00716_;
wire _00717_;
wire _00718_;
wire _00719_;
wire _00720_;
wire _00721_;
wire _00722_;
wire _00723_;
wire _00724_;
wire _00725_;
wire _00726_;
wire _00727_;
wire _00728_;
wire _00729_;
wire _00730_;
wire _00731_;
wire _00732_;
wire _00733_;
wire _00734_;
wire _00735_;
wire _00736_;
wire _00737_;
wire _00738_;
wire _00739_;
wire _00740_;
wire _00741_;
wire _00742_;
wire _00743_;
wire _00744_;
wire _00745_;
wire _00746_;
wire _00747_;
wire _00748_;
wire _00749_;
wire _00750_;
wire _00751_;
wire _00752_;
wire _00753_;
wire _00754_;
wire _00755_;
wire _00756_;
wire _00757_;
wire _00758_;
wire _00759_;
wire _00760_;
wire _00761_;
wire _00762_;
wire _00763_;
wire _00764_;
wire _00765_;
wire _00766_;
wire _00767_;
wire _00768_;
wire _00769_;
wire _00770_;
wire _00771_;
wire _00772_;
wire _00773_;
wire _00774_;
wire _00775_;
wire _00776_;
wire _00777_;
wire _00778_;
wire _00779_;
wire _00780_;
wire _00781_;
wire _00782_;
wire _00783_;
wire _00784_;
wire _00785_;
wire _00786_;
wire _00787_;
wire _00788_;
wire _00789_;
wire _00790_;
wire _00791_;
wire _00792_;
wire _00793_;
wire _00794_;
wire _00795_;
wire _00796_;
wire _00797_;
wire _00798_;
wire _00799_;
wire _00800_;
wire _00801_;
wire _00802_;
wire _00803_;
wire _00804_;
wire _00805_;
wire _00806_;
wire _00807_;
wire _00808_;
wire _00809_;
wire _00810_;
wire _00811_;
wire _00812_;
wire _00813_;
wire _00814_;
wire _00815_;
wire _00816_;
wire _00817_;
wire _00818_;
wire _00819_;
wire _00820_;
wire _00821_;
wire _00822_;
wire _00823_;
wire _00824_;
wire _00825_;
wire _00826_;
wire _00827_;
wire _00828_;
wire _00829_;
wire _00830_;
wire _00831_;
wire _00832_;
wire _00833_;
wire _00834_;
wire _00835_;
wire _00836_;
wire _00837_;
wire _00838_;
wire _00839_;
wire _00840_;
wire _00841_;
wire _00842_;
wire _00843_;
wire _00844_;
wire _00845_;
wire _00846_;
wire _00847_;
wire _00848_;
wire _00849_;
wire _00850_;
wire _00851_;
wire _00852_;
wire _00853_;
wire _00854_;
wire _00855_;
wire _00856_;
wire _00857_;
wire _00858_;
wire _00859_;
wire _00860_;
wire _00861_;
wire _00862_;
wire _00863_;
wire _00864_;
wire _00865_;
wire _00866_;
wire _00867_;
wire _00868_;
wire _00869_;
wire _00870_;
wire _00871_;
wire _00872_;
wire _00873_;
wire _00874_;
wire _00875_;
wire _00876_;
wire _00877_;
wire _00878_;
wire _00879_;
wire _00880_;
wire _00881_;
wire _00882_;
wire _00883_;
wire _00884_;
wire _00885_;
wire _00886_;
wire _00887_;
wire _00888_;
wire _00889_;
wire _00890_;
wire _00891_;
wire _00892_;
wire _00893_;
wire _00894_;
wire _00895_;
wire _00896_;
wire _00897_;
wire _00898_;
wire _00899_;
wire _00900_;
wire _00901_;
wire _00902_;
wire _00903_;
wire _00904_;
wire _00905_;
wire _00906_;
wire _00907_;
wire _00908_;
wire _00909_;
wire _00910_;
wire _00911_;
wire _00912_;
wire _00913_;
wire _00914_;
wire _00915_;
wire _00916_;
wire _00917_;
wire _00918_;
wire _00919_;
wire _00920_;
wire _00921_;
wire _00922_;
wire _00923_;
wire _00924_;
wire _00925_;
wire _00926_;
wire _00927_;
wire _00928_;
wire _00929_;
wire _00930_;
wire _00931_;
wire _00932_;
wire _00933_;
wire _00934_;
wire _00935_;
wire _00936_;
wire _00937_;
wire _00938_;
wire _00939_;
wire _00940_;
wire _00941_;
wire _00942_;
wire _00943_;
wire _00944_;
wire _00945_;
wire _00946_;
wire _00947_;
wire _00948_;
wire _00949_;
wire _00950_;
wire _00951_;
wire _00952_;
wire _00953_;
wire _00954_;
wire _00955_;
wire _00956_;
wire _00957_;
wire _00958_;
wire _00959_;
wire _00960_;
wire _00961_;
wire _00962_;
wire _00963_;
wire _00964_;
wire _00965_;
wire _00966_;
wire _00967_;
wire _00968_;
wire _00969_;
wire _00970_;
wire _00971_;
wire _00972_;
wire _00973_;
wire _00974_;
wire _00975_;
wire _00976_;
wire _00977_;
wire _00978_;
wire _00979_;
wire _00980_;
wire _00981_;
wire _00982_;
wire _00983_;
wire _00984_;
wire _00985_;
wire _00986_;
wire _00987_;
wire _00988_;
wire _00989_;
wire _00990_;
wire _00991_;
wire _00992_;
wire _00993_;
wire _00994_;
wire _00995_;
wire _00996_;
wire _00997_;
wire _00998_;
wire _00999_;
wire _01000_;
wire _01001_;
wire _01002_;
wire _01003_;
wire _01004_;
wire _01005_;
wire _01006_;
wire _01007_;
wire _01008_;
wire _01009_;
wire _01010_;
wire _01011_;
wire _01012_;
wire _01013_;
wire _01014_;
wire _01015_;
wire _01016_;
wire _01017_;
wire _01018_;
wire _01019_;
wire _01020_;
wire _01021_;
wire _01022_;
wire _01023_;
wire _01024_;
wire _01025_;
wire _01026_;
wire _01027_;
wire _01028_;
wire _01029_;
wire _01030_;
wire _01031_;
wire _01032_;
wire _01033_;
wire _01034_;
wire _01035_;
wire _01036_;
wire _01037_;
wire _01038_;
wire _01039_;
wire _01040_;
wire _01041_;
wire _01042_;
wire _01043_;
wire _01044_;
wire _01045_;
wire _01046_;
wire _01047_;
wire _01048_;
wire _01049_;
wire _01050_;
wire _01051_;
wire _01052_;
wire _01053_;
wire _01054_;
wire _01055_;
wire _01056_;
wire _01057_;
wire _01058_;
wire _01059_;
wire _01060_;
wire _01061_;
wire _01062_;
wire _01063_;
wire _01064_;
wire _01065_;
wire _01066_;
wire _01067_;
wire _01068_;
wire _01069_;
wire _01070_;
wire _01071_;
wire _01072_;
wire _01073_;
wire _01074_;
wire _01075_;
wire _01076_;
wire _01077_;
wire _01078_;
wire _01079_;
wire _01080_;
wire _01081_;
wire _01082_;
wire _01083_;
wire _01084_;
wire _01085_;
wire _01086_;
wire _01087_;
wire _01088_;
wire _01089_;
wire _01090_;
wire _01091_;
wire _01092_;
wire _01093_;
wire _01094_;
wire _01095_;
wire _01096_;
wire _01097_;
wire _01098_;
wire _01099_;
wire _01100_;
wire _01101_;
wire _01102_;
wire _01103_;
wire _01104_;
wire _01105_;
wire _01106_;
wire _01107_;
wire _01108_;
wire _01109_;
wire _01110_;
wire _01111_;
wire _01112_;
wire _01113_;
wire _01114_;
wire _01115_;
wire _01116_;
wire _01117_;
wire _01118_;
wire _01119_;
wire _01120_;
wire _01121_;
wire _01122_;
wire _01123_;
wire _01124_;
wire _01125_;
wire _01126_;
wire _01127_;
wire _01128_;
wire _01129_;
wire _01130_;
wire _01131_;
wire _01132_;
wire _01133_;
wire _01134_;
wire _01135_;
wire _01136_;
wire _01137_;
wire _01138_;
wire _01139_;
wire _01140_;
wire _01141_;
wire _01142_;
wire _01143_;
wire _01144_;
wire _01145_;
wire _01146_;
wire _01147_;
wire _01148_;
wire _01149_;
wire _01150_;
wire _01151_;
wire _01152_;
wire _01153_;
wire _01154_;
wire _01155_;
wire _01156_;
wire _01157_;
wire _01158_;
wire _01159_;
wire _01160_;
wire _01161_;
wire _01162_;
wire _01163_;
wire _01164_;
wire _01165_;
wire _01166_;
wire _01167_;
wire _01168_;
wire _01169_;
wire _01170_;
wire _01171_;
wire _01172_;
wire _01173_;
wire _01174_;
wire _01175_;
wire _01176_;
wire _01177_;
wire _01178_;
wire _01179_;
wire _01180_;
wire _01181_;
wire _01182_;
wire _01183_;
wire _01184_;
wire _01185_;
wire _01186_;
wire _01187_;
wire _01188_;
wire _01189_;
wire _01190_;
wire _01191_;
wire _01192_;
wire _01193_;
wire _01194_;
wire _01195_;
wire _01196_;
wire _01197_;
wire _01198_;
wire _01199_;
wire _01200_;
wire _01201_;
wire _01202_;
wire _01203_;
wire _01204_;
wire _01205_;
wire _01206_;
wire _01207_;
wire _01208_;
wire _01209_;
wire _01210_;
wire _01211_;
wire _01212_;
wire _01213_;
wire _01214_;
wire _01215_;
wire _01216_;
wire _01217_;
wire _01218_;
wire _01219_;
wire _01220_;
wire _01221_;
wire _01222_;
wire _01223_;
wire _01224_;
wire _01225_;
wire _01226_;
wire _01227_;
wire _01228_;
wire _01229_;
wire _01230_;
wire _01231_;
wire _01232_;
wire _01233_;
wire _01234_;
wire _01235_;
wire _01236_;
wire _01237_;
wire _01238_;
wire _01239_;
wire _01240_;
wire _01241_;
wire _01242_;
wire _01243_;
wire _01244_;
wire _01245_;
wire _01246_;
wire _01247_;
wire _01248_;
wire _01249_;
wire _01250_;
wire _01251_;
wire _01252_;
wire _01253_;
wire _01254_;
wire _01255_;
wire _01256_;
wire _01257_;
wire _01258_;
wire _01259_;
wire _01260_;
wire _01261_;
wire _01262_;
wire _01263_;
wire _01264_;
wire _01265_;
wire _01266_;
wire _01267_;
wire _01268_;
wire _01269_;
wire _01270_;
wire _01271_;
wire _01272_;
wire _01273_;
wire _01274_;
wire _01275_;
wire _01276_;
wire _01277_;
wire _01278_;
wire _01279_;
wire _01280_;
wire _01281_;
wire _01282_;
wire _01283_;
wire _01284_;
wire _01285_;
wire _01286_;
wire _01287_;
wire _01288_;
wire _01289_;
wire _01290_;
wire _01291_;
wire _01292_;
wire _01293_;
wire _01294_;
wire _01295_;
wire _01296_;
wire _01297_;
wire _01298_;
wire _01299_;
wire _01300_;
wire _01301_;
wire _01302_;
wire _01303_;
wire _01304_;
wire _01305_;
wire _01306_;
wire _01307_;
wire _01308_;
wire _01309_;
wire _01310_;
wire _01311_;
wire _01312_;
wire _01313_;
wire _01314_;
wire _01315_;
wire _01316_;
wire _01317_;
wire _01318_;
wire _01319_;
wire _01320_;
wire _01321_;
wire _01322_;
wire _01323_;
wire _01324_;
wire _01325_;
wire _01326_;
wire _01327_;
wire _01328_;
wire _01329_;
wire _01330_;
wire _01331_;
wire _01332_;
wire _01333_;
wire _01334_;
wire _01335_;
wire _01336_;
wire _01337_;
wire _01338_;
wire _01339_;
wire _01340_;
wire _01341_;
wire _01342_;
wire _01343_;
wire _01344_;
wire _01345_;
wire _01346_;
wire _01347_;
wire _01348_;
wire _01349_;
wire _01350_;
wire _01351_;
wire _01352_;
wire _01353_;
wire _01354_;
wire _01355_;
wire _01356_;
wire _01357_;
wire _01358_;
wire _01359_;
wire _01360_;
wire _01361_;
wire _01362_;
wire _01363_;
wire _01364_;
wire _01365_;
wire _01366_;
wire _01367_;
wire _01368_;
wire _01369_;
wire _01370_;
wire _01371_;
wire _01372_;
wire _01373_;
wire _01374_;
wire _01375_;
wire _01376_;
wire _01377_;
wire _01378_;
wire _01379_;
wire _01380_;
wire _01381_;
wire _01382_;
wire _01383_;
wire _01384_;
wire _01385_;
wire _01386_;
wire _01387_;
wire _01388_;
wire _01389_;
wire _01390_;
wire _01391_;
wire _01392_;
wire _01393_;
wire _01394_;
wire _01395_;
wire _01396_;
wire _01397_;
wire _01398_;
wire _01399_;
wire _01400_;
wire _01401_;
wire _01402_;
wire _01403_;
wire _01404_;
wire _01405_;
wire _01406_;
wire _01407_;
wire _01408_;
wire _01409_;
wire _01410_;
wire _01411_;
wire _01412_;
wire _01413_;
wire _01414_;
wire _01415_;
wire _01416_;
wire _01417_;
wire _01418_;
wire _01419_;
wire _01420_;
wire _01421_;
wire _01422_;
wire _01423_;
wire _01424_;
wire _01425_;
wire _01426_;
wire _01427_;
wire _01428_;
wire _01429_;
wire _01430_;
wire _01431_;
wire _01432_;
wire _01433_;
wire _01434_;
wire _01435_;
wire _01436_;
wire _01437_;
wire _01438_;
wire _01439_;
wire _01440_;
wire _01441_;
wire _01442_;
wire _01443_;
wire _01444_;
wire _01445_;
wire _01446_;
wire _01447_;
wire _01448_;
wire _01449_;
wire _01450_;
wire _01451_;
wire _01452_;
wire _01453_;
wire _01454_;
wire _01455_;
wire _01456_;
wire _01457_;
wire _01458_;
wire _01459_;
wire _01460_;
wire _01461_;
wire _01462_;
wire _01463_;
wire _01464_;
wire _01465_;
wire _01466_;
wire _01467_;
wire _01468_;
wire _01469_;
wire _01470_;
wire _01471_;
wire _01472_;
wire _01473_;
wire _01474_;
wire _01475_;
wire _01476_;
wire _01477_;
wire _01478_;
wire _01479_;
wire _01480_;
wire _01481_;
wire _01482_;
wire _01483_;
wire _01484_;
wire _01485_;
wire _01486_;
wire _01487_;
wire _01488_;
wire _01489_;
wire _01490_;
wire _01491_;
wire _01492_;
wire _01493_;
wire _01494_;
wire _01495_;
wire _01496_;
wire _01497_;
wire _01498_;
wire _01499_;
wire _01500_;
wire _01501_;
wire _01502_;
wire _01503_;
wire _01504_;
wire _01505_;
wire _01506_;
wire _01507_;
wire _01508_;
wire _01509_;
wire _01510_;
wire _01511_;
wire _01512_;
wire _01513_;
wire _01514_;
wire _01515_;
wire _01516_;
wire _01517_;
wire _01518_;
wire _01519_;
wire _01520_;
wire _01521_;
wire _01522_;
wire _01523_;
wire _01524_;
wire _01525_;
wire _01526_;
wire _01527_;
wire _01528_;
wire _01529_;
wire _01530_;
wire _01531_;
wire _01532_;
wire _01533_;
wire _01534_;
wire _01535_;
wire _01536_;
wire _01537_;
wire _01538_;
wire _01539_;
wire _01540_;
wire _01541_;
wire _01542_;
wire _01543_;
wire _01544_;
wire _01545_;
wire _01546_;
wire _01547_;
wire _01548_;
wire _01549_;
wire _01550_;
wire _01551_;
wire _01552_;
wire _01553_;
wire _01554_;
wire _01555_;
wire _01556_;
wire _01557_;
wire _01558_;
wire _01559_;
wire _01560_;
wire _01561_;
wire _01562_;
wire _01563_;
wire _01564_;
wire _01565_;
wire _01566_;
wire _01567_;
wire _01568_;
wire _01569_;
wire _01570_;
wire _01571_;
wire _01572_;
wire _01573_;
wire _01574_;
wire _01575_;
wire _01576_;
wire _01577_;
wire _01578_;
wire _01579_;
wire _01580_;
wire _01581_;
wire _01582_;
wire _01583_;
wire _01584_;
wire _01585_;
wire _01586_;
wire _01587_;
wire _01588_;
wire _01589_;
wire _01590_;
wire _01591_;
wire _01592_;
wire _01593_;
wire _01594_;
wire _01595_;
wire _01596_;
wire _01597_;
wire _01598_;
wire _01599_;
wire _01600_;
wire _01601_;
wire _01602_;
wire _01603_;
wire _01604_;
wire _01605_;
wire _01606_;
wire _01607_;
wire _01608_;
wire _01609_;
wire _01610_;
wire _01611_;
wire _01612_;
wire _01613_;
wire _01614_;
wire _01615_;
wire _01616_;
wire _01617_;
wire _01618_;
wire _01619_;
wire _01620_;
wire _01621_;
wire _01622_;
wire _01623_;
wire _01624_;
wire _01625_;
wire _01626_;
wire _01627_;
wire _01628_;
wire _01629_;
wire _01630_;
wire _01631_;
wire _01632_;
wire _01633_;
wire _01634_;
wire _01635_;
wire _01636_;
wire _01637_;
wire _01638_;
wire _01639_;
wire _01640_;
wire _01641_;
wire _01642_;
wire _01643_;
wire _01644_;
wire _01645_;
wire _01646_;
wire _01647_;
wire _01648_;
wire _01649_;
wire _01650_;
wire _01651_;
wire _01652_;
wire _01653_;
wire _01654_;
wire _01655_;
wire _01656_;
wire _01657_;
wire _01658_;
wire _01659_;
wire _01660_;
wire _01661_;
wire _01662_;
wire _01663_;
wire _01664_;
wire _01665_;
wire _01666_;
wire _01667_;
wire _01668_;
wire _01669_;
wire _01670_;
wire _01671_;
wire _01672_;
wire _01673_;
wire _01674_;
wire _01675_;
wire _01676_;
wire _01677_;
wire _01678_;
wire _01679_;
wire _01680_;
wire _01681_;
wire _01682_;
wire _01683_;
wire _01684_;
wire _01685_;
wire _01686_;
wire _01687_;
wire _01688_;
wire _01689_;
wire _01690_;
wire _01691_;
wire _01692_;
wire _01693_;
wire _01694_;
wire _01695_;
wire _01696_;
wire _01697_;
wire _01698_;
wire _01699_;
wire _01700_;
wire _01701_;
wire _01702_;
wire _01703_;
wire _01704_;
wire _01705_;
wire _01706_;
wire _01707_;
wire _01708_;
wire _01709_;
wire _01710_;
wire _01711_;
wire _01712_;
wire _01713_;
wire _01714_;
wire _01715_;
wire _01716_;
wire _01717_;
wire _01718_;
wire _01719_;
wire _01720_;
wire _01721_;
wire _01722_;
wire _01723_;
wire _01724_;
wire _01725_;
wire _01726_;
wire _01727_;
wire _01728_;
wire _01729_;
wire _01730_;
wire _01731_;
wire _01732_;
wire _01733_;
wire _01734_;
wire _01735_;
wire _01736_;
wire _01737_;
wire _01738_;
wire _01739_;
wire _01740_;
wire _01741_;
wire _01742_;
wire _01743_;
wire _01744_;
wire _01745_;
wire _01746_;
wire _01747_;
wire _01748_;
wire _01749_;
wire _01750_;
wire _01751_;
wire _01752_;
wire _01753_;
wire _01754_;
wire _01755_;
wire _01756_;
wire _01757_;
wire _01758_;
wire _01759_;
wire _01760_;
wire _01761_;
wire _01762_;
wire _01763_;
wire _01764_;
wire _01765_;
wire _01766_;
wire _01767_;
wire _01768_;
wire _01769_;
wire _01770_;
wire _01771_;
wire _01772_;
wire _01773_;
wire _01774_;
wire _01775_;
wire _01776_;
wire _01777_;
wire _01778_;
wire _01779_;
wire _01780_;
wire _01781_;
wire _01782_;
wire _01783_;
wire _01784_;
wire _01785_;
wire _01786_;
wire _01787_;
wire _01788_;
wire _01789_;
wire _01790_;
wire _01791_;
wire _01792_;
wire _01793_;
wire _01794_;
wire _01795_;
wire _01796_;
wire _01797_;
wire _01798_;
wire _01799_;
wire _01800_;
wire _01801_;
wire _01802_;
wire _01803_;
wire _01804_;
wire _01805_;
wire _01806_;
wire _01807_;
wire _01808_;
wire _01809_;
wire _01810_;
wire _01811_;
wire _01812_;
wire _01813_;
wire _01814_;
wire _01815_;
wire _01816_;
wire _01817_;
wire _01818_;
wire _01819_;
wire _01820_;
wire _01821_;
wire _01822_;
wire _01823_;
wire _01824_;
wire _01825_;
wire _01826_;
wire _01827_;
wire _01828_;
wire _01829_;
wire _01830_;
wire _01831_;
wire _01832_;
wire _01833_;
wire _01834_;
wire _01835_;
wire _01836_;
wire _01837_;
wire _01838_;
wire _01839_;
wire _01840_;
wire _01841_;
wire _01842_;
wire _01843_;
wire _01844_;
wire _01845_;
wire _01846_;
wire _01847_;
wire _01848_;
wire _01849_;
wire _01850_;
wire _01851_;
wire _01852_;
wire _01853_;
wire _01854_;
wire _01855_;
wire _01856_;
wire _01857_;
wire _01858_;
wire _01859_;
wire _01860_;
wire _01861_;
wire _01862_;
wire _01863_;
wire _01864_;
wire _01865_;
wire _01866_;
wire _01867_;
wire _01868_;
wire _01869_;
wire _01870_;
wire _01871_;
wire _01872_;
wire _01873_;
wire _01874_;
wire _01875_;
wire _01876_;
wire _01877_;
wire _01878_;
wire _01879_;
wire _01880_;
wire _01881_;
wire _01882_;
wire _01883_;
wire _01884_;
wire _01885_;
wire _01886_;
wire _01887_;
wire _01888_;
wire _01889_;
wire _01890_;
wire _01891_;
wire _01892_;
wire _01893_;
wire _01894_;
wire _01895_;
wire _01896_;
wire _01897_;
wire _01898_;
wire _01899_;
wire _01900_;
wire _01901_;
wire _01902_;
wire _01903_;
wire _01904_;
wire _01905_;
wire _01906_;
wire _01907_;
wire _01908_;
wire _01909_;
wire _01910_;
wire _01911_;
wire _01912_;
wire _01913_;
wire _01914_;
wire _01915_;
wire _01916_;
wire _01917_;
wire _01918_;
wire _01919_;
wire _01920_;
wire _01921_;
wire _01922_;
wire _01923_;
wire _01924_;
wire _01925_;
wire _01926_;
wire _01927_;
wire _01928_;
wire _01929_;
wire _01930_;
wire _01931_;
wire _01932_;
wire _01933_;
wire _01934_;
wire _01935_;
wire _01936_;
wire _01937_;
wire _01938_;
wire _01939_;
wire _01940_;
wire _01941_;
wire _01942_;
wire _01943_;
wire _01944_;
wire _01945_;
wire _01946_;
wire _01947_;
wire _01948_;
wire _01949_;
wire _01950_;
wire _01951_;
wire _01952_;
wire _01953_;
wire _01954_;
wire _01955_;
wire _01956_;
wire _01957_;
wire _01958_;
wire _01959_;
wire _01960_;
wire _01961_;
wire _01962_;
wire _01963_;
wire _01964_;
wire _01965_;
wire _01966_;
wire _01967_;
wire _01968_;
wire _01969_;
wire _01970_;
wire _01971_;
wire _01972_;
wire _01973_;
wire _01974_;
wire _01975_;
wire _01976_;
wire _01977_;
wire _01978_;
wire _01979_;
wire _01980_;
wire _01981_;
wire _01982_;
wire _01983_;
wire _01984_;
wire _01985_;
wire _01986_;
wire _01987_;
wire _01988_;
wire _01989_;
wire _01990_;
wire _01991_;
wire _01992_;
wire _01993_;
wire _01994_;
wire _01995_;
wire _01996_;
wire _01997_;
wire _01998_;
wire _01999_;
wire _02000_;
wire _02001_;
wire _02002_;
wire _02003_;
wire _02004_;
wire _02005_;
wire _02006_;
wire _02007_;
wire _02008_;
wire _02009_;
wire _02010_;
wire _02011_;
wire _02012_;
wire _02013_;
wire _02014_;
wire _02015_;
wire _02016_;
wire _02017_;
wire _02018_;
wire _02019_;
wire _02020_;
wire _02021_;
wire _02022_;
wire _02023_;
wire _02024_;
wire _02025_;
wire _02026_;
wire _02027_;
wire _02028_;
wire _02029_;
wire _02030_;
wire _02031_;
wire _02032_;
wire _02033_;
wire _02034_;
wire _02035_;
wire _02036_;
wire _02037_;
wire _02038_;
wire _02039_;
wire _02040_;
wire _02041_;
wire _02042_;
wire _02043_;
wire _02044_;
wire _02045_;
wire _02046_;
wire _02047_;
wire _02048_;
wire _02049_;
wire _02050_;
wire _02051_;
wire _02052_;
wire _02053_;
wire _02054_;
wire _02055_;
wire _02056_;
wire _02057_;
wire _02058_;
wire _02059_;
wire _02060_;
wire _02061_;
wire _02062_;
wire _02063_;
wire _02064_;
wire _02065_;
wire _02066_;
wire _02067_;
wire _02068_;
wire _02069_;
wire _02070_;
wire _02071_;
wire _02072_;
wire _02073_;
wire _02074_;
wire _02075_;
wire _02076_;
wire _02077_;
wire _02078_;
wire _02079_;
wire _02080_;
wire _02081_;
wire _02082_;
wire _02083_;
wire _02084_;
wire _02085_;
wire _02086_;
wire _02087_;
wire _02088_;
wire _02089_;
wire _02090_;
wire _02091_;
wire _02092_;
wire _02093_;
wire _02094_;
wire _02095_;
wire _02096_;
wire _02097_;
wire _02098_;
wire _02099_;
wire _02100_;
wire _02101_;
wire _02102_;
wire _02103_;
wire _02104_;
wire _02105_;
wire _02106_;
wire _02107_;
wire _02108_;
wire _02109_;
wire _02110_;
wire _02111_;
wire _02112_;
wire _02113_;
wire _02114_;
wire _02115_;
wire _02116_;
wire _02117_;
wire _02118_;
wire _02119_;
wire _02120_;
wire _02121_;
wire _02122_;
wire _02123_;
wire _02124_;
wire _02125_;
wire _02126_;
wire _02127_;
wire _02128_;
wire _02129_;
wire _02130_;
wire _02131_;
wire _02132_;
wire _02133_;
wire _02134_;
wire _02135_;
wire _02136_;
wire _02137_;
wire _02138_;
wire _02139_;
wire _02140_;
wire _02141_;
wire _02142_;
wire _02143_;
wire _02144_;
wire _02145_;
wire _02146_;
wire _02147_;
wire _02148_;
wire _02149_;
wire _02150_;
wire _02151_;
wire _02152_;
wire _02153_;
wire _02154_;
wire _02155_;
wire _02156_;
wire _02157_;
wire _02158_;
wire _02159_;
wire _02160_;
wire _02161_;
wire _02162_;
wire _02163_;
wire _02164_;
wire _02165_;
wire _02166_;
wire _02167_;
wire _02168_;
wire _02169_;
wire _02170_;
wire _02171_;
wire _02172_;
wire _02173_;
wire _02174_;
wire _02175_;
wire _02176_;
wire _02177_;
wire _02178_;
wire _02179_;
wire _02180_;
wire _02181_;
wire _02182_;
wire _02183_;
wire _02184_;
wire _02185_;
wire _02186_;
wire _02187_;
wire _02188_;
wire _02189_;
wire _02190_;
wire _02191_;
wire _02192_;
wire _02193_;
wire _02194_;
wire _02195_;
wire _02196_;
wire _02197_;
wire _02198_;
wire _02199_;
wire _02200_;
wire _02201_;
wire _02202_;
wire _02203_;
wire _02204_;
wire _02205_;
wire _02206_;
wire _02207_;
wire _02208_;
wire _02209_;
wire _02210_;
wire _02211_;
wire _02212_;
wire _02213_;
wire _02214_;
wire _02215_;
wire _02216_;
wire _02217_;
wire _02218_;
wire _02219_;
wire _02220_;
wire _02221_;
wire _02222_;
wire _02223_;
wire _02224_;
wire _02225_;
wire _02226_;
wire _02227_;
wire _02228_;
wire _02229_;
wire _02230_;
wire _02231_;
wire _02232_;
wire _02233_;
wire _02234_;
wire _02235_;
wire _02236_;
wire _02237_;
wire _02238_;
wire _02239_;
wire _02240_;
wire _02241_;
wire _02242_;
wire _02243_;
wire _02244_;
wire _02245_;
wire _02246_;
wire _02247_;
wire _02248_;
wire _02249_;
wire _02250_;
wire _02251_;
wire _02252_;
wire _02253_;
wire _02254_;
wire _02255_;
wire _02256_;
wire _02257_;
wire _02258_;
wire _02259_;
wire _02260_;
wire _02261_;
wire _02262_;
wire _02263_;
wire _02264_;
wire _02265_;
wire _02266_;
wire _02267_;
wire _02268_;
wire _02269_;
wire _02270_;
wire _02271_;
wire _02272_;
wire _02273_;
wire _02274_;
wire _02275_;
wire _02276_;
wire _02277_;
wire _02278_;
wire _02279_;
wire _02280_;
wire _02281_;
wire _02282_;
wire _02283_;
wire _02284_;
wire _02285_;
wire _02286_;
wire _02287_;
wire _02288_;
wire _02289_;
wire _02290_;
wire _02291_;
wire _02292_;
wire _02293_;
wire _02294_;
wire _02295_;
wire _02296_;
wire _02297_;
wire _02298_;
wire _02299_;
wire _02300_;
wire _02301_;
wire _02302_;
wire _02303_;
wire _02304_;
wire _02305_;
wire _02306_;
wire _02307_;
wire _02308_;
wire _02309_;
wire _02310_;
wire _02311_;
wire _02312_;
wire _02313_;
wire _02314_;
wire _02315_;
wire _02316_;
wire _02317_;
wire _02318_;
wire _02319_;
wire _02320_;
wire _02321_;
wire _02322_;
wire _02323_;
wire _02324_;
wire _02325_;
wire _02326_;
wire _02327_;
wire _02328_;
wire _02329_;
wire _02330_;
wire _02331_;
wire _02332_;
wire _02333_;
wire _02334_;
wire _02335_;
wire _02336_;
wire _02337_;
wire _02338_;
wire _02339_;
wire _02340_;
wire _02341_;
wire _02342_;
wire _02343_;
wire _02344_;
wire _02345_;
wire _02346_;
wire _02347_;
wire _02348_;
wire _02349_;
wire _02350_;
wire _02351_;
wire _02352_;
wire _02353_;
wire _02354_;
wire _02355_;
wire _02356_;
wire _02357_;
wire _02358_;
wire _02359_;
wire _02360_;
wire _02361_;
wire _02362_;
wire _02363_;
wire _02364_;
wire _02365_;
wire _02366_;
wire _02367_;
wire _02368_;
wire _02369_;
wire _02370_;
wire _02371_;
wire _02372_;
wire _02373_;
wire _02374_;
wire _02375_;
wire _02376_;
wire _02377_;
wire _02378_;
wire _02379_;
wire _02380_;
wire _02381_;
wire _02382_;
wire _02383_;
wire _02384_;
wire _02385_;
wire _02386_;
wire _02387_;
wire _02388_;
wire _02389_;
wire _02390_;
wire _02391_;
wire _02392_;
wire _02393_;
wire _02394_;
wire _02395_;
wire _02396_;
wire _02397_;
wire _02398_;
wire _02399_;
wire _02400_;
wire _02401_;
wire _02402_;
wire _02403_;
wire _02404_;
wire _02405_;
wire _02406_;
wire _02407_;
wire _02408_;
wire _02409_;
wire _02410_;
wire _02411_;
wire _02412_;
wire _02413_;
wire _02414_;
wire _02415_;
wire _02416_;
wire _02417_;
wire _02418_;
wire _02419_;
wire _02420_;
wire _02421_;
wire _02422_;
wire _02423_;
wire _02424_;
wire _02425_;
wire _02426_;
wire _02427_;
wire _02428_;
wire _02429_;
wire _02430_;
wire _02431_;
wire _02432_;
wire _02433_;
wire _02434_;
wire _02435_;
wire _02436_;
wire _02437_;
wire _02438_;
wire _02439_;
wire _02440_;
wire _02441_;
wire _02442_;
wire _02443_;
wire _02444_;
wire _02445_;
wire _02446_;
wire _02447_;
wire _02448_;
wire _02449_;
wire _02450_;
wire _02451_;
wire _02452_;
wire _02453_;
wire _02454_;
wire _02455_;
wire _02456_;
wire _02457_;
wire _02458_;
wire _02459_;
wire _02460_;
wire _02461_;
wire _02462_;
wire _02463_;
wire _02464_;
wire _02465_;
wire _02466_;
wire _02467_;
wire _02468_;
wire _02469_;
wire _02470_;
wire _02471_;
wire _02472_;
wire _02473_;
wire _02474_;
wire _02475_;
wire _02476_;
wire _02477_;
wire _02478_;
wire _02479_;
wire _02480_;
wire _02481_;
wire _02482_;
wire _02483_;
wire _02484_;
wire _02485_;
wire _02486_;
wire _02487_;
wire _02488_;
wire _02489_;
wire _02490_;
wire _02491_;
wire _02492_;
wire _02493_;
wire _02494_;
wire _02495_;
wire _02496_;
wire _02497_;
wire _02498_;
wire _02499_;
wire _02500_;
wire _02501_;
wire _02502_;
wire _02503_;
wire _02504_;
wire _02505_;
wire _02506_;
wire _02507_;
wire _02508_;
wire _02509_;
wire _02510_;
wire _02511_;
wire _02512_;
wire _02513_;
wire _02514_;
wire _02515_;
wire _02516_;
wire _02517_;
wire _02518_;
wire _02519_;
wire _02520_;
wire _02521_;
wire _02522_;
wire _02523_;
wire _02524_;
wire _02525_;
wire _02526_;
wire _02527_;
wire _02528_;
wire _02529_;
wire _02530_;
wire _02531_;
wire _02532_;
wire _02533_;
wire _02534_;
wire _02535_;
wire _02536_;
wire _02537_;
wire _02538_;
wire _02539_;
wire _02540_;
wire _02541_;
wire _02542_;
wire _02543_;
wire _02544_;
wire _02545_;
wire _02546_;
wire _02547_;
wire _02548_;
wire _02549_;
wire _02550_;
wire _02551_;
wire _02552_;
wire _02553_;
wire _02554_;
wire _02555_;
wire _02556_;
wire _02557_;
wire _02558_;
wire _02559_;
wire _02560_;
wire _02561_;
wire _02562_;
wire _02563_;
wire _02564_;
wire _02565_;
wire _02566_;
wire _02567_;
wire _02568_;
wire _02569_;
wire _02570_;
wire _02571_;
wire _02572_;
wire _02573_;
wire _02574_;
wire _02575_;
wire _02576_;
wire _02577_;
wire _02578_;
wire _02579_;
wire _02580_;
wire _02581_;
wire _02582_;
wire _02583_;
wire _02584_;
wire _02585_;
wire _02586_;
wire _02587_;
wire _02588_;
wire _02589_;
wire _02590_;
wire _02591_;
wire _02592_;
wire _02593_;
wire _02594_;
wire _02595_;
wire _02596_;
wire _02597_;
wire _02598_;
wire _02599_;
wire _02600_;
wire _02601_;
wire _02602_;
wire _02603_;
wire _02604_;
wire _02605_;
wire _02606_;
wire _02607_;
wire _02608_;
wire _02609_;
wire _02610_;
wire _02611_;
wire _02612_;
wire _02613_;
wire _02614_;
wire _02615_;
wire _02616_;
wire _02617_;
wire _02618_;
wire _02619_;
wire _02620_;
wire _02621_;
wire _02622_;
wire _02623_;
wire _02624_;
wire _02625_;
wire _02626_;
wire _02627_;
wire _02628_;
wire _02629_;
wire _02630_;
wire _02631_;
wire _02632_;
wire _02633_;
wire _02634_;
wire _02635_;
wire _02636_;
wire _02637_;
wire _02638_;
wire _02639_;
wire _02640_;
wire _02641_;
wire _02642_;
wire _02643_;
wire _02644_;
wire _02645_;
wire _02646_;
wire _02647_;
wire _02648_;
wire _02649_;
wire _02650_;
wire _02651_;
wire _02652_;
wire _02653_;
wire _02654_;
wire _02655_;
wire _02656_;
wire _02657_;
wire _02658_;
wire _02659_;
wire _02660_;
wire _02661_;
wire _02662_;
wire _02663_;
wire _02664_;
wire _02665_;
wire _02666_;
wire _02667_;
wire _02668_;
wire _02669_;
wire _02670_;
wire _02671_;
wire _02672_;
wire _02673_;
wire _02674_;
wire _02675_;
wire _02676_;
wire _02677_;
wire _02678_;
wire _02679_;
wire _02680_;
wire _02681_;
wire _02682_;
wire _02683_;
wire _02684_;
wire _02685_;
wire _02686_;
wire _02687_;
wire _02688_;
wire _02689_;
wire _02690_;
wire _02691_;
wire _02692_;
wire _02693_;
wire _02694_;
wire _02695_;
wire _02696_;
wire _02697_;
wire _02698_;
wire _02699_;
wire _02700_;
wire _02701_;
wire _02702_;
wire _02703_;
wire _02704_;
wire _02705_;
wire _02706_;
wire _02707_;
wire _02708_;
wire _02709_;
wire _02710_;
wire _02711_;
wire _02712_;
wire _02713_;
wire _02714_;
wire _02715_;
wire _02716_;
wire _02717_;
wire _02718_;
wire _02719_;
wire _02720_;
wire _02721_;
wire _02722_;
wire _02723_;
wire _02724_;
wire _02725_;
wire _02726_;
wire _02727_;
wire _02728_;
wire _02729_;
wire _02730_;
wire _02731_;
wire _02732_;
wire _02733_;
wire _02734_;
wire _02735_;
wire _02736_;
wire _02737_;
wire _02738_;
wire _02739_;
wire _02740_;
wire _02741_;
wire _02742_;
wire _02743_;
wire _02744_;
wire _02745_;
wire _02746_;
wire _02747_;
wire _02748_;
wire _02749_;
wire _02750_;
wire _02751_;
wire _02752_;
wire _02753_;
wire _02754_;
wire _02755_;
wire _02756_;
wire _02757_;
wire _02758_;
wire _02759_;
wire _02760_;
wire _02761_;
wire _02762_;
wire _02763_;
wire _02764_;
wire _02765_;
wire _02766_;
wire _02767_;
wire _02768_;
wire _02769_;
wire _02770_;
wire _02771_;
wire _02772_;
wire _02773_;
wire _02774_;
wire _02775_;
wire _02776_;
wire _02777_;
wire _02778_;
wire _02779_;
wire _02780_;
wire _02781_;
wire _02782_;
wire _02783_;
wire _02784_;
wire _02785_;
wire _02786_;
wire _02787_;
wire _02788_;
wire _02789_;
wire _02790_;
wire _02791_;
wire _02792_;
wire _02793_;
wire _02794_;
wire _02795_;
wire _02796_;
wire _02797_;
wire _02798_;
wire _02799_;
wire _02800_;
wire _02801_;
wire _02802_;
wire _02803_;
wire _02804_;
wire _02805_;
wire _02806_;
wire _02807_;
wire _02808_;
wire _02809_;
wire _02810_;
wire _02811_;
wire _02812_;
wire _02813_;
wire _02814_;
wire _02815_;
wire _02816_;
wire _02817_;
wire _02818_;
wire _02819_;
wire _02820_;
wire _02821_;
wire _02822_;
wire _02823_;
wire _02824_;
wire _02825_;
wire _02826_;
wire _02827_;
wire _02828_;
wire _02829_;
wire _02830_;
wire _02831_;
wire _02832_;
wire _02833_;
wire _02834_;
wire _02835_;
wire _02836_;
wire _02837_;
wire _02838_;
wire _02839_;
wire _02840_;
wire _02841_;
wire _02842_;
wire _02843_;
wire _02844_;
wire _02845_;
wire _02846_;
wire _02847_;
wire _02848_;
wire _02849_;
wire _02850_;
wire _02851_;
wire _02852_;
wire _02853_;
wire _02854_;
wire _02855_;
wire _02856_;
wire _02857_;
wire _02858_;
wire _02859_;
wire _02860_;
wire _02861_;
wire _02862_;
wire _02863_;
wire _02864_;
wire _02865_;
wire _02866_;
wire _02867_;
wire _02868_;
wire _02869_;
wire _02870_;
wire _02871_;
wire _02872_;
wire _02873_;
wire _02874_;
wire _02875_;
wire _02876_;
wire _02877_;
wire _02878_;
wire _02879_;
wire _02880_;
wire _02881_;
wire _02882_;
wire _02883_;
wire _02884_;
wire _02885_;
wire _02886_;
wire _02887_;
wire _02888_;
wire _02889_;
wire _02890_;
wire _02891_;
wire _02892_;
wire _02893_;
wire _02894_;
wire _02895_;
wire _02896_;
wire _02897_;
wire _02898_;
wire _02899_;
wire _02900_;
wire _02901_;
wire _02902_;
wire _02903_;
wire _02904_;
wire _02905_;
wire _02906_;
wire _02907_;
wire _02908_;
wire _02909_;
wire _02910_;
wire _02911_;
wire _02912_;
wire _02913_;
wire _02914_;
wire _02915_;
wire _02916_;
wire _02917_;
wire _02918_;
wire _02919_;
wire _02920_;
wire _02921_;
wire _02922_;
wire _02923_;
wire _02924_;
wire _02925_;
wire _02926_;
wire _02927_;
wire _02928_;
wire _02929_;
wire _02930_;
wire _02931_;
wire _02932_;
wire _02933_;
wire _02934_;
wire _02935_;
wire _02936_;
wire _02937_;
wire _02938_;
wire _02939_;
wire _02940_;
wire _02941_;
wire _02942_;
wire _02943_;
wire _02944_;
wire _02945_;
wire _02946_;
wire _02947_;
wire _02948_;
wire _02949_;
wire _02950_;
wire _02951_;
wire _02952_;
wire _02953_;
wire _02954_;
wire _02955_;
wire _02956_;
wire _02957_;
wire _02958_;
wire _02959_;
wire _02960_;
wire _02961_;
wire _02962_;
wire _02963_;
wire _02964_;
wire _02965_;
wire _02966_;
wire _02967_;
wire _02968_;
wire _02969_;
wire _02970_;
wire _02971_;
wire _02972_;
wire _02973_;
wire _02974_;
wire _02975_;
wire _02976_;
wire _02977_;
wire _02978_;
wire _02979_;
wire _02980_;
wire _02981_;
wire _02982_;
wire _02983_;
wire _02984_;
wire _02985_;
wire _02986_;
wire _02987_;
wire _02988_;
wire _02989_;
wire _02990_;
wire _02991_;
wire _02992_;
wire _02993_;
wire _02994_;
wire _02995_;
wire _02996_;
wire _02997_;
wire _02998_;
wire _02999_;
wire _03000_;
wire _03001_;
wire _03002_;
wire _03003_;
wire _03004_;
wire _03005_;
wire _03006_;
wire _03007_;
wire _03008_;
wire _03009_;
wire _03010_;
wire _03011_;
wire _03012_;
wire _03013_;
wire _03014_;
wire _03015_;
wire _03016_;
wire _03017_;
wire _03018_;
wire _03019_;
wire _03020_;
wire _03021_;
wire _03022_;
wire _03023_;
wire _03024_;
wire _03025_;
wire _03026_;
wire _03027_;
wire _03028_;
wire _03029_;
wire _03030_;
wire _03031_;
wire _03032_;
wire _03033_;
wire _03034_;
wire _03035_;
wire _03036_;
wire _03037_;
wire _03038_;
wire _03039_;
wire _03040_;
wire _03041_;
wire _03042_;
wire _03043_;
wire _03044_;
wire _03045_;
wire _03046_;
wire _03047_;
wire _03048_;
wire _03049_;
wire _03050_;
wire _03051_;
wire _03052_;
wire _03053_;
wire _03054_;
wire _03055_;
wire _03056_;
wire _03057_;
wire _03058_;
wire _03059_;
wire _03060_;
wire _03061_;
wire _03062_;
wire _03063_;
wire _03064_;
wire _03065_;
wire _03066_;
wire _03067_;
wire _03068_;
wire _03069_;
wire _03070_;
wire _03071_;
wire _03072_;
wire _03073_;
wire _03074_;
wire _03075_;
wire _03076_;
wire _03077_;
wire _03078_;
wire _03079_;
wire _03080_;
wire _03081_;
wire _03082_;
wire _03083_;
wire _03084_;
wire _03085_;
wire _03086_;
wire _03087_;
wire _03088_;
wire _03089_;
wire _03090_;
wire _03091_;
wire _03092_;
wire _03093_;
wire _03094_;
wire _03095_;
wire _03096_;
wire _03097_;
wire _03098_;
wire _03099_;
wire _03100_;
wire _03101_;
wire _03102_;
wire _03103_;
wire _03104_;
wire _03105_;
wire _03106_;
wire _03107_;
wire _03108_;
wire _03109_;
wire _03110_;
wire _03111_;
wire _03112_;
wire _03113_;
wire _03114_;
wire _03115_;
wire _03116_;
wire _03117_;
wire _03118_;
wire _03119_;
wire _03120_;
wire _03121_;
wire _03122_;
wire _03123_;
wire _03124_;
wire _03125_;
wire _03126_;
wire _03127_;
wire _03128_;
wire _03129_;
wire _03130_;
wire _03131_;
wire _03132_;
wire _03133_;
wire _03134_;
wire _03135_;
wire _03136_;
wire _03137_;
wire _03138_;
wire _03139_;
wire _03140_;
wire _03141_;
wire _03142_;
wire _03143_;
wire _03144_;
wire _03145_;
wire _03146_;
wire _03147_;
wire _03148_;
wire _03149_;
wire _03150_;
wire _03151_;
wire _03152_;
wire _03153_;
wire _03154_;
wire _03155_;
wire _03156_;
wire _03157_;
wire _03158_;
wire _03159_;
wire _03160_;
wire _03161_;
wire _03162_;
wire _03163_;
wire _03164_;
wire _03165_;
wire _03166_;
wire _03167_;
wire _03168_;
wire _03169_;
wire _03170_;
wire _03171_;
wire _03172_;
wire _03173_;
wire _03174_;
wire _03175_;
wire _03176_;
wire _03177_;
wire _03178_;
wire _03179_;
wire _03180_;
wire _03181_;
wire _03182_;
wire _03183_;
wire _03184_;
wire _03185_;
wire _03186_;
wire _03187_;
wire _03188_;
wire _03189_;
wire _03190_;
wire _03191_;
wire _03192_;
wire _03193_;
wire _03194_;
wire _03195_;
wire _03196_;
wire _03197_;
wire _03198_;
wire _03199_;
wire _03200_;
wire _03201_;
wire _03202_;
wire _03203_;
wire _03204_;
wire _03205_;
wire _03206_;
wire _03207_;
wire _03208_;
wire _03209_;
wire _03210_;
wire _03211_;
wire _03212_;
wire _03213_;
wire _03214_;
wire _03215_;
wire _03216_;
wire _03217_;
wire _03218_;
wire _03219_;
wire _03220_;
wire _03221_;
wire _03222_;
wire _03223_;
wire _03224_;
wire _03225_;
wire _03226_;
wire _03227_;
wire _03228_;
wire _03229_;
wire _03230_;
wire _03231_;
wire _03232_;
wire _03233_;
wire _03234_;
wire _03235_;
wire _03236_;
wire _03237_;
wire _03238_;
wire _03239_;
wire _03240_;
wire _03241_;
wire _03242_;
wire _03243_;
wire _03244_;
wire _03245_;
wire _03246_;
wire _03247_;
wire _03248_;
wire _03249_;
wire _03250_;
wire _03251_;
wire _03252_;
wire _03253_;
wire _03254_;
wire _03255_;
wire _03256_;
wire _03257_;
wire _03258_;
wire _03259_;
wire _03260_;
wire _03261_;
wire _03262_;
wire _03263_;
wire _03264_;
wire _03265_;
wire _03266_;
wire _03267_;
wire _03268_;
wire _03269_;
wire _03270_;
wire _03271_;
wire _03272_;
wire _03273_;
wire _03274_;
wire _03275_;
wire _03276_;
wire _03277_;
wire _03278_;
wire _03279_;
wire _03280_;
wire _03281_;
wire _03282_;
wire _03283_;
wire _03284_;
wire _03285_;
wire _03286_;
wire _03287_;
wire _03288_;
wire _03289_;
wire _03290_;
wire _03291_;
wire _03292_;
wire _03293_;
wire _03294_;
wire _03295_;
wire _03296_;
wire _03297_;
wire _03298_;
wire _03299_;
wire _03300_;
wire _03301_;
wire _03302_;
wire _03303_;
wire _03304_;
wire _03305_;
wire _03306_;
wire _03307_;
wire _03308_;
wire _03309_;
wire _03310_;
wire _03311_;
wire _03312_;
wire _03313_;
wire _03314_;
wire _03315_;
wire _03316_;
wire _03317_;
wire _03318_;
wire _03319_;
wire _03320_;
wire _03321_;
wire _03322_;
wire _03323_;
wire _03324_;
wire _03325_;
wire _03326_;
wire _03327_;
wire _03328_;
wire _03329_;
wire _03330_;
wire _03331_;
wire _03332_;
wire _03333_;
wire _03334_;
wire _03335_;
wire _03336_;
wire _03337_;
wire _03338_;
wire _03339_;
wire _03340_;
wire _03341_;
wire _03342_;
wire _03343_;
wire _03344_;
wire _03345_;
wire _03346_;
wire _03347_;
wire _03348_;
wire _03349_;
wire _03350_;
wire _03351_;
wire _03352_;
wire _03353_;
wire _03354_;
wire _03355_;
wire _03356_;
wire _03357_;
wire _03358_;
wire _03359_;
wire _03360_;
wire _03361_;
wire _03362_;
wire _03363_;
wire _03364_;
wire _03365_;
wire _03366_;
wire _03367_;
wire _03368_;
wire _03369_;
wire _03370_;
wire _03371_;
wire _03372_;
wire _03373_;
wire _03374_;
wire _03375_;
wire _03376_;
wire _03377_;
wire _03378_;
wire _03379_;
wire _03380_;
wire _03381_;
wire _03382_;
wire _03383_;
wire _03384_;
wire _03385_;
wire _03386_;
wire _03387_;
wire _03388_;
wire _03389_;
wire _03390_;
wire _03391_;
wire _03392_;
wire _03393_;
wire _03394_;
wire _03395_;
wire _03396_;
wire _03397_;
wire _03398_;
wire _03399_;
wire _03400_;
wire _03401_;
wire _03402_;
wire _03403_;
wire _03404_;
wire _03405_;
wire _03406_;
wire _03407_;
wire _03408_;
wire _03409_;
wire _03410_;
wire _03411_;
wire _03412_;
wire _03413_;
wire _03414_;
wire _03415_;
wire _03416_;
wire _03417_;
wire _03418_;
wire _03419_;
wire _03420_;
wire _03421_;
wire _03422_;
wire _03423_;
wire _03424_;
wire _03425_;
wire _03426_;
wire _03427_;
wire _03428_;
wire _03429_;
wire _03430_;
wire _03431_;
wire _03432_;
wire _03433_;
wire _03434_;
wire _03435_;
wire _03436_;
wire _03437_;
wire _03438_;
wire _03439_;
wire _03440_;
wire _03441_;
wire _03442_;
wire _03443_;
wire _03444_;
wire _03445_;
wire _03446_;
wire _03447_;
wire _03448_;
wire _03449_;
wire _03450_;
wire _03451_;
wire _03452_;
wire _03453_;
wire _03454_;
wire _03455_;
wire _03456_;
wire _03457_;
wire _03458_;
wire _03459_;
wire _03460_;
wire _03461_;
wire _03462_;
wire _03463_;
wire _03464_;
wire _03465_;
wire _03466_;
wire _03467_;
wire _03468_;
wire _03469_;
wire _03470_;
wire _03471_;
wire _03472_;
wire _03473_;
wire _03474_;
wire _03475_;
wire _03476_;
wire _03477_;
wire _03478_;
wire _03479_;
wire _03480_;
wire _03481_;
wire _03482_;
wire _03483_;
wire _03484_;
wire _03485_;
wire _03486_;
wire _03487_;
wire _03488_;
wire _03489_;
wire _03490_;
wire _03491_;
wire _03492_;
wire _03493_;
wire _03494_;
wire _03495_;
wire _03496_;
wire _03497_;
wire _03498_;
wire _03499_;
wire _03500_;
wire _03501_;
wire _03502_;
wire _03503_;
wire _03504_;
wire _03505_;
wire _03506_;
wire _03507_;
wire _03508_;
wire _03509_;
wire _03510_;
wire _03511_;
wire _03512_;
wire _03513_;
wire _03514_;
wire _03515_;
wire _03516_;
wire _03517_;
wire _03518_;
wire _03519_;
wire _03520_;
wire _03521_;
wire _03522_;
wire _03523_;
wire _03524_;
wire _03525_;
wire _03526_;
wire _03527_;
wire _03528_;
wire _03529_;
wire _03530_;
wire _03531_;
wire _03532_;
wire _03533_;
wire _03534_;
wire _03535_;
wire _03536_;
wire _03537_;
wire _03538_;
wire _03539_;
wire _03540_;
wire _03541_;
wire _03542_;
wire _03543_;
wire _03544_;
wire _03545_;
wire _03546_;
wire _03547_;
wire _03548_;
wire _03549_;
wire _03550_;
wire _03551_;
wire _03552_;
wire _03553_;
wire _03554_;
wire _03555_;
wire _03556_;
wire _03557_;
wire _03558_;
wire _03559_;
wire _03560_;
wire _03561_;
wire _03562_;
wire _03563_;
wire _03564_;
wire _03565_;
wire _03566_;
wire _03567_;
wire _03568_;
wire _03569_;
wire _03570_;
wire _03571_;
wire _03572_;
wire _03573_;
wire _03574_;
wire _03575_;
wire _03576_;
wire _03577_;
wire _03578_;
wire _03579_;
wire _03580_;
wire _03581_;
wire _03582_;
wire _03583_;
wire _03584_;
wire _03585_;
wire _03586_;
wire _03587_;
wire _03588_;
wire _03589_;
wire _03590_;
wire _03591_;
wire _03592_;
wire _03593_;
wire _03594_;
wire _03595_;
wire _03596_;
wire _03597_;
wire _03598_;
wire _03599_;
wire _03600_;
wire _03601_;
wire _03602_;
wire _03603_;
wire _03604_;
wire _03605_;
wire _03606_;
wire _03607_;
wire _03608_;
wire _03609_;
wire _03610_;
wire _03611_;
wire _03612_;
wire _03613_;
wire _03614_;
wire _03615_;
wire _03616_;
wire _03617_;
wire _03618_;
wire _03619_;
wire _03620_;
wire _03621_;
wire _03622_;
wire _03623_;
wire _03624_;
wire _03625_;
wire _03626_;
wire _03627_;
wire _03628_;
wire _03629_;
wire _03630_;
wire _03631_;
wire _03632_;
wire _03633_;
wire _03634_;
wire _03635_;
wire _03636_;
wire _03637_;
wire _03638_;
wire _03639_;
wire _03640_;
wire _03641_;
wire _03642_;
wire _03643_;
wire _03644_;
wire _03645_;
wire _03646_;
wire _03647_;
wire _03648_;
wire _03649_;
wire _03650_;
wire _03651_;
wire _03652_;
wire _03653_;
wire _03654_;
wire _03655_;
wire _03656_;
wire _03657_;
wire _03658_;
wire _03659_;
wire _03660_;
wire _03661_;
wire _03662_;
wire _03663_;
wire _03664_;
wire _03665_;
wire _03666_;
wire _03667_;
wire _03668_;
wire _03669_;
wire _03670_;
wire _03671_;
wire _03672_;
wire _03673_;
wire _03674_;
wire _03675_;
wire _03676_;
wire _03677_;
wire _03678_;
wire _03679_;
wire _03680_;
wire _03681_;
wire _03682_;
wire _03683_;
wire _03684_;
wire _03685_;
wire _03686_;
wire _03687_;
wire _03688_;
wire _03689_;
wire _03690_;
wire _03691_;
wire _03692_;
wire _03693_;
wire _03694_;
wire _03695_;
wire _03696_;
wire _03697_;
wire _03698_;
wire _03699_;
wire _03700_;
wire _03701_;
wire _03702_;
wire _03703_;
wire _03704_;
wire _03705_;
wire _03706_;
wire _03707_;
wire _03708_;
wire _03709_;
wire _03710_;
wire _03711_;
wire _03712_;
wire _03713_;
wire _03714_;
wire _03715_;
wire _03716_;
wire _03717_;
wire _03718_;
wire _03719_;
wire _03720_;
wire _03721_;
wire _03722_;
wire _03723_;
wire _03724_;
wire _03725_;
wire _03726_;
wire _03727_;
wire _03728_;
wire _03729_;
wire _03730_;
wire _03731_;
wire _03732_;
wire _03733_;
wire _03734_;
wire _03735_;
wire _03736_;
wire _03737_;
wire _03738_;
wire _03739_;
wire _03740_;
wire _03741_;
wire _03742_;
wire _03743_;
wire _03744_;
wire _03745_;
wire _03746_;
wire _03747_;
wire _03748_;
wire _03749_;
wire _03750_;
wire _03751_;
wire _03752_;
wire _03753_;
wire _03754_;
wire _03755_;
wire _03756_;
wire _03757_;
wire _03758_;
wire _03759_;
wire _03760_;
wire _03761_;
wire _03762_;
wire _03763_;
wire _03764_;
wire _03765_;
wire _03766_;
wire _03767_;
wire _03768_;
wire _03769_;
wire _03770_;
wire _03771_;
wire _03772_;
wire _03773_;
wire _03774_;
wire _03775_;
wire _03776_;
wire _03777_;
wire _03778_;
wire _03779_;
wire _03780_;
wire _03781_;
wire _03782_;
wire _03783_;
wire _03784_;
wire _03785_;
wire _03786_;
wire _03787_;
wire _03788_;
wire _03789_;
wire _03790_;
wire _03791_;
wire _03792_;
wire _03793_;
wire _03794_;
wire _03795_;
wire _03796_;
wire _03797_;
wire _03798_;
wire _03799_;
wire _03800_;
wire _03801_;
wire _03802_;
wire _03803_;
wire _03804_;
wire _03805_;
wire _03806_;
wire _03807_;
wire _03808_;
wire _03809_;
wire _03810_;
wire _03811_;
wire _03812_;
wire _03813_;
wire _03814_;
wire _03815_;
wire _03816_;
wire _03817_;
wire _03818_;
wire _03819_;
wire _03820_;
wire _03821_;
wire _03822_;
wire _03823_;
wire _03824_;
wire _03825_;
wire _03826_;
wire _03827_;
wire _03828_;
wire _03829_;
wire _03830_;
wire _03831_;
wire _03832_;
wire _03833_;
wire _03834_;
wire _03835_;
wire _03836_;
wire _03837_;
wire _03838_;
wire _03839_;
wire _03840_;
wire _03841_;
wire _03842_;
wire _03843_;
wire _03844_;
wire _03845_;
wire _03846_;
wire _03847_;
wire _03848_;
wire _03849_;
wire _03850_;
wire _03851_;
wire _03852_;
wire _03853_;
wire _03854_;
wire _03855_;
wire _03856_;
wire _03857_;
wire _03858_;
wire _03859_;
wire _03860_;
wire _03861_;
wire _03862_;
wire _03863_;
wire _03864_;
wire _03865_;
wire _03866_;
wire _03867_;
wire _03868_;
wire _03869_;
wire _03870_;
wire _03871_;
wire _03872_;
wire _03873_;
wire _03874_;
wire _03875_;
wire _03876_;
wire _03877_;
wire _03878_;
wire _03879_;
wire _03880_;
wire _03881_;
wire _03882_;
wire _03883_;
wire _03884_;
wire _03885_;
wire _03886_;
wire _03887_;
wire _03888_;
wire _03889_;
wire _03890_;
wire _03891_;
wire _03892_;
wire _03893_;
wire _03894_;
wire _03895_;
wire _03896_;
wire _03897_;
wire _03898_;
wire _03899_;
wire _03900_;
wire _03901_;
wire _03902_;
wire _03903_;
wire _03904_;
wire _03905_;
wire _03906_;
wire _03907_;
wire _03908_;
wire _03909_;
wire _03910_;
wire _03911_;
wire _03912_;
wire _03913_;
wire _03914_;
wire _03915_;
wire _03916_;
wire _03917_;
wire _03918_;
wire _03919_;
wire _03920_;
wire _03921_;
wire _03922_;
wire _03923_;
wire _03924_;
wire _03925_;
wire _03926_;
wire _03927_;
wire _03928_;
wire _03929_;
wire _03930_;
wire _03931_;
wire _03932_;
wire _03933_;
wire _03934_;
wire _03935_;
wire _03936_;
wire _03937_;
wire _03938_;
wire _03939_;
wire _03940_;
wire _03941_;
wire _03942_;
wire _03943_;
wire _03944_;
wire _03945_;
wire _03946_;
wire _03947_;
wire _03948_;
wire _03949_;
wire _03950_;
wire _03951_;
wire _03952_;
wire _03953_;
wire _03954_;
wire _03955_;
wire _03956_;
wire _03957_;
wire _03958_;
wire _03959_;
wire _03960_;
wire _03961_;
wire _03962_;
wire _03963_;
wire _03964_;
wire _03965_;
wire _03966_;
wire _03967_;
wire _03968_;
wire _03969_;
wire _03970_;
wire _03971_;
wire _03972_;
wire _03973_;
wire _03974_;
wire _03975_;
wire _03976_;
wire _03977_;
wire _03978_;
wire _03979_;
wire _03980_;
wire _03981_;
wire _03982_;
wire _03983_;
wire _03984_;
wire _03985_;
wire _03986_;
wire _03987_;
wire _03988_;
wire _03989_;
wire _03990_;
wire _03991_;
wire _03992_;
wire _03993_;
wire _03994_;
wire _03995_;
wire _03996_;
wire _03997_;
wire _03998_;
wire _03999_;
wire _04000_;
wire _04001_;
wire _04002_;
wire _04003_;
wire _04004_;
wire _04005_;
wire _04006_;
wire _04007_;
wire _04008_;
wire _04009_;
wire _04010_;
wire _04011_;
wire _04012_;
wire _04013_;
wire _04014_;
wire _04015_;
wire _04016_;
wire _04017_;
wire _04018_;
wire _04019_;
wire _04020_;
wire _04021_;
wire _04022_;
wire _04023_;
wire _04024_;
wire _04025_;
wire _04026_;
wire _04027_;
wire _04028_;
wire _04029_;
wire _04030_;
wire _04031_;
wire _04032_;
wire _04033_;
wire _04034_;
wire _04035_;
wire _04036_;
wire _04037_;
wire _04038_;
wire _04039_;
wire _04040_;
wire _04041_;
wire _04042_;
wire _04043_;
wire _04044_;
wire _04045_;
wire _04046_;
wire _04047_;
wire _04048_;
wire _04049_;
wire _04050_;
wire _04051_;
wire _04052_;
wire _04053_;
wire _04054_;
wire _04055_;
wire _04056_;
wire _04057_;
wire _04058_;
wire _04059_;
wire _04060_;
wire _04061_;
wire _04062_;
wire _04063_;
wire _04064_;
wire _04065_;
wire _04066_;
wire _04067_;
wire _04068_;
wire _04069_;
wire _04070_;
wire _04071_;
wire _04072_;
wire _04073_;
wire _04074_;
wire _04075_;
wire _04076_;
wire _04077_;
wire _04078_;
wire _04079_;
wire _04080_;
wire _04081_;
wire _04082_;
wire _04083_;
wire _04084_;
wire _04085_;
wire _04086_;
wire _04087_;
wire _04088_;
wire _04089_;
wire _04090_;
wire _04091_;
wire _04092_;
wire _04093_;
wire _04094_;
wire _04095_;
wire _04096_;
wire _04097_;
wire _04098_;
wire _04099_;
wire _04100_;
wire _04101_;
wire _04102_;
wire _04103_;
wire _04104_;
wire _04105_;
wire _04106_;
wire _04107_;
wire _04108_;
wire _04109_;
wire _04110_;
wire _04111_;
wire _04112_;
wire _04113_;
wire _04114_;
wire _04115_;
wire _04116_;
wire _04117_;
wire _04118_;
wire _04119_;
wire _04120_;
wire _04121_;
wire _04122_;
wire _04123_;
wire _04124_;
wire _04125_;
wire _04126_;
wire _04127_;
wire _04128_;
wire _04129_;
wire _04130_;
wire _04131_;
wire _04132_;
wire _04133_;
wire _04134_;
wire _04135_;
wire _04136_;
wire _04137_;
wire _04138_;
wire _04139_;
wire _04140_;
wire _04141_;
wire _04142_;
wire _04143_;
wire _04144_;
wire _04145_;
wire _04146_;
wire _04147_;
wire _04148_;
wire _04149_;
wire _04150_;
wire _04151_;
wire _04152_;
wire _04153_;
wire _04154_;
wire _04155_;
wire _04156_;
wire _04157_;
wire _04158_;
wire _04159_;
wire _04160_;
wire _04161_;
wire _04162_;
wire _04163_;
wire _04164_;
wire _04165_;
wire _04166_;
wire _04167_;
wire _04168_;
wire _04169_;
wire _04170_;
wire _04171_;
wire _04172_;
wire _04173_;
wire _04174_;
wire _04175_;
wire _04176_;
wire _04177_;
wire _04178_;
wire _04179_;
wire _04180_;
wire _04181_;
wire _04182_;
wire _04183_;
wire _04184_;
wire _04185_;
wire _04186_;
wire _04187_;
wire _04188_;
wire _04189_;
wire _04190_;
wire _04191_;
wire _04192_;
wire _04193_;
wire _04194_;
wire _04195_;
wire _04196_;
wire _04197_;
wire _04198_;
wire _04199_;
wire _04200_;
wire _04201_;
wire _04202_;
wire _04203_;
wire _04204_;
wire _04205_;
wire _04206_;
wire _04207_;
wire _04208_;
wire _04209_;
wire _04210_;
wire _04211_;
wire _04212_;
wire _04213_;
wire _04214_;
wire _04215_;
wire _04216_;
wire _04217_;
wire _04218_;
wire _04219_;
wire _04220_;
wire _04221_;
wire _04222_;
wire _04223_;
wire _04224_;
wire _04225_;
wire _04226_;
wire _04227_;
wire _04228_;
wire _04229_;
wire _04230_;
wire _04231_;
wire _04232_;
wire _04233_;
wire _04234_;
wire _04235_;
wire _04236_;
wire _04237_;
wire _04238_;
wire _04239_;
wire _04240_;
wire _04241_;
wire _04242_;
wire _04243_;
wire _04244_;
wire _04245_;
wire _04246_;
wire _04247_;
wire _04248_;
wire _04249_;
wire _04250_;
wire _04251_;
wire _04252_;
wire _04253_;
wire _04254_;
wire _04255_;
wire _04256_;
wire _04257_;
wire _04258_;
wire _04259_;
wire _04260_;
wire _04261_;
wire _04262_;
wire _04263_;
wire _04264_;
wire _04265_;
wire _04266_;
wire _04267_;
wire _04268_;
wire _04269_;
wire _04270_;
wire _04271_;
wire _04272_;
wire _04273_;
wire _04274_;
wire _04275_;
wire _04276_;
wire _04277_;
wire _04278_;
wire _04279_;
wire _04280_;
wire _04281_;
wire _04282_;
wire _04283_;
wire _04284_;
wire _04285_;
wire _04286_;
wire _04287_;
wire _04288_;
wire _04289_;
wire _04290_;
wire _04291_;
wire _04292_;
wire _04293_;
wire _04294_;
wire _04295_;
wire _04296_;
wire _04297_;
wire _04298_;
wire _04299_;
wire _04300_;
wire _04301_;
wire _04302_;
wire _04303_;
wire _04304_;
wire _04305_;
wire _04306_;
wire _04307_;
wire _04308_;
wire _04309_;
wire _04310_;
wire _04311_;
wire _04312_;
wire _04313_;
wire _04314_;
wire _04315_;
wire _04316_;
wire _04317_;
wire _04318_;
wire _04319_;
wire _04320_;
wire _04321_;
wire _04322_;
wire _04323_;
wire _04324_;
wire _04325_;
wire _04326_;
wire _04327_;
wire _04328_;
wire _04329_;
wire _04330_;
wire _04331_;
wire _04332_;
wire _04333_;
wire _04334_;
wire _04335_;
wire _04336_;
wire _04337_;
wire _04338_;
wire _04339_;
wire _04340_;
wire _04341_;
wire _04342_;
wire _04343_;
wire _04344_;
wire _04345_;
wire _04346_;
wire _04347_;
wire _04348_;
wire _04349_;
wire _04350_;
wire _04351_;
wire _04352_;
wire _04353_;
wire _04354_;
wire _04355_;
wire _04356_;
wire _04357_;
wire _04358_;
wire _04359_;
wire _04360_;
wire _04361_;
wire _04362_;
wire _04363_;
wire _04364_;
wire _04365_;
wire _04366_;
wire _04367_;
wire _04368_;
wire _04369_;
wire _04370_;
wire _04371_;
wire _04372_;
wire _04373_;
wire _04374_;
wire _04375_;
wire _04376_;
wire _04377_;
wire _04378_;
wire _04379_;
wire _04380_;
wire _04381_;
wire _04382_;
wire _04383_;
wire _04384_;
wire _04385_;
wire _04386_;
wire _04387_;
wire _04388_;
wire _04389_;
wire _04390_;
wire _04391_;
wire _04392_;
wire _04393_;
wire _04394_;
wire _04395_;
wire _04396_;
wire _04397_;
wire _04398_;
wire _04399_;
wire _04400_;
wire _04401_;
wire _04402_;
wire _04403_;
wire _04404_;
wire _04405_;
wire _04406_;
wire _04407_;
wire _04408_;
wire _04409_;
wire _04410_;
wire _04411_;
wire _04412_;
wire _04413_;
wire _04414_;
wire _04415_;
wire _04416_;
wire _04417_;
wire _04418_;
wire _04419_;
wire _04420_;
wire _04421_;
wire _04422_;
wire _04423_;
wire _04424_;
wire _04425_;
wire _04426_;
wire _04427_;
wire _04428_;
wire _04429_;
wire _04430_;
wire _04431_;
wire _04432_;
wire _04433_;
wire _04434_;
wire _04435_;
wire _04436_;
wire _04437_;
wire _04438_;
wire _04439_;
wire _04440_;
wire _04441_;
wire _04442_;
wire _04443_;
wire _04444_;
wire _04445_;
wire _04446_;
wire _04447_;
wire _04448_;
wire _04449_;
wire _04450_;
wire _04451_;
wire _04452_;
wire _04453_;
wire _04454_;
wire _04455_;
wire _04456_;
wire _04457_;
wire _04458_;
wire _04459_;
wire _04460_;
wire _04461_;
wire _04462_;
wire _04463_;
wire _04464_;
wire _04465_;
wire _04466_;
wire _04467_;
wire _04468_;
wire _04469_;
wire _04470_;
wire _04471_;
wire _04472_;
wire _04473_;
wire _04474_;
wire _04475_;
wire _04476_;
wire _04477_;
wire _04478_;
wire _04479_;
wire _04480_;
wire _04481_;
wire _04482_;
wire _04483_;
wire _04484_;
wire _04485_;
wire _04486_;
wire _04487_;
wire _04488_;
wire _04489_;
wire _04490_;
wire _04491_;
wire _04492_;
wire _04493_;
wire _04494_;
wire _04495_;
wire _04496_;
wire _04497_;
wire _04498_;
wire _04499_;
wire _04500_;
wire _04501_;
wire _04502_;
wire _04503_;
wire _04504_;
wire _04505_;
wire _04506_;
wire _04507_;
wire _04508_;
wire _04509_;
wire _04510_;
wire _04511_;
wire _04512_;
wire _04513_;
wire _04514_;
wire _04515_;
wire _04516_;
wire _04517_;
wire _04518_;
wire _04519_;
wire _04520_;
wire _04521_;
wire _04522_;
wire _04523_;
wire _04524_;
wire _04525_;
wire _04526_;
wire _04527_;
wire _04528_;
wire _04529_;
wire _04530_;
wire _04531_;
wire _04532_;
wire _04533_;
wire _04534_;
wire _04535_;
wire _04536_;
wire _04537_;
wire _04538_;
wire _04539_;
wire _04540_;
wire _04541_;
wire _04542_;
wire _04543_;
wire _04544_;
wire _04545_;
wire _04546_;
wire _04547_;
wire _04548_;
wire _04549_;
wire _04550_;
wire _04551_;
wire _04552_;
wire _04553_;
wire _04554_;
wire _04555_;
wire _04556_;
wire _04557_;
wire _04558_;
wire _04559_;
wire _04560_;
wire _04561_;
wire _04562_;
wire _04563_;
wire _04564_;
wire _04565_;
wire _04566_;
wire _04567_;
wire _04568_;
wire _04569_;
wire _04570_;
wire _04571_;
wire _04572_;
wire _04573_;
wire _04574_;
wire _04575_;
wire _04576_;
wire _04577_;
wire _04578_;
wire _04579_;
wire _04580_;
wire _04581_;
wire _04582_;
wire _04583_;
wire _04584_;
wire _04585_;
wire _04586_;
wire _04587_;
wire _04588_;
wire _04589_;
wire _04590_;
wire _04591_;
wire _04592_;
wire _04593_;
wire _04594_;
wire _04595_;
wire _04596_;
wire _04597_;
wire _04598_;
wire _04599_;
wire _04600_;
wire _04601_;
wire _04602_;
wire _04603_;
wire _04604_;
wire _04605_;
wire _04606_;
wire _04607_;
wire _04608_;
wire _04609_;
wire _04610_;
wire _04611_;
wire _04612_;
wire _04613_;
wire _04614_;
wire _04615_;
wire _04616_;
wire _04617_;
wire _04618_;
wire _04619_;
wire _04620_;
wire _04621_;
wire _04622_;
wire _04623_;
wire _04624_;
wire _04625_;
wire _04626_;
wire _04627_;
wire _04628_;
wire _04629_;
wire _04630_;
wire _04631_;
wire _04632_;
wire _04633_;
wire _04634_;
wire _04635_;
wire _04636_;
wire _04637_;
wire _04638_;
wire _04639_;
wire _04640_;
wire _04641_;
wire _04642_;
wire _04643_;
wire _04644_;
wire _04645_;
wire _04646_;
wire _04647_;
wire _04648_;
wire _04649_;
wire _04650_;
wire _04651_;
wire _04652_;
wire _04653_;
wire _04654_;
wire _04655_;
wire _04656_;
wire _04657_;
wire _04658_;
wire _04659_;
wire _04660_;
wire _04661_;
wire _04662_;
wire _04663_;
wire _04664_;
wire _04665_;
wire _04666_;
wire _04667_;
wire _04668_;
wire _04669_;
wire _04670_;
wire _04671_;
wire _04672_;
wire _04673_;
wire _04674_;
wire _04675_;
wire _04676_;
wire _04677_;
wire _04678_;
wire _04679_;
wire _04680_;
wire _04681_;
wire _04682_;
wire _04683_;
wire _04684_;
wire _04685_;
wire _04686_;
wire _04687_;
wire _04688_;
wire _04689_;
wire _04690_;
wire _04691_;
wire _04692_;
wire _04693_;
wire _04694_;
wire _04695_;
wire _04696_;
wire _04697_;
wire _04698_;
wire _04699_;
wire _04700_;
wire _04701_;
wire _04702_;
wire _04703_;
wire _04704_;
wire _04705_;
wire _04706_;
wire _04707_;
wire _04708_;
wire _04709_;
wire _04710_;
wire _04711_;
wire _04712_;
wire _04713_;
wire _04714_;
wire _04715_;
wire _04716_;
wire _04717_;
wire _04718_;
wire _04719_;
wire _04720_;
wire _04721_;
wire _04722_;
wire _04723_;
wire _04724_;
wire _04725_;
wire _04726_;
wire _04727_;
wire _04728_;
wire _04729_;
wire _04730_;
wire _04731_;
wire _04732_;
wire _04733_;
wire _04734_;
wire _04735_;
wire _04736_;
wire _04737_;
wire _04738_;
wire _04739_;
wire _04740_;
wire _04741_;
wire _04742_;
wire _04743_;
wire _04744_;
wire _04745_;
wire _04746_;
wire _04747_;
wire _04748_;
wire _04749_;
wire _04750_;
wire _04751_;
wire _04752_;
wire _04753_;
wire _04754_;
wire _04755_;
wire _04756_;
wire _04757_;
wire _04758_;
wire _04759_;
wire _04760_;
wire _04761_;
wire _04762_;
wire _04763_;
wire _04764_;
wire _04765_;
wire _04766_;
wire _04767_;
wire _04768_;
wire _04769_;
wire _04770_;
wire _04771_;
wire _04772_;
wire _04773_;
wire _04774_;
wire _04775_;
wire _04776_;
wire _04777_;
wire _04778_;
wire _04779_;
wire _04780_;
wire _04781_;
wire _04782_;
wire _04783_;
wire _04784_;
wire _04785_;
wire _04786_;
wire _04787_;
wire _04788_;
wire _04789_;
wire _04790_;
wire _04791_;
wire _04792_;
wire _04793_;
wire _04794_;
wire _04795_;
wire _04796_;
wire _04797_;
wire _04798_;
wire _04799_;
wire _04800_;
wire _04801_;
wire _04802_;
wire _04803_;
wire _04804_;
wire _04805_;
wire _04806_;
wire _04807_;
wire _04808_;
wire _04809_;
wire _04810_;
wire _04811_;
wire _04812_;
wire _04813_;
wire _04814_;
wire _04815_;
wire _04816_;
wire _04817_;
wire _04818_;
wire _04819_;
wire _04820_;
wire _04821_;
wire _04822_;
wire _04823_;
wire _04824_;
wire _04825_;
wire _04826_;
wire _04827_;
wire _04828_;
wire _04829_;
wire _04830_;
wire _04831_;
wire _04832_;
wire _04833_;
wire _04834_;
wire _04835_;
wire _04836_;
wire _04837_;
wire _04838_;
wire _04839_;
wire _04840_;
wire _04841_;
wire _04842_;
wire _04843_;
wire _04844_;
wire _04845_;
wire _04846_;
wire _04847_;
wire _04848_;
wire _04849_;
wire _04850_;
wire _04851_;
wire _04852_;
wire _04853_;
wire _04854_;
wire _04855_;
wire _04856_;
wire _04857_;
wire _04858_;
wire _04859_;
wire _04860_;
wire _04861_;
wire _04862_;
wire _04863_;
wire _04864_;
wire _04865_;
wire _04866_;
wire _04867_;
wire _04868_;
wire _04869_;
wire _04870_;
wire _04871_;
wire _04872_;
wire _04873_;
wire _04874_;
wire _04875_;
wire _04876_;
wire _04877_;
wire _04878_;
wire _04879_;
wire _04880_;
wire _04881_;
wire _04882_;
wire _04883_;
wire _04884_;
wire _04885_;
wire _04886_;
wire _04887_;
wire _04888_;
wire _04889_;
wire _04890_;
wire _04891_;
wire _04892_;
wire _04893_;
wire _04894_;
wire _04895_;
wire _04896_;
wire _04897_;
wire _04898_;
wire _04899_;
wire _04900_;
wire _04901_;
wire _04902_;
wire _04903_;
wire _04904_;
wire _04905_;
wire _04906_;
wire _04907_;
wire _04908_;
wire _04909_;
wire _04910_;
wire _04911_;
wire _04912_;
wire _04913_;
wire _04914_;
wire _04915_;
wire _04916_;
wire _04917_;
wire _04918_;
wire _04919_;
wire _04920_;
wire _04921_;
wire _04922_;
wire _04923_;
wire _04924_;
wire _04925_;
wire _04926_;
wire _04927_;
wire _04928_;
wire _04929_;
wire _04930_;
wire _04931_;
wire _04932_;
wire _04933_;
wire _04934_;
wire _04935_;
wire _04936_;
wire _04937_;
wire _04938_;
wire _04939_;
wire _04940_;
wire _04941_;
wire _04942_;
wire _04943_;
wire _04944_;
wire _04945_;
wire _04946_;
wire _04947_;
wire _04948_;
wire _04949_;
wire _04950_;
wire _04951_;
wire _04952_;
wire _04953_;
wire _04954_;
wire _04955_;
wire _04956_;
wire _04957_;
wire _04958_;
wire _04959_;
wire _04960_;
wire _04961_;
wire _04962_;
wire _04963_;
wire _04964_;
wire _04965_;
wire _04966_;
wire _04967_;
wire _04968_;
wire _04969_;
wire _04970_;
wire _04971_;
wire _04972_;
wire _04973_;
wire _04974_;
wire _04975_;
wire _04976_;
wire _04977_;
wire _04978_;
wire _04979_;
wire _04980_;
wire _04981_;
wire _04982_;
wire _04983_;
wire _04984_;
wire _04985_;
wire _04986_;
wire _04987_;
wire _04988_;
wire _04989_;
wire _04990_;
wire _04991_;
wire _04992_;
wire _04993_;
wire _04994_;
wire _04995_;
wire _04996_;
wire _04997_;
wire _04998_;
wire _04999_;
wire _05000_;
wire _05001_;
wire _05002_;
wire _05003_;
wire _05004_;
wire _05005_;
wire _05006_;
wire _05007_;
wire _05008_;
wire _05009_;
wire _05010_;
wire _05011_;
wire _05012_;
wire _05013_;
wire _05014_;
wire _05015_;
wire _05016_;
wire _05017_;
wire _05018_;
wire _05019_;
wire _05020_;
wire _05021_;
wire _05022_;
wire _05023_;
wire _05024_;
wire _05025_;
wire _05026_;
wire _05027_;
wire _05028_;
wire _05029_;
wire _05030_;
wire _05031_;
wire _05032_;
wire _05033_;
wire _05034_;
wire _05035_;
wire _05036_;
wire _05037_;
wire _05038_;
wire _05039_;
wire _05040_;
wire _05041_;
wire _05042_;
wire _05043_;
wire _05044_;
wire _05045_;
wire _05046_;
wire _05047_;
wire _05048_;
wire _05049_;
wire _05050_;
wire _05051_;
wire _05052_;
wire _05053_;
wire _05054_;
wire _05055_;
wire _05056_;
wire _05057_;
wire _05058_;
wire _05059_;
wire _05060_;
wire _05061_;
wire _05062_;
wire _05063_;
wire _05064_;
wire _05065_;
wire _05066_;
wire _05067_;
wire _05068_;
wire _05069_;
wire _05070_;
wire _05071_;
wire _05072_;
wire _05073_;
wire _05074_;
wire _05075_;
wire _05076_;
wire _05077_;
wire _05078_;
wire _05079_;
wire _05080_;
wire _05081_;
wire _05082_;
wire _05083_;
wire _05084_;
wire _05085_;
wire _05086_;
wire _05087_;
wire _05088_;
wire _05089_;
wire _05090_;
wire _05091_;
wire _05092_;
wire _05093_;
wire _05094_;
wire _05095_;
wire _05096_;
wire _05097_;
wire _05098_;
wire _05099_;
wire _05100_;
wire _05101_;
wire _05102_;
wire _05103_;
wire _05104_;
wire _05105_;
wire _05106_;
wire _05107_;
wire _05108_;
wire _05109_;
wire _05110_;
wire _05111_;
wire _05112_;
wire _05113_;
wire _05114_;
wire _05115_;
wire _05116_;
wire _05117_;
wire _05118_;
wire _05119_;
wire _05120_;
wire _05121_;
wire _05122_;
wire _05123_;
wire _05124_;
wire _05125_;
wire _05126_;
wire _05127_;
wire _05128_;
wire _05129_;
wire _05130_;
wire _05131_;
wire _05132_;
wire _05133_;
wire _05134_;
wire _05135_;
wire _05136_;
wire _05137_;
wire _05138_;
wire _05139_;
wire _05140_;
wire _05141_;
wire _05142_;
wire _05143_;
wire _05144_;
wire _05145_;
wire _05146_;
wire _05147_;
wire _05148_;
wire _05149_;
wire _05150_;
wire _05151_;
wire _05152_;
wire _05153_;
wire _05154_;
wire _05155_;
wire _05156_;
wire _05157_;
wire _05158_;
wire _05159_;
wire _05160_;
wire _05161_;
wire _05162_;
wire _05163_;
wire _05164_;
wire _05165_;
wire _05166_;
wire _05167_;
wire _05168_;
wire _05169_;
wire _05170_;
wire _05171_;
wire _05172_;
wire _05173_;
wire _05174_;
wire _05175_;
wire _05176_;
wire _05177_;
wire _05178_;
wire _05179_;
wire _05180_;
wire _05181_;
wire _05182_;
wire _05183_;
wire _05184_;
wire _05185_;
wire _05186_;
wire _05187_;
wire _05188_;
wire _05189_;
wire _05190_;
wire _05191_;
wire _05192_;
wire _05193_;
wire _05194_;
wire _05195_;
wire _05196_;
wire _05197_;
wire _05198_;
wire _05199_;
wire _05200_;
wire _05201_;
wire _05202_;
wire _05203_;
wire _05204_;
wire _05205_;
wire _05206_;
wire _05207_;
wire _05208_;
wire _05209_;
wire _05210_;
wire _05211_;
wire _05212_;
wire _05213_;
wire _05214_;
wire _05215_;
wire _05216_;
wire _05217_;
wire _05218_;
wire _05219_;
wire _05220_;
wire _05221_;
wire _05222_;
wire _05223_;
wire _05224_;
wire _05225_;
wire _05226_;
wire _05227_;
wire _05228_;
wire _05229_;
wire _05230_;
wire _05231_;
wire _05232_;
wire _05233_;
wire _05234_;
wire _05235_;
wire _05236_;
wire _05237_;
wire _05238_;
wire _05239_;
wire _05240_;
wire _05241_;
wire _05242_;
wire _05243_;
wire _05244_;
wire _05245_;
wire _05246_;
wire _05247_;
wire _05248_;
wire _05249_;
wire _05250_;
wire _05251_;
wire _05252_;
wire _05253_;
wire _05254_;
wire _05255_;
wire _05256_;
wire _05257_;
wire _05258_;
wire _05259_;
wire _05260_;
wire _05261_;
wire _05262_;
wire _05263_;
wire _05264_;
wire _05265_;
wire _05266_;
wire _05267_;
wire _05268_;
wire _05269_;
wire _05270_;
wire _05271_;
wire _05272_;
wire _05273_;
wire _05274_;
wire _05275_;
wire _05276_;
wire _05277_;
wire _05278_;
wire _05279_;
wire _05280_;
wire _05281_;
wire _05282_;
wire _05283_;
wire _05284_;
wire _05285_;
wire _05286_;
wire _05287_;
wire _05288_;
wire _05289_;
wire _05290_;
wire _05291_;
wire _05292_;
wire _05293_;
wire _05294_;
wire _05295_;
wire _05296_;
wire _05297_;
wire _05298_;
wire _05299_;
wire _05300_;
wire _05301_;
wire _05302_;
wire _05303_;
wire _05304_;
wire _05305_;
wire _05306_;
wire _05307_;
wire _05308_;
wire _05309_;
wire _05310_;
wire _05311_;
wire _05312_;
wire _05313_;
wire _05314_;
wire _05315_;
wire _05316_;
wire _05317_;
wire _05318_;
wire _05319_;
wire _05320_;
wire _05321_;
wire _05322_;
wire _05323_;
wire _05324_;
wire _05325_;
wire _05326_;
wire _05327_;
wire _05328_;
wire _05329_;
wire _05330_;
wire _05331_;
wire _05332_;
wire _05333_;
wire _05334_;
wire _05335_;
wire _05336_;
wire _05337_;
wire _05338_;
wire _05339_;
wire _05340_;
wire _05341_;
wire _05342_;
wire _05343_;
wire _05344_;
wire _05345_;
wire _05346_;
wire _05347_;
wire _05348_;
wire _05349_;
wire _05350_;
wire _05351_;
wire _05352_;
wire _05353_;
wire _05354_;
wire _05355_;
wire _05356_;
wire _05357_;
wire _05358_;
wire _05359_;
wire _05360_;
wire _05361_;
wire _05362_;
wire _05363_;
wire _05364_;
wire _05365_;
wire _05366_;
wire _05367_;
wire _05368_;
wire _05369_;
wire _05370_;
wire _05371_;
wire _05372_;
wire _05373_;
wire _05374_;
wire _05375_;
wire _05376_;
wire _05377_;
wire _05378_;
wire _05379_;
wire _05380_;
wire _05381_;
wire _05382_;
wire _05383_;
wire _05384_;
wire _05385_;
wire _05386_;
wire _05387_;
wire _05388_;
wire _05389_;
wire _05390_;
wire _05391_;
wire _05392_;
wire _05393_;
wire _05394_;
wire _05395_;
wire _05396_;
wire _05397_;
wire _05398_;
wire _05399_;
wire _05400_;
wire _05401_;
wire _05402_;
wire _05403_;
wire _05404_;
wire _05405_;
wire _05406_;
wire _05407_;
wire _05408_;
wire _05409_;
wire _05410_;
wire _05411_;
wire _05412_;
wire _05413_;
wire _05414_;
wire _05415_;
wire _05416_;
wire _05417_;
wire _05418_;
wire _05419_;
wire _05420_;
wire _05421_;
wire _05422_;
wire _05423_;
wire _05424_;
wire _05425_;
wire _05426_;
wire _05427_;
wire _05428_;
wire _05429_;
wire _05430_;
wire _05431_;
wire _05432_;
wire _05433_;
wire _05434_;
wire _05435_;
wire _05436_;
wire _05437_;
wire _05438_;
wire _05439_;
wire _05440_;
wire _05441_;
wire _05442_;
wire _05443_;
wire _05444_;
wire _05445_;
wire _05446_;
wire _05447_;
wire _05448_;
wire _05449_;
wire _05450_;
wire _05451_;
wire _05452_;
wire _05453_;
wire _05454_;
wire _05455_;
wire _05456_;
wire _05457_;
wire _05458_;
wire _05459_;
wire _05460_;
wire _05461_;
wire _05462_;
wire _05463_;
wire _05464_;
wire _05465_;
wire _05466_;
wire _05467_;
wire _05468_;
wire _05469_;
wire _05470_;
wire _05471_;
wire _05472_;
wire _05473_;
wire _05474_;
wire _05475_;
wire _05476_;
wire _05477_;
wire _05478_;
wire _05479_;
wire _05480_;
wire _05481_;
wire _05482_;
wire _05483_;
wire _05484_;
wire _05485_;
wire _05486_;
wire _05487_;
wire _05488_;
wire _05489_;
wire _05490_;
wire _05491_;
wire _05492_;
wire _05493_;
wire _05494_;
wire _05495_;
wire _05496_;
wire _05497_;
wire _05498_;
wire _05499_;
wire _05500_;
wire _05501_;
wire _05502_;
wire _05503_;
wire _05504_;
wire _05505_;
wire _05506_;
wire _05507_;
wire _05508_;
wire _05509_;
wire _05510_;
wire _05511_;
wire _05512_;
wire _05513_;
wire _05514_;
wire _05515_;
wire _05516_;
wire _05517_;
wire _05518_;
wire _05519_;
wire _05520_;
wire _05521_;
wire _05522_;
wire _05523_;
wire _05524_;
wire _05525_;
wire _05526_;
wire _05527_;
wire _05528_;
wire _05529_;
wire _05530_;
wire _05531_;
wire _05532_;
wire _05533_;
wire _05534_;
wire _05535_;
wire _05536_;
wire _05537_;
wire _05538_;
wire _05539_;
wire _05540_;
wire _05541_;
wire _05542_;
wire _05543_;
wire _05544_;
wire _05545_;
wire _05546_;
wire _05547_;
wire _05548_;
wire _05549_;
wire _05550_;
wire _05551_;
wire _05552_;
wire _05553_;
wire _05554_;
wire _05555_;
wire _05556_;
wire _05557_;
wire _05558_;
wire _05559_;
wire _05560_;
wire _05561_;
wire _05562_;
wire _05563_;
wire _05564_;
wire _05565_;
wire _05566_;
wire _05567_;
wire _05568_;
wire _05569_;
wire _05570_;
wire _05571_;
wire _05572_;
wire _05573_;
wire _05574_;
wire _05575_;
wire _05576_;
wire _05577_;
wire _05578_;
wire _05579_;
wire _05580_;
wire _05581_;
wire _05582_;
wire _05583_;
wire _05584_;
wire _05585_;
wire _05586_;
wire _05587_;
wire _05588_;
wire _05589_;
wire _05590_;
wire _05591_;
wire _05592_;
wire _05593_;
wire _05594_;
wire _05595_;
wire _05596_;
wire _05597_;
wire _05598_;
wire _05599_;
wire _05600_;
wire _05601_;
wire _05602_;
wire _05603_;
wire _05604_;
wire _05605_;
wire _05606_;
wire _05607_;
wire _05608_;
wire _05609_;
wire _05610_;
wire _05611_;
wire _05612_;
wire _05613_;
wire _05614_;
wire _05615_;
wire _05616_;
wire _05617_;
wire _05618_;
wire _05619_;
wire _05620_;
wire _05621_;
wire _05622_;
wire _05623_;
wire _05624_;
wire _05625_;
wire _05626_;
wire _05627_;
wire _05628_;
wire _05629_;
wire _05630_;
wire _05631_;
wire _05632_;
wire _05633_;
wire _05634_;
wire _05635_;
wire _05636_;
wire _05637_;
wire _05638_;
wire _05639_;
wire _05640_;
wire _05641_;
wire _05642_;
wire _05643_;
wire _05644_;
wire _05645_;
wire _05646_;
wire _05647_;
wire _05648_;
wire _05649_;
wire _05650_;
wire _05651_;
wire _05652_;
wire _05653_;
wire _05654_;
wire _05655_;
wire _05656_;
wire _05657_;
wire _05658_;
wire _05659_;
wire _05660_;
wire _05661_;
wire _05662_;
wire _05663_;
wire _05664_;
wire _05665_;
wire _05666_;
wire _05667_;
wire _05668_;
wire _05669_;
wire _05670_;
wire _05671_;
wire _05672_;
wire _05673_;
wire _05674_;
wire _05675_;
wire _05676_;
wire _05677_;
wire _05678_;
wire _05679_;
wire _05680_;
wire _05681_;
wire _05682_;
wire _05683_;
wire _05684_;
wire _05685_;
wire _05686_;
wire _05687_;
wire _05688_;
wire _05689_;
wire _05690_;
wire _05691_;
wire _05692_;
wire _05693_;
wire _05694_;
wire _05695_;
wire _05696_;
wire _05697_;
wire _05698_;
wire _05699_;
wire _05700_;
wire _05701_;
wire _05702_;
wire _05703_;
wire _05704_;
wire _05705_;
wire _05706_;
wire _05707_;
wire _05708_;
wire _05709_;
wire _05710_;
wire _05711_;
wire _05712_;
wire _05713_;
wire _05714_;
wire _05715_;
wire _05716_;
wire _05717_;
wire _05718_;
wire _05719_;
wire _05720_;
wire _05721_;
wire _05722_;
wire _05723_;
wire _05724_;
wire _05725_;
wire _05726_;
wire _05727_;
wire _05728_;
wire _05729_;
wire _05730_;
wire _05731_;
wire _05732_;
wire _05733_;
wire _05734_;
wire _05735_;
wire _05736_;
wire _05737_;
wire _05738_;
wire _05739_;
wire _05740_;
wire _05741_;
wire _05742_;
wire _05743_;
wire _05744_;
wire _05745_;
wire _05746_;
wire _05747_;
wire _05748_;
wire _05749_;
wire _05750_;
wire _05751_;
wire _05752_;
wire _05753_;
wire _05754_;
wire _05755_;
wire _05756_;
wire _05757_;
wire _05758_;
wire _05759_;
wire _05760_;
wire _05761_;
wire _05762_;
wire _05763_;
wire _05764_;
wire _05765_;
wire _05766_;
wire _05767_;
wire _05768_;
wire _05769_;
wire _05770_;
wire _05771_;
wire _05772_;
wire _05773_;
wire _05774_;
wire _05775_;
wire _05776_;
wire _05777_;
wire _05778_;
wire _05779_;
wire _05780_;
wire _05781_;
wire _05782_;
wire _05783_;
wire _05784_;
wire _05785_;
wire _05786_;
wire _05787_;
wire _05788_;
wire _05789_;
wire _05790_;
wire _05791_;
wire _05792_;
wire _05793_;
wire _05794_;
wire _05795_;
wire _05796_;
wire _05797_;
wire _05798_;
wire _05799_;
wire _05800_;
wire _05801_;
wire _05802_;
wire _05803_;
wire _05804_;
wire _05805_;
wire _05806_;
wire _05807_;
wire _05808_;
wire _05809_;
wire _05810_;
wire _05811_;
wire _05812_;
wire _05813_;
wire _05814_;
wire _05815_;
wire _05816_;
wire _05817_;
wire _05818_;
wire _05819_;
wire _05820_;
wire _05821_;
wire _05822_;
wire _05823_;
wire _05824_;
wire _05825_;
wire _05826_;
wire _05827_;
wire _05828_;
wire _05829_;
wire _05830_;
wire _05831_;
wire _05832_;
wire _05833_;
wire _05834_;
wire _05835_;
wire _05836_;
wire _05837_;
wire _05838_;
wire _05839_;
wire _05840_;
wire _05841_;
wire _05842_;
wire _05843_;
wire _05844_;
wire _05845_;
wire _05846_;
wire _05847_;
wire _05848_;
wire _05849_;
wire _05850_;
wire _05851_;
wire _05852_;
wire _05853_;
wire _05854_;
wire _05855_;
wire _05856_;
wire _05857_;
wire _05858_;
wire _05859_;
wire _05860_;
wire _05861_;
wire _05862_;
wire _05863_;
wire _05864_;
wire _05865_;
wire _05866_;
wire _05867_;
wire _05868_;
wire _05869_;
wire _05870_;
wire _05871_;
wire _05872_;
wire _05873_;
wire _05874_;
wire _05875_;
wire _05876_;
wire _05877_;
wire _05878_;
wire _05879_;
wire _05880_;
wire _05881_;
wire _05882_;
wire _05883_;
wire _05884_;
wire _05885_;
wire _05886_;
wire _05887_;
wire _05888_;
wire _05889_;
wire _05890_;
wire _05891_;
wire _05892_;
wire _05893_;
wire _05894_;
wire _05895_;
wire _05896_;
wire _05897_;
wire _05898_;
wire _05899_;
wire _05900_;
wire _05901_;
wire _05902_;
wire _05903_;
wire _05904_;
wire _05905_;
wire _05906_;
wire _05907_;
wire _05908_;
wire _05909_;
wire _05910_;
wire _05911_;
wire _05912_;
wire _05913_;
wire _05914_;
wire _05915_;
wire _05916_;
wire _05917_;
wire _05918_;
wire _05919_;
wire _05920_;
wire _05921_;
wire _05922_;
wire _05923_;
wire _05924_;
wire _05925_;
wire _05926_;
wire _05927_;
wire _05928_;
wire _05929_;
wire _05930_;
wire _05931_;
wire _05932_;
wire _05933_;
wire _05934_;
wire _05935_;
wire _05936_;
wire _05937_;
wire _05938_;
wire _05939_;
wire _05940_;
wire _05941_;
wire _05942_;
wire _05943_;
wire _05944_;
wire _05945_;
wire _05946_;
wire _05947_;
wire _05948_;
wire _05949_;
wire _05950_;
wire _05951_;
wire _05952_;
wire _05953_;
wire _05954_;
wire _05955_;
wire _05956_;
wire _05957_;
wire _05958_;
wire _05959_;
wire _05960_;
wire _05961_;
wire _05962_;
wire _05963_;
wire _05964_;
wire _05965_;
wire _05966_;
wire _05967_;
wire _05968_;
wire _05969_;
wire _05970_;
wire _05971_;
wire _05972_;
wire _05973_;
wire _05974_;
wire _05975_;
wire _05976_;
wire _05977_;
wire _05978_;
wire _05979_;
wire _05980_;
wire _05981_;
wire _05982_;
wire _05983_;
wire _05984_;
wire _05985_;
wire _05986_;
wire _05987_;
wire _05988_;
wire _05989_;
wire _05990_;
wire _05991_;
wire _05992_;
wire _05993_;
wire _05994_;
wire _05995_;
wire _05996_;
wire _05997_;
wire _05998_;
wire _05999_;
wire _06000_;
wire _06001_;
wire _06002_;
wire _06003_;
wire _06004_;
wire _06005_;
wire _06006_;
wire _06007_;
wire _06008_;
wire _06009_;
wire _06010_;
wire _06011_;
wire _06012_;
wire _06013_;
wire _06014_;
wire _06015_;
wire _06016_;
wire _06017_;
wire _06018_;
wire _06019_;
wire _06020_;
wire _06021_;
wire _06022_;
wire _06023_;
wire _06024_;
wire _06025_;
wire _06026_;
wire _06027_;
wire _06028_;
wire _06029_;
wire _06030_;
wire _06031_;
wire _06032_;
wire _06033_;
wire _06034_;
wire _06035_;
wire _06036_;
wire _06037_;
wire _06038_;
wire _06039_;
wire _06040_;
wire _06041_;
wire _06042_;
wire _06043_;
wire _06044_;
wire _06045_;
wire _06046_;
wire _06047_;
wire _06048_;
wire _06049_;
wire _06050_;
wire _06051_;
wire _06052_;
wire _06053_;
wire _06054_;
wire _06055_;
wire _06056_;
wire _06057_;
wire _06058_;
wire _06059_;
wire _06060_;
wire _06061_;
wire _06062_;
wire _06063_;
wire _06064_;
wire _06065_;
wire _06066_;
wire _06067_;
wire _06068_;
wire _06069_;
wire _06070_;
wire _06071_;
wire _06072_;
wire _06073_;
wire _06074_;
wire _06075_;
wire _06076_;
wire _06077_;
wire _06078_;
wire _06079_;
wire _06080_;
wire _06081_;
wire _06082_;
wire _06083_;
wire _06084_;
wire _06085_;
wire _06086_;
wire _06087_;
wire _06088_;
wire _06089_;
wire _06090_;
wire _06091_;
wire _06092_;
wire _06093_;
wire _06094_;
wire _06095_;
wire _06096_;
wire _06097_;
wire _06098_;
wire _06099_;
wire _06100_;
wire _06101_;
wire _06102_;
wire _06103_;
wire _06104_;
wire _06105_;
wire _06106_;
wire _06107_;
wire _06108_;
wire _06109_;
wire _06110_;
wire _06111_;
wire _06112_;
wire _06113_;
wire _06114_;
wire _06115_;
wire _06116_;
wire _06117_;
wire _06118_;
wire _06119_;
wire _06120_;
wire _06121_;
wire _06122_;
wire _06123_;
wire _06124_;
wire _06125_;
wire _06126_;
wire _06127_;
wire _06128_;
wire _06129_;
wire _06130_;
wire _06131_;
wire _06132_;
wire _06133_;
wire _06134_;
wire _06135_;
wire _06136_;
wire _06137_;
wire _06138_;
wire _06139_;
wire _06140_;
wire _06141_;
wire _06142_;
wire _06143_;
wire _06144_;
wire _06145_;
wire _06146_;
wire _06147_;
wire _06148_;
wire _06149_;
wire _06150_;
wire _06151_;
wire _06152_;
wire _06153_;
wire _06154_;
wire _06155_;
wire _06156_;
wire _06157_;
wire _06158_;
wire _06159_;
wire _06160_;
wire _06161_;
wire _06162_;
wire _06163_;
wire _06164_;
wire _06165_;
wire _06166_;
wire _06167_;
wire _06168_;
wire _06169_;
wire _06170_;
wire _06171_;
wire _06172_;
wire _06173_;
wire _06174_;
wire _06175_;
wire _06176_;
wire _06177_;
wire _06178_;
wire _06179_;
wire _06180_;
wire _06181_;
wire _06182_;
wire _06183_;
wire _06184_;
wire _06185_;
wire _06186_;
wire _06187_;
wire _06188_;
wire _06189_;
wire _06190_;
wire _06191_;
wire _06192_;
wire _06193_;
wire _06194_;
wire _06195_;
wire _06196_;
wire _06197_;
wire _06198_;
wire _06199_;
wire _06200_;
wire _06201_;
wire _06202_;
wire _06203_;
wire _06204_;
wire _06205_;
wire _06206_;
wire _06207_;
wire _06208_;
wire _06209_;
wire _06210_;
wire _06211_;
wire _06212_;
wire _06213_;
wire _06214_;
wire _06215_;
wire _06216_;
wire _06217_;
wire _06218_;
wire _06219_;
wire _06220_;
wire _06221_;
wire _06222_;
wire _06223_;
wire _06224_;
wire _06225_;
wire _06226_;
wire _06227_;
wire _06228_;
wire _06229_;
wire _06230_;
wire _06231_;
wire _06232_;
wire _06233_;
wire _06234_;
wire _06235_;
wire _06236_;
wire _06237_;
wire _06238_;
wire _06239_;
wire _06240_;
wire _06241_;
wire _06242_;
wire _06243_;
wire _06244_;
wire _06245_;
wire _06246_;
wire _06247_;
wire _06248_;
wire _06249_;
wire _06250_;
wire _06251_;
wire _06252_;
wire _06253_;
wire _06254_;
wire _06255_;
wire _06256_;
wire _06257_;
wire _06258_;
wire _06259_;
wire _06260_;
wire _06261_;
wire _06262_;
wire _06263_;
wire _06264_;
wire _06265_;
wire _06266_;
wire _06267_;
wire _06268_;
wire _06269_;
wire _06270_;
wire _06271_;
wire _06272_;
wire _06273_;
wire _06274_;
wire _06275_;
wire _06276_;
wire _06277_;
wire _06278_;
wire _06279_;
wire _06280_;
wire _06281_;
wire _06282_;
wire _06283_;
wire _06284_;
wire _06285_;
wire _06286_;
wire _06287_;
wire _06288_;
wire _06289_;
wire _06290_;
wire _06291_;
wire _06292_;
wire _06293_;
wire _06294_;
wire _06295_;
wire _06296_;
wire _06297_;
wire _06298_;
wire _06299_;
wire _06300_;
wire _06301_;
wire _06302_;
wire _06303_;
wire _06304_;
wire _06305_;
wire _06306_;
wire _06307_;
wire _06308_;
wire _06309_;
wire _06310_;
wire _06311_;
wire _06312_;
wire _06313_;
wire _06314_;
wire _06315_;
wire _06316_;
wire _06317_;
wire _06318_;
wire _06319_;
wire _06320_;
wire _06321_;
wire _06322_;
wire _06323_;
wire _06324_;
wire _06325_;
wire _06326_;
wire _06327_;
wire _06328_;
wire _06329_;
wire _06330_;
wire _06331_;
wire _06332_;
wire _06333_;
wire _06334_;
wire _06335_;
wire _06336_;
wire _06337_;
wire _06338_;
wire _06339_;
wire _06340_;
wire _06341_;
wire _06342_;
wire _06343_;
wire _06344_;
wire _06345_;
wire _06346_;
wire _06347_;
wire _06348_;
wire _06349_;
wire _06350_;
wire _06351_;
wire _06352_;
wire _06353_;
wire _06354_;
wire _06355_;
wire _06356_;
wire _06357_;
wire _06358_;
wire _06359_;
wire _06360_;
wire _06361_;
wire _06362_;
wire _06363_;
wire _06364_;
wire _06365_;
wire _06366_;
wire _06367_;
wire _06368_;
wire _06369_;
wire _06370_;
wire _06371_;
wire _06372_;
wire _06373_;
wire _06374_;
wire _06375_;
wire _06376_;
wire _06377_;
wire _06378_;
wire _06379_;
wire _06380_;
wire _06381_;
wire _06382_;
wire _06383_;
wire _06384_;
wire _06385_;
wire _06386_;
wire _06387_;
wire _06388_;
wire _06389_;
wire _06390_;
wire _06391_;
wire _06392_;
wire _06393_;
wire _06394_;
wire _06395_;
wire _06396_;
wire _06397_;
wire _06398_;
wire _06399_;
wire _06400_;
wire _06401_;
wire _06402_;
wire _06403_;
wire _06404_;
wire _06405_;
wire _06406_;
wire _06407_;
wire _06408_;
wire _06409_;
wire _06410_;
wire _06411_;
wire _06412_;
wire _06413_;
wire _06414_;
wire _06415_;
wire _06416_;
wire _06417_;
wire _06418_;
wire _06419_;
wire _06420_;
wire _06421_;
wire _06422_;
wire _06423_;
wire _06424_;
wire _06425_;
wire _06426_;
wire _06427_;
wire _06428_;
wire _06429_;
wire _06430_;
wire _06431_;
wire _06432_;
wire _06433_;
wire _06434_;
wire _06435_;
wire _06436_;
wire _06437_;
wire _06438_;
wire _06439_;
wire _06440_;
wire _06441_;
wire _06442_;
wire _06443_;
wire _06444_;
wire _06445_;
wire _06446_;
wire _06447_;
wire _06448_;
wire _06449_;
wire _06450_;
wire _06451_;
wire _06452_;
wire _06453_;
wire _06454_;
wire _06455_;
wire _06456_;
wire _06457_;
wire _06458_;
wire _06459_;
wire _06460_;
wire _06461_;
wire _06462_;
wire _06463_;
wire _06464_;
wire _06465_;
wire _06466_;
wire _06467_;
wire _06468_;
wire _06469_;
wire _06470_;
wire _06471_;
wire _06472_;
wire _06473_;
wire _06474_;
wire _06475_;
wire _06476_;
wire _06477_;
wire _06478_;
wire _06479_;
wire _06480_;
wire _06481_;
wire _06482_;
wire _06483_;
wire _06484_;
wire _06485_;
wire _06486_;
wire _06487_;
wire _06488_;
wire _06489_;
wire _06490_;
wire _06491_;
wire _06492_;
wire _06493_;
wire _06494_;
wire _06495_;
wire _06496_;
wire _06497_;
wire _06498_;
wire _06499_;
wire _06500_;
wire _06501_;
wire _06502_;
wire _06503_;
wire _06504_;
wire _06505_;
wire _06506_;
wire _06507_;
wire _06508_;
wire _06509_;
wire _06510_;
wire _06511_;
wire _06512_;
wire _06513_;
wire _06514_;
wire _06515_;
wire _06516_;
wire _06517_;
wire _06518_;
wire _06519_;
wire _06520_;
wire _06521_;
wire _06522_;
wire _06523_;
wire _06524_;
wire _06525_;
wire _06526_;
wire _06527_;
wire _06528_;
wire _06529_;
wire _06530_;
wire _06531_;
wire _06532_;
wire _06533_;
wire _06534_;
wire _06535_;
wire _06536_;
wire _06537_;
wire _06538_;
wire _06539_;
wire _06540_;
wire _06541_;
wire _06542_;
wire _06543_;
wire _06544_;
wire _06545_;
wire _06546_;
wire _06547_;
wire _06548_;
wire _06549_;
wire _06550_;
wire _06551_;
wire _06552_;
wire _06553_;
wire _06554_;
wire _06555_;
wire _06556_;
wire _06557_;
wire _06558_;
wire _06559_;
wire _06560_;
wire _06561_;
wire _06562_;
wire _06563_;
wire _06564_;
wire _06565_;
wire _06566_;
wire _06567_;
wire _06568_;
wire _06569_;
wire _06570_;
wire _06571_;
wire _06572_;
wire _06573_;
wire _06574_;
wire _06575_;
wire _06576_;
wire _06577_;
wire _06578_;
wire _06579_;
wire _06580_;
wire _06581_;
wire _06582_;
wire _06583_;
wire _06584_;
wire _06585_;
wire _06586_;
wire _06587_;
wire _06588_;
wire _06589_;
wire _06590_;
wire _06591_;
wire _06592_;
wire _06593_;
wire _06594_;
wire _06595_;
wire _06596_;
wire _06597_;
wire _06598_;
wire _06599_;
wire _06600_;
wire _06601_;
wire _06602_;
wire _06603_;
wire _06604_;
wire _06605_;
wire _06606_;
wire _06607_;
wire _06608_;
wire _06609_;
wire _06610_;
wire _06611_;
wire _06612_;
wire _06613_;
wire _06614_;
wire _06615_;
wire _06616_;
wire _06617_;
wire _06618_;
wire _06619_;
wire _06620_;
wire _06621_;
wire _06622_;
wire _06623_;
wire _06624_;
wire _06625_;
wire _06626_;
wire _06627_;
wire _06628_;
wire _06629_;
wire _06630_;
wire _06631_;
wire _06632_;
wire _06633_;
wire _06634_;
wire _06635_;
wire _06636_;
wire _06637_;
wire _06638_;
wire _06639_;
wire _06640_;
wire _06641_;
wire _06642_;
wire _06643_;
wire _06644_;
wire _06645_;
wire _06646_;
wire _06647_;
wire _06648_;
wire _06649_;
wire _06650_;
wire _06651_;
wire _06652_;
wire _06653_;
wire _06654_;
wire _06655_;
wire _06656_;
wire _06657_;
wire _06658_;
wire _06659_;
wire _06660_;
wire _06661_;
wire _06662_;
wire _06663_;
wire _06664_;
wire _06665_;
wire _06666_;
wire _06667_;
wire _06668_;
wire _06669_;
wire _06670_;
wire _06671_;
wire _06672_;
wire _06673_;
wire _06674_;
wire _06675_;
wire _06676_;
wire _06677_;
wire _06678_;
wire _06679_;
wire _06680_;
wire _06681_;
wire _06682_;
wire _06683_;
wire _06684_;
wire _06685_;
wire _06686_;
wire _06687_;
wire _06688_;
wire _06689_;
wire _06690_;
wire _06691_;
wire _06692_;
wire _06693_;
wire _06694_;
wire _06695_;
wire _06696_;
wire _06697_;
wire _06698_;
wire _06699_;
wire _06700_;
wire _06701_;
wire _06702_;
wire _06703_;
wire _06704_;
wire _06705_;
wire _06706_;
wire _06707_;
wire _06708_;
wire _06709_;
wire _06710_;
wire _06711_;
wire _06712_;
wire _06713_;
wire _06714_;
wire _06715_;
wire _06716_;
wire _06717_;
wire _06718_;
wire _06719_;
wire _06720_;
wire _06721_;
wire _06722_;
wire _06723_;
wire _06724_;
wire _06725_;
wire _06726_;
wire _06727_;
wire _06728_;
wire _06729_;
wire _06730_;
wire _06731_;
wire _06732_;
wire _06733_;
wire _06734_;
wire _06735_;
wire _06736_;
wire _06737_;
wire _06738_;
wire _06739_;
wire _06740_;
wire _06741_;
wire _06742_;
wire _06743_;
wire _06744_;
wire _06745_;
wire _06746_;
wire _06747_;
wire _06748_;
wire _06749_;
wire _06750_;
wire _06751_;
wire _06752_;
wire _06753_;
wire _06754_;
wire _06755_;
wire _06756_;
wire _06757_;
wire _06758_;
wire _06759_;
wire _06760_;
wire _06761_;
wire _06762_;
wire _06763_;
wire _06764_;
wire _06765_;
wire _06766_;
wire _06767_;
wire _06768_;
wire _06769_;
wire _06770_;
wire _06771_;
wire _06772_;
wire _06773_;
wire _06774_;
wire _06775_;
wire _06776_;
wire _06777_;
wire _06778_;
wire _06779_;
wire _06780_;
wire _06781_;
wire _06782_;
wire _06783_;
wire _06784_;
wire _06785_;
wire _06786_;
wire _06787_;
wire _06788_;
wire _06789_;
wire _06790_;
wire _06791_;
wire _06792_;
wire _06793_;
wire _06794_;
wire _06795_;
wire _06796_;
wire _06797_;
wire _06798_;
wire _06799_;
wire _06800_;
wire _06801_;
wire _06802_;
wire _06803_;
wire _06804_;
wire _06805_;
wire _06806_;
wire _06807_;
wire _06808_;
wire _06809_;
wire _06810_;
wire _06811_;
wire _06812_;
wire _06813_;
wire _06814_;
wire _06815_;
wire _06816_;
wire _06817_;
wire _06818_;
wire _06819_;
wire _06820_;
wire _06821_;
wire _06822_;
wire _06823_;
wire _06824_;
wire _06825_;
wire _06826_;
wire _06827_;
wire _06828_;
wire _06829_;
wire _06830_;
wire _06831_;
wire _06832_;
wire _06833_;
wire _06834_;
wire _06835_;
wire _06836_;
wire _06837_;
wire _06838_;
wire _06839_;
wire _06840_;
wire _06841_;
wire _06842_;
wire _06843_;
wire _06844_;
wire _06845_;
wire _06846_;
wire _06847_;
wire _06848_;
wire _06849_;
wire _06850_;
wire _06851_;
wire _06852_;
wire _06853_;
wire _06854_;
wire _06855_;
wire _06856_;
wire _06857_;
wire _06858_;
wire _06859_;
wire _06860_;
wire _06861_;
wire _06862_;
wire _06863_;
wire _06864_;
wire _06865_;
wire _06866_;
wire _06867_;
wire _06868_;
wire _06869_;
wire _06870_;
wire _06871_;
wire _06872_;
wire _06873_;
wire _06874_;
wire _06875_;
wire _06876_;
wire _06877_;
wire _06878_;
wire _06879_;
wire _06880_;
wire _06881_;
wire _06882_;
wire _06883_;
wire _06884_;
wire _06885_;
wire _06886_;
wire _06887_;
wire _06888_;
wire _06889_;
wire _06890_;
wire _06891_;
wire _06892_;
wire _06893_;
wire _06894_;
wire _06895_;
wire _06896_;
wire _06897_;
wire _06898_;
wire _06899_;
wire _06900_;
wire _06901_;
wire _06902_;
wire _06903_;
wire _06904_;
wire _06905_;
wire _06906_;
wire _06907_;
wire _06908_;
wire _06909_;
wire _06910_;
wire _06911_;
wire _06912_;
wire _06913_;
wire _06914_;
wire _06915_;
wire _06916_;
wire _06917_;
wire _06918_;
wire _06919_;
wire _06920_;
wire _06921_;
wire _06922_;
wire _06923_;
wire _06924_;
wire _06925_;
wire _06926_;
wire _06927_;
wire _06928_;
wire _06929_;
wire _06930_;
wire _06931_;
wire _06932_;
wire _06933_;
wire _06934_;
wire _06935_;
wire _06936_;
wire _06937_;
wire _06938_;
wire _06939_;
wire _06940_;
wire _06941_;
wire _06942_;
wire _06943_;
wire _06944_;
wire _06945_;
wire _06946_;
wire _06947_;
wire _06948_;
wire _06949_;
wire _06950_;
wire _06951_;
wire _06952_;
wire _06953_;
wire _06954_;
wire _06955_;
wire _06956_;
wire _06957_;
wire _06958_;
wire _06959_;
wire _06960_;
wire _06961_;
wire _06962_;
wire _06963_;
wire _06964_;
wire _06965_;
wire _06966_;
wire _06967_;
wire _06968_;
wire _06969_;
wire _06970_;
wire _06971_;
wire _06972_;
wire _06973_;
wire _06974_;
wire _06975_;
wire _06976_;
wire _06977_;
wire _06978_;
wire _06979_;
wire _06980_;
wire _06981_;
wire _06982_;
wire _06983_;
wire _06984_;
wire _06985_;
wire _06986_;
wire _06987_;
wire _06988_;
wire _06989_;
wire _06990_;
wire _06991_;
wire _06992_;
wire _06993_;
wire _06994_;
wire _06995_;
wire _06996_;
wire _06997_;
wire _06998_;
wire _06999_;
wire _07000_;
wire _07001_;
wire _07002_;
wire _07003_;
wire _07004_;
wire _07005_;
wire _07006_;
wire _07007_;
wire _07008_;
wire _07009_;
wire _07010_;
wire _07011_;
wire _07012_;
wire _07013_;
wire _07014_;
wire _07015_;
wire _07016_;
wire _07017_;
wire _07018_;
wire _07019_;
wire _07020_;
wire _07021_;
wire _07022_;
wire _07023_;
wire _07024_;
wire _07025_;
wire _07026_;
wire _07027_;
wire _07028_;
wire _07029_;
wire _07030_;
wire _07031_;
wire _07032_;
wire _07033_;
wire _07034_;
wire _07035_;
wire _07036_;
wire _07037_;
wire _07038_;
wire _07039_;
wire _07040_;
wire _07041_;
wire _07042_;
wire _07043_;
wire _07044_;
wire _07045_;
wire _07046_;
wire _07047_;
wire _07048_;
wire _07049_;
wire _07050_;
wire _07051_;
wire _07052_;
wire _07053_;
wire _07054_;
wire _07055_;
wire _07056_;
wire _07057_;
wire _07058_;
wire _07059_;
wire _07060_;
wire _07061_;
wire _07062_;
wire _07063_;
wire _07064_;
wire _07065_;
wire _07066_;
wire _07067_;
wire _07068_;
wire _07069_;
wire _07070_;
wire _07071_;
wire _07072_;
wire _07073_;
wire _07074_;
wire _07075_;
wire _07076_;
wire _07077_;
wire _07078_;
wire _07079_;
wire _07080_;
wire _07081_;
wire _07082_;
wire _07083_;
wire _07084_;
wire _07085_;
wire _07086_;
wire _07087_;
wire _07088_;
wire _07089_;
wire _07090_;
wire _07091_;
wire _07092_;
wire _07093_;
wire _07094_;
wire _07095_;
wire _07096_;
wire _07097_;
wire _07098_;
wire _07099_;
wire _07100_;
wire _07101_;
wire _07102_;
wire _07103_;
wire _07104_;
wire _07105_;
wire _07106_;
wire _07107_;
wire _07108_;
wire _07109_;
wire _07110_;
wire _07111_;
wire _07112_;
wire _07113_;
wire _07114_;
wire _07115_;
wire _07116_;
wire _07117_;
wire _07118_;
wire _07119_;
wire _07120_;
wire _07121_;
wire _07122_;
wire _07123_;
wire _07124_;
wire _07125_;
wire _07126_;
wire _07127_;
wire _07128_;
wire _07129_;
wire _07130_;
wire _07131_;
wire _07132_;
wire _07133_;
wire _07134_;
wire _07135_;
wire _07136_;
wire _07137_;
wire _07138_;
wire _07139_;
wire _07140_;
wire _07141_;
wire _07142_;
wire _07143_;
wire _07144_;
wire _07145_;
wire _07146_;
wire _07147_;
wire _07148_;
wire _07149_;
wire _07150_;
wire _07151_;
wire _07152_;
wire _07153_;
wire _07154_;
wire _07155_;
wire _07156_;
wire _07157_;
wire _07158_;
wire _07159_;
wire _07160_;
wire _07161_;
wire _07162_;
wire _07163_;
wire _07164_;
wire _07165_;
wire _07166_;
wire _07167_;
wire _07168_;
wire _07169_;
wire _07170_;
wire _07171_;
wire _07172_;
wire _07173_;
wire _07174_;
wire _07175_;
wire _07176_;
wire _07177_;
wire _07178_;
wire _07179_;
wire _07180_;
wire _07181_;
wire _07182_;
wire _07183_;
wire _07184_;
wire _07185_;
wire _07186_;
wire _07187_;
wire _07188_;
wire _07189_;
wire _07190_;
wire _07191_;
wire _07192_;
wire _07193_;
wire _07194_;
wire _07195_;
wire _07196_;
wire _07197_;
wire _07198_;
wire _07199_;
wire _07200_;
wire _07201_;
wire _07202_;
wire _07203_;
wire _07204_;
wire _07205_;
wire _07206_;
wire _07207_;
wire _07208_;
wire _07209_;
wire _07210_;
wire _07211_;
wire _07212_;
wire _07213_;
wire _07214_;
wire _07215_;
wire _07216_;
wire _07217_;
wire _07218_;
wire _07219_;
wire _07220_;
wire _07221_;
wire _07222_;
wire _07223_;
wire _07224_;
wire _07225_;
wire _07226_;
wire _07227_;
wire _07228_;
wire _07229_;
wire _07230_;
wire _07231_;
wire _07232_;
wire _07233_;
wire _07234_;
wire _07235_;
wire _07236_;
wire _07237_;
wire _07238_;
wire _07239_;
wire _07240_;
wire _07241_;
wire _07242_;
wire _07243_;
wire _07244_;
wire _07245_;
wire _07246_;
wire _07247_;
wire _07248_;
wire _07249_;
wire _07250_;
wire _07251_;
wire _07252_;
wire _07253_;
wire _07254_;
wire _07255_;
wire _07256_;
wire _07257_;
wire _07258_;
wire _07259_;
wire _07260_;
wire _07261_;
wire _07262_;
wire _07263_;
wire _07264_;
wire _07265_;
wire _07266_;
wire _07267_;
wire _07268_;
wire _07269_;
wire _07270_;
wire _07271_;
wire _07272_;
wire _07273_;
wire _07274_;
wire _07275_;
wire _07276_;
wire _07277_;
wire _07278_;
wire _07279_;
wire _07280_;
wire _07281_;
wire _07282_;
wire _07283_;
wire _07284_;
wire _07285_;
wire _07286_;
wire _07287_;
wire _07288_;
wire _07289_;
wire _07290_;
wire _07291_;
wire _07292_;
wire _07293_;
wire _07294_;
wire _07295_;
wire _07296_;
wire _07297_;
wire _07298_;
wire _07299_;
wire _07300_;
wire _07301_;
wire _07302_;
wire _07303_;
wire _07304_;
wire _07305_;
wire _07306_;
wire _07307_;
wire _07308_;
wire _07309_;
wire _07310_;
wire _07311_;
wire _07312_;
wire _07313_;
wire _07314_;
wire _07315_;
wire _07316_;
wire _07317_;
wire _07318_;
wire _07319_;
wire _07320_;
wire _07321_;
wire _07322_;
wire _07323_;
wire _07324_;
wire _07325_;
wire _07326_;
wire _07327_;
wire _07328_;
wire _07329_;
wire _07330_;
wire _07331_;
wire _07332_;
wire _07333_;
wire _07334_;
wire _07335_;
wire _07336_;
wire _07337_;
wire _07338_;
wire _07339_;
wire _07340_;
wire _07341_;
wire _07342_;
wire _07343_;
wire _07344_;
wire _07345_;
wire _07346_;
wire _07347_;
wire _07348_;
wire _07349_;
wire _07350_;
wire _07351_;
wire _07352_;
wire _07353_;
wire _07354_;
wire _07355_;
wire _07356_;
wire _07357_;
wire _07358_;
wire _07359_;
wire _07360_;
wire _07361_;
wire _07362_;
wire _07363_;
wire _07364_;
wire _07365_;
wire _07366_;
wire _07367_;
wire _07368_;
wire _07369_;
wire _07370_;
wire _07371_;
wire _07372_;
wire _07373_;
wire _07374_;
wire _07375_;
wire _07376_;
wire _07377_;
wire _07378_;
wire _07379_;
wire _07380_;
wire _07381_;
wire _07382_;
wire _07383_;
wire _07384_;
wire _07385_;
wire _07386_;
wire _07387_;
wire _07388_;
wire _07389_;
wire _07390_;
wire _07391_;
wire _07392_;
wire _07393_;
wire _07394_;
wire _07395_;
wire _07396_;
wire _07397_;
wire _07398_;
wire _07399_;
wire _07400_;
wire _07401_;
wire _07402_;
wire _07403_;
wire _07404_;
wire _07405_;
wire _07406_;
wire _07407_;
wire _07408_;
wire _07409_;
wire _07410_;
wire _07411_;
wire _07412_;
wire _07413_;
wire _07414_;
wire _07415_;
wire _07416_;
wire _07417_;
wire _07418_;
wire _07419_;
wire _07420_;
wire _07421_;
wire _07422_;
wire _07423_;
wire _07424_;
wire _07425_;
wire _07426_;
wire _07427_;
wire _07428_;
wire _07429_;
wire _07430_;
wire _07431_;
wire _07432_;
wire _07433_;
wire _07434_;
wire _07435_;
wire _07436_;
wire _07437_;
wire _07438_;
wire _07439_;
wire _07440_;
wire _07441_;
wire _07442_;
wire _07443_;
wire _07444_;
wire _07445_;
wire _07446_;
wire _07447_;
wire _07448_;
wire _07449_;
wire _07450_;
wire _07451_;
wire _07452_;
wire _07453_;
wire _07454_;
wire _07455_;
wire _07456_;
wire _07457_;
wire _07458_;
wire _07459_;
wire _07460_;
wire _07461_;
wire _07462_;
wire _07463_;
wire _07464_;
wire _07465_;
wire _07466_;
wire _07467_;
wire _07468_;
wire _07469_;
wire _07470_;
wire _07471_;
wire _07472_;
wire _07473_;
wire _07474_;
wire _07475_;
wire _07476_;
wire _07477_;
wire _07478_;
wire _07479_;
wire _07480_;
wire _07481_;
wire _07482_;
wire _07483_;
wire _07484_;
wire _07485_;
wire _07486_;
wire _07487_;
wire _07488_;
wire _07489_;
wire _07490_;
wire _07491_;
wire _07492_;
wire _07493_;
wire _07494_;
wire _07495_;
wire _07496_;
wire _07497_;
wire _07498_;
wire _07499_;
wire _07500_;
wire _07501_;
wire _07502_;
wire _07503_;
wire _07504_;
wire _07505_;
wire _07506_;
wire _07507_;
wire _07508_;
wire _07509_;
wire _07510_;
wire _07511_;
wire _07512_;
wire _07513_;
wire _07514_;
wire _07515_;
wire _07516_;
wire _07517_;
wire _07518_;
wire _07519_;
wire _07520_;
wire _07521_;
wire _07522_;
wire _07523_;
wire _07524_;
wire _07525_;
wire _07526_;
wire _07527_;
wire _07528_;
wire _07529_;
wire _07530_;
wire _07531_;
wire _07532_;
wire _07533_;
wire _07534_;
wire _07535_;
wire _07536_;
wire _07537_;
wire _07538_;
wire _07539_;
wire _07540_;
wire _07541_;
wire _07542_;
wire _07543_;
wire _07544_;
wire _07545_;
wire _07546_;
wire _07547_;
wire _07548_;
wire _07549_;
wire _07550_;
wire _07551_;
wire _07552_;
wire _07553_;
wire _07554_;
wire _07555_;
wire _07556_;
wire _07557_;
wire _07558_;
wire _07559_;
wire _07560_;
wire _07561_;
wire _07562_;
wire _07563_;
wire _07564_;
wire _07565_;
wire _07566_;
wire _07567_;
wire _07568_;
wire _07569_;
wire _07570_;
wire _07571_;
wire _07572_;
wire _07573_;
wire _07574_;
wire _07575_;
wire _07576_;
wire _07577_;
wire _07578_;
wire _07579_;
wire _07580_;
wire _07581_;
wire _07582_;
wire _07583_;
wire _07584_;
wire _07585_;
wire _07586_;
wire _07587_;
wire _07588_;
wire _07589_;
wire _07590_;
wire _07591_;
wire _07592_;
wire _07593_;
wire _07594_;
wire _07595_;
wire _07596_;
wire _07597_;
wire _07598_;
wire _07599_;
wire _07600_;
wire _07601_;
wire _07602_;
wire _07603_;
wire _07604_;
wire _07605_;
wire _07606_;
wire _07607_;
wire _07608_;
wire _07609_;
wire _07610_;
wire _07611_;
wire _07612_;
wire _07613_;
wire _07614_;
wire _07615_;
wire _07616_;
wire _07617_;
wire _07618_;
wire _07619_;
wire _07620_;
wire _07621_;
wire _07622_;
wire _07623_;
wire _07624_;
wire _07625_;
wire _07626_;
wire _07627_;
wire _07628_;
wire _07629_;
wire _07630_;
wire _07631_;
wire _07632_;
wire _07633_;
wire _07634_;
wire _07635_;
wire _07636_;
wire _07637_;
wire _07638_;
wire _07639_;
wire _07640_;
wire _07641_;
wire _07642_;
wire _07643_;
wire _07644_;
wire _07645_;
wire _07646_;
wire _07647_;
wire _07648_;
wire _07649_;
wire _07650_;
wire _07651_;
wire _07652_;
wire _07653_;
wire _07654_;
wire _07655_;
wire _07656_;
wire _07657_;
wire _07658_;
wire _07659_;
wire _07660_;
wire _07661_;
wire _07662_;
wire _07663_;
wire _07664_;
wire _07665_;
wire _07666_;
wire _07667_;
wire _07668_;
wire _07669_;
wire _07670_;
wire _07671_;
wire _07672_;
wire _07673_;
wire _07674_;
wire _07675_;
wire _07676_;
wire _07677_;
wire _07678_;
wire _07679_;
wire _07680_;
wire _07681_;
wire _07682_;
wire _07683_;
wire _07684_;
wire _07685_;
wire _07686_;
wire _07687_;
wire _07688_;
wire _07689_;
wire _07690_;
wire _07691_;
wire _07692_;
wire _07693_;
wire _07694_;
wire _07695_;
wire _07696_;
wire _07697_;
wire _07698_;
wire _07699_;
wire _07700_;
wire _07701_;
wire _07702_;
wire _07703_;
wire _07704_;
wire _07705_;
wire _07706_;
wire _07707_;
wire _07708_;
wire _07709_;
wire _07710_;
wire _07711_;
wire _07712_;
wire _07713_;
wire _07714_;
wire _07715_;
wire _07716_;
wire _07717_;
wire _07718_;
wire _07719_;
wire _07720_;
wire _07721_;
wire _07722_;
wire _07723_;
wire _07724_;
wire _07725_;
wire _07726_;
wire _07727_;
wire _07728_;
wire _07729_;
wire _07730_;
wire _07731_;
wire _07732_;
wire _07733_;
wire _07734_;
wire _07735_;
wire _07736_;
wire _07737_;
wire _07738_;
wire _07739_;
wire _07740_;
wire _07741_;
wire _07742_;
wire _07743_;
wire _07744_;
wire _07745_;
wire _07746_;
wire _07747_;
wire _07748_;
wire _07749_;
wire _07750_;
wire _07751_;
wire _07752_;
wire _07753_;
wire _07754_;
wire _07755_;
wire _07756_;
wire _07757_;
wire _07758_;
wire _07759_;
wire _07760_;
wire _07761_;
wire _07762_;
wire _07763_;
wire _07764_;
wire _07765_;
wire _07766_;
wire _07767_;
wire _07768_;
wire _07769_;
wire _07770_;
wire _07771_;
wire _07772_;
wire _07773_;
wire _07774_;
wire _07775_;
wire _07776_;
wire _07777_;
wire _07778_;
wire _07779_;
wire _07780_;
wire _07781_;
wire _07782_;
wire _07783_;
wire _07784_;
wire _07785_;
wire _07786_;
wire _07787_;
wire _07788_;
wire _07789_;
wire _07790_;
wire _07791_;
wire _07792_;
wire _07793_;
wire _07794_;
wire _07795_;
wire _07796_;
wire _07797_;
wire _07798_;
wire _07799_;
wire _07800_;
wire _07801_;
wire _07802_;
wire _07803_;
wire _07804_;
wire _07805_;
wire _07806_;
wire _07807_;
wire _07808_;
wire _07809_;
wire _07810_;
wire _07811_;
wire _07812_;
wire _07813_;
wire _07814_;
wire _07815_;
wire _07816_;
wire _07817_;
wire _07818_;
wire _07819_;
wire _07820_;
wire _07821_;
wire _07822_;
wire _07823_;
wire _07824_;
wire _07825_;
wire _07826_;
wire _07827_;
wire _07828_;
wire _07829_;
wire _07830_;
wire _07831_;
wire _07832_;
wire _07833_;
wire _07834_;
wire _07835_;
wire _07836_;
wire _07837_;
wire _07838_;
wire _07839_;
wire _07840_;
wire _07841_;
wire _07842_;
wire _07843_;
wire _07844_;
wire _07845_;
wire _07846_;
wire _07847_;
wire _07848_;
wire _07849_;
wire _07850_;
wire _07851_;
wire _07852_;
wire _07853_;
wire _07854_;
wire _07855_;
wire _07856_;
wire _07857_;
wire _07858_;
wire _07859_;
wire _07860_;
wire _07861_;
wire _07862_;
wire _07863_;
wire _07864_;
wire _07865_;
wire _07866_;
wire _07867_;
wire _07868_;
wire _07869_;
wire _07870_;
wire _07871_;
wire _07872_;
wire _07873_;
wire _07874_;
wire _07875_;
wire _07876_;
wire _07877_;
wire _07878_;
wire _07879_;
wire _07880_;
wire _07881_;
wire _07882_;
wire _07883_;
wire _07884_;
wire _07885_;
wire _07886_;
wire _07887_;
wire _07888_;
wire _07889_;
wire _07890_;
wire _07891_;
wire _07892_;
wire _07893_;
wire _07894_;
wire _07895_;
wire _07896_;
wire _07897_;
wire _07898_;
wire _07899_;
wire _07900_;
wire _07901_;
wire _07902_;
wire _07903_;
wire _07904_;
wire _07905_;
wire _07906_;
wire _07907_;
wire _07908_;
wire _07909_;
wire _07910_;
wire _07911_;
wire _07912_;
wire _07913_;
wire _07914_;
wire _07915_;
wire _07916_;
wire _07917_;
wire _07918_;
wire _07919_;
wire _07920_;
wire _07921_;
wire _07922_;
wire _07923_;
wire _07924_;
wire _07925_;
wire _07926_;
wire _07927_;
wire _07928_;
wire _07929_;
wire _07930_;
wire _07931_;
wire _07932_;
wire _07933_;
wire _07934_;
wire _07935_;
wire _07936_;
wire _07937_;
wire _07938_;
wire _07939_;
wire _07940_;
wire _07941_;
wire _07942_;
wire _07943_;
wire _07944_;
wire _07945_;
wire _07946_;
wire _07947_;
wire _07948_;
wire _07949_;
wire _07950_;
wire _07951_;
wire _07952_;
wire _07953_;
wire _07954_;
wire _07955_;
wire _07956_;
wire _07957_;
wire _07958_;
wire _07959_;
wire _07960_;
wire _07961_;
wire _07962_;
wire _07963_;
wire _07964_;
wire _07965_;
wire _07966_;
wire _07967_;
wire _07968_;
wire _07969_;
wire _07970_;
wire _07971_;
wire _07972_;
wire _07973_;
wire _07974_;
wire _07975_;
wire _07976_;
wire _07977_;
wire _07978_;
wire _07979_;
wire _07980_;
wire _07981_;
wire _07982_;
wire _07983_;
wire _07984_;
wire _07985_;
wire _07986_;
wire _07987_;
wire _07988_;
wire _07989_;
wire _07990_;
wire _07991_;
wire _07992_;
wire _07993_;
wire _07994_;
wire _07995_;
wire _07996_;
wire _07997_;
wire _07998_;
wire _07999_;
wire _08000_;
wire _08001_;
wire _08002_;
wire _08003_;
wire _08004_;
wire _08005_;
wire _08006_;
wire _08007_;
wire _08008_;
wire _08009_;
wire _08010_;
wire _08011_;
wire _08012_;
wire _08013_;
wire _08014_;
wire _08015_;
wire _08016_;
wire _08017_;
wire _08018_;
wire _08019_;
wire _08020_;
wire _08021_;
wire _08022_;
wire _08023_;
wire _08024_;
wire _08025_;
wire _08026_;
wire _08027_;
wire _08028_;
wire _08029_;
wire _08030_;
wire _08031_;
wire _08032_;
wire _08033_;
wire _08034_;
wire _08035_;
wire _08036_;
wire _08037_;
wire _08038_;
wire _08039_;
wire _08040_;
wire _08041_;
wire _08042_;
wire _08043_;
wire _08044_;
wire _08045_;
wire _08046_;
wire _08047_;
wire _08048_;
wire _08049_;
wire _08050_;
wire _08051_;
wire _08052_;
wire _08053_;
wire _08054_;
wire _08055_;
wire _08056_;
wire _08057_;
wire _08058_;
wire _08059_;
wire _08060_;
wire _08061_;
wire _08062_;
wire _08063_;
wire _08064_;
wire _08065_;
wire _08066_;
wire _08067_;
wire _08068_;
wire _08069_;
wire _08070_;
wire _08071_;
wire _08072_;
wire _08073_;
wire _08074_;
wire _08075_;
wire _08076_;
wire _08077_;
wire _08078_;
wire _08079_;
wire _08080_;
wire _08081_;
wire _08082_;
wire _08083_;
wire _08084_;
wire _08085_;
wire _08086_;
wire _08087_;
wire _08088_;
wire _08089_;
wire _08090_;
wire _08091_;
wire _08092_;
wire _08093_;
wire _08094_;
wire _08095_;
wire _08096_;
wire _08097_;
wire _08098_;
wire _08099_;
wire _08100_;
wire _08101_;
wire _08102_;
wire _08103_;
wire _08104_;
wire _08105_;
wire _08106_;
wire _08107_;
wire _08108_;
wire _08109_;
wire _08110_;
wire _08111_;
wire _08112_;
wire _08113_;
wire _08114_;
wire _08115_;
wire _08116_;
wire _08117_;
wire _08118_;
wire _08119_;
wire _08120_;
wire _08121_;
wire _08122_;
wire _08123_;
wire _08124_;
wire _08125_;
wire _08126_;
wire _08127_;
wire _08128_;
wire _08129_;
wire _08130_;
wire _08131_;
wire _08132_;
wire _08133_;
wire _08134_;
wire _08135_;
wire _08136_;
wire _08137_;
wire _08138_;
wire _08139_;
wire _08140_;
wire _08141_;
wire _08142_;
wire _08143_;
wire _08144_;
wire _08145_;
wire _08146_;
wire _08147_;
wire _08148_;
wire _08149_;
wire _08150_;
wire _08151_;
wire _08152_;
wire _08153_;
wire _08154_;
wire _08155_;
wire _08156_;
wire _08157_;
wire _08158_;
wire _08159_;
wire _08160_;
wire _08161_;
wire _08162_;
wire _08163_;
wire _08164_;
wire _08165_;
wire _08166_;
wire _08167_;
wire _08168_;
wire _08169_;
wire _08170_;
wire _08171_;
wire _08172_;
wire _08173_;
wire _08174_;
wire _08175_;
wire _08176_;
wire _08177_;
wire _08178_;
wire _08179_;
wire _08180_;
wire _08181_;
wire _08182_;
wire _08183_;
wire _08184_;
wire _08185_;
wire _08186_;
wire _08187_;
wire _08188_;
wire _08189_;
wire _08190_;
wire _08191_;
wire _08192_;
wire _08193_;
wire _08194_;
wire _08195_;
wire _08196_;
wire _08197_;
wire _08198_;
wire _08199_;
wire _08200_;
wire _08201_;
wire _08202_;
wire _08203_;
wire _08204_;
wire _08205_;
wire _08206_;
wire _08207_;
wire _08208_;
wire _08209_;
wire _08210_;
wire _08211_;
wire _08212_;
wire _08213_;
wire _08214_;
wire _08215_;
wire _08216_;
wire _08217_;
wire _08218_;
wire _08219_;
wire _08220_;
wire _08221_;
wire _08222_;
wire _08223_;
wire _08224_;
wire _08225_;
wire _08226_;
wire _08227_;
wire _08228_;
wire _08229_;
wire _08230_;
wire _08231_;
wire _08232_;
wire _08233_;
wire _08234_;
wire _08235_;
wire _08236_;
wire _08237_;
wire _08238_;
wire _08239_;
wire _08240_;
wire _08241_;
wire _08242_;
wire _08243_;
wire _08244_;
wire _08245_;
wire _08246_;
wire _08247_;
wire _08248_;
wire _08249_;
wire _08250_;
wire _08251_;
wire _08252_;
wire _08253_;
wire _08254_;
wire _08255_;
wire _08256_;
wire _08257_;
wire _08258_;
wire _08259_;
wire _08260_;
wire _08261_;
wire _08262_;
wire _08263_;
wire _08264_;
wire _08265_;
wire _08266_;
wire _08267_;
wire _08268_;
wire _08269_;
wire _08270_;
wire _08271_;
wire _08272_;
wire _08273_;
wire _08274_;
wire _08275_;
wire _08276_;
wire _08277_;
wire _08278_;
wire _08279_;
wire _08280_;
wire _08281_;
wire _08282_;
wire _08283_;
wire _08284_;
wire _08285_;
wire _08286_;
wire _08287_;
wire _08288_;
wire _08289_;
wire _08290_;
wire _08291_;
wire _08292_;
wire _08293_;
wire _08294_;
wire _08295_;
wire _08296_;
wire _08297_;
wire _08298_;
wire _08299_;
wire _08300_;
wire _08301_;
wire _08302_;
wire _08303_;
wire _08304_;
wire _08305_;
wire _08306_;
wire _08307_;
wire _08308_;
wire _08309_;
wire _08310_;
wire _08311_;
wire _08312_;
wire _08313_;
wire _08314_;
wire _08315_;
wire _08316_;
wire _08317_;
wire _08318_;
wire _08319_;
wire _08320_;
wire _08321_;
wire _08322_;
wire _08323_;
wire _08324_;
wire _08325_;
wire _08326_;
wire _08327_;
wire _08328_;
wire _08329_;
wire _08330_;
wire _08331_;
wire _08332_;
wire _08333_;
wire _08334_;
wire _08335_;
wire _08336_;
wire _08337_;
wire _08338_;
wire _08339_;
wire _08340_;
wire _08341_;
wire _08342_;
wire _08343_;
wire _08344_;
wire _08345_;
wire _08346_;
wire _08347_;
wire _08348_;
wire _08349_;
wire _08350_;
wire _08351_;
wire _08352_;
wire _08353_;
wire _08354_;
wire _08355_;
wire _08356_;
wire _08357_;
wire _08358_;
wire _08359_;
wire _08360_;
wire _08361_;
wire _08362_;
wire _08363_;
wire _08364_;
wire _08365_;
wire _08366_;
wire _08367_;
wire _08368_;
wire _08369_;
wire _08370_;
wire _08371_;
wire _08372_;
wire _08373_;
wire _08374_;
wire _08375_;
wire _08376_;
wire _08377_;
wire _08378_;
wire _08379_;
wire _08380_;
wire _08381_;
wire _08382_;
wire _08383_;
wire _08384_;
wire _08385_;
wire _08386_;
wire _08387_;
wire _08388_;
wire _08389_;
wire _08390_;
wire _08391_;
wire _08392_;
wire _08393_;
wire _08394_;
wire _08395_;
wire _08396_;
wire _08397_;
wire _08398_;
wire _08399_;
wire _08400_;
wire _08401_;
wire _08402_;
wire _08403_;
wire _08404_;
wire _08405_;
wire _08406_;
wire _08407_;
wire _08408_;
wire _08409_;
wire _08410_;
wire _08411_;
wire _08412_;
wire _08413_;
wire _08414_;
wire _08415_;
wire _08416_;
wire _08417_;
wire _08418_;
wire _08419_;
wire _08420_;
wire _08421_;
wire _08422_;
wire _08423_;
wire _08424_;
wire _08425_;
wire _08426_;
wire _08427_;
wire _08428_;
wire _08429_;
wire _08430_;
wire _08431_;
wire _08432_;
wire _08433_;
wire _08434_;
wire _08435_;
wire _08436_;
wire _08437_;
wire _08438_;
wire _08439_;
wire _08440_;
wire _08441_;
wire _08442_;
wire _08443_;
wire _08444_;
wire _08445_;
wire _08446_;
wire _08447_;
wire _08448_;
wire _08449_;
wire _08450_;
wire _08451_;
wire _08452_;
wire _08453_;
wire _08454_;
wire _08455_;
wire _08456_;
wire _08457_;
wire _08458_;
wire _08459_;
wire _08460_;
wire _08461_;
wire _08462_;
wire _08463_;
wire _08464_;
wire _08465_;
wire _08466_;
wire _08467_;
wire _08468_;
wire _08469_;
wire _08470_;
wire _08471_;
wire _08472_;
wire _08473_;
wire _08474_;
wire _08475_;
wire _08476_;
wire _08477_;
wire _08478_;
wire _08479_;
wire _08480_;
wire _08481_;
wire _08482_;
wire _08483_;
wire _08484_;
wire _08485_;
wire _08486_;
wire _08487_;
wire _08488_;
wire _08489_;
wire _08490_;
wire _08491_;
wire _08492_;
wire _08493_;
wire _08494_;
wire _08495_;
wire _08496_;
wire _08497_;
wire _08498_;
wire _08499_;
wire _08500_;
wire _08501_;
wire _08502_;
wire _08503_;
wire _08504_;
wire _08505_;
wire _08506_;
wire _08507_;
wire _08508_;
wire _08509_;
wire _08510_;
wire _08511_;
wire _08512_;
wire _08513_;
wire _08514_;
wire _08515_;
wire _08516_;
wire _08517_;
wire _08518_;
wire _08519_;
wire _08520_;
wire _08521_;
wire _08522_;
wire _08523_;
wire _08524_;
wire _08525_;
wire _08526_;
wire _08527_;
wire _08528_;
wire _08529_;
wire _08530_;
wire _08531_;
wire _08532_;
wire _08533_;
wire _08534_;
wire _08535_;
wire _08536_;
wire _08537_;
wire _08538_;
wire _08539_;
wire _08540_;
wire _08541_;
wire _08542_;
wire _08543_;
wire _08544_;
wire _08545_;
wire _08546_;
wire _08547_;
wire _08548_;
wire _08549_;
wire _08550_;
wire _08551_;
wire _08552_;
wire _08553_;
wire _08554_;
wire _08555_;
wire _08556_;
wire _08557_;
wire _08558_;
wire _08559_;
wire _08560_;
wire _08561_;
wire _08562_;
wire _08563_;
wire _08564_;
wire _08565_;
wire _08566_;
wire _08567_;
wire _08568_;
wire _08569_;
wire _08570_;
wire _08571_;
wire _08572_;
wire _08573_;
wire _08574_;
wire _08575_;
wire _08576_;
wire _08577_;
wire _08578_;
wire _08579_;
wire _08580_;
wire _08581_;
wire _08582_;
wire _08583_;
wire _08584_;
wire _08585_;
wire _08586_;
wire _08587_;
wire _08588_;
wire _08589_;
wire _08590_;
wire _08591_;
wire _08592_;
wire _08593_;
wire _08594_;
wire _08595_;
wire _08596_;
wire _08597_;
wire _08598_;
wire _08599_;
wire _08600_;
wire _08601_;
wire _08602_;
wire _08603_;
wire _08604_;
wire _08605_;
wire _08606_;
wire _08607_;
wire _08608_;
wire _08609_;
wire _08610_;
wire _08611_;
wire _08612_;
wire _08613_;
wire _08614_;
wire _08615_;
wire _08616_;
wire _08617_;
wire _08618_;
wire _08619_;
wire _08620_;
wire _08621_;
wire _08622_;
wire _08623_;
wire _08624_;
wire _08625_;
wire _08626_;
wire _08627_;
wire _08628_;
wire _08629_;
wire _08630_;
wire _08631_;
wire _08632_;
wire _08633_;
wire _08634_;
wire _08635_;
wire _08636_;
wire _08637_;
wire _08638_;
wire _08639_;
wire _08640_;
wire _08641_;
wire _08642_;
wire _08643_;
wire _08644_;
wire _08645_;
wire _08646_;
wire _08647_;
wire _08648_;
wire _08649_;
wire _08650_;
wire _08651_;
wire _08652_;
wire _08653_;
wire _08654_;
wire _08655_;
wire _08656_;
wire _08657_;
wire _08658_;
wire _08659_;
wire _08660_;
wire _08661_;
wire _08662_;
wire _08663_;
wire _08664_;
wire _08665_;
wire _08666_;
wire _08667_;
wire _08668_;
wire _08669_;
wire _08670_;
wire _08671_;
wire _08672_;
wire _08673_;
wire _08674_;
wire _08675_;
wire _08676_;
wire _08677_;
wire _08678_;
wire _08679_;
wire _08680_;
wire _08681_;
wire _08682_;
wire _08683_;
wire _08684_;
wire _08685_;
wire _08686_;
wire _08687_;
wire _08688_;
wire _08689_;
wire _08690_;
wire _08691_;
wire _08692_;
wire _08693_;
wire _08694_;
wire _08695_;
wire _08696_;
wire _08697_;
wire _08698_;
wire _08699_;
wire _08700_;
wire _08701_;
wire _08702_;
wire _08703_;
wire _08704_;
wire _08705_;
wire _08706_;
wire _08707_;
wire _08708_;
wire _08709_;
wire _08710_;
wire _08711_;
wire _08712_;
wire _08713_;
wire _08714_;
wire _08715_;
wire _08716_;
wire _08717_;
wire _08718_;
wire _08719_;
wire _08720_;
wire _08721_;
wire _08722_;
wire _08723_;
wire _08724_;
wire _08725_;
wire _08726_;
wire _08727_;
wire _08728_;
wire _08729_;
wire _08730_;
wire _08731_;
wire _08732_;
wire _08733_;
wire _08734_;
wire _08735_;
wire _08736_;
wire _08737_;
wire _08738_;
wire _08739_;
wire _08740_;
wire _08741_;
wire _08742_;
wire _08743_;
wire _08744_;
wire _08745_;
wire _08746_;
wire _08747_;
wire _08748_;
wire _08749_;
wire _08750_;
wire _08751_;
wire _08752_;
wire _08753_;
wire _08754_;
wire _08755_;
wire _08756_;
wire _08757_;
wire _08758_;
wire _08759_;
wire _08760_;
wire _08761_;
wire _08762_;
wire _08763_;
wire _08764_;
wire _08765_;
wire _08766_;
wire _08767_;
wire _08768_;
wire _08769_;
wire _08770_;
wire _08771_;
wire _08772_;
wire _08773_;
wire _08774_;
wire _08775_;
wire _08776_;
wire _08777_;
wire _08778_;
wire _08779_;
wire _08780_;
wire _08781_;
wire _08782_;
wire _08783_;
wire _08784_;
wire _08785_;
wire _08786_;
wire _08787_;
wire _08788_;
wire _08789_;
wire _08790_;
wire _08791_;
wire _08792_;
wire _08793_;
wire _08794_;
wire _08795_;
wire _08796_;
wire _08797_;
wire _08798_;
wire _08799_;
wire _08800_;
wire _08801_;
wire _08802_;
wire _08803_;
wire _08804_;
wire _08805_;
wire _08806_;
wire _08807_;
wire _08808_;
wire _08809_;
wire _08810_;
wire _08811_;
wire _08812_;
wire _08813_;
wire _08814_;
wire _08815_;
wire _08816_;
wire _08817_;
wire _08818_;
wire _08819_;
wire _08820_;
wire _08821_;
wire _08822_;
wire _08823_;
wire _08824_;
wire _08825_;
wire _08826_;
wire _08827_;
wire _08828_;
wire _08829_;
wire _08830_;
wire _08831_;
wire _08832_;
wire _08833_;
wire _08834_;
wire _08835_;
wire _08836_;
wire _08837_;
wire _08838_;
wire _08839_;
wire _08840_;
wire _08841_;
wire _08842_;
wire _08843_;
wire _08844_;
wire _08845_;
wire _08846_;
wire _08847_;
wire _08848_;
wire _08849_;
wire _08850_;
wire _08851_;
wire _08852_;
wire _08853_;
wire _08854_;
wire _08855_;
wire _08856_;
wire _08857_;
wire _08858_;
wire _08859_;
wire _08860_;
wire _08861_;
wire _08862_;
wire _08863_;
wire _08864_;
wire _08865_;
wire _08866_;
wire _08867_;
wire _08868_;
wire _08869_;
wire _08870_;
wire _08871_;
wire _08872_;
wire _08873_;
wire _08874_;
wire _08875_;
wire _08876_;
wire _08877_;
wire _08878_;
wire _08879_;
wire _08880_;
wire _08881_;
wire _08882_;
wire _08883_;
wire _08884_;
wire _08885_;
wire _08886_;
wire _08887_;
wire _08888_;
wire _08889_;
wire _08890_;
wire _08891_;
wire _08892_;
wire _08893_;
wire _08894_;
wire _08895_;
wire _08896_;
wire _08897_;
wire _08898_;
wire _08899_;
wire _08900_;
wire _08901_;
wire _08902_;
wire _08903_;
wire _08904_;
wire _08905_;
wire _08906_;
wire _08907_;
wire _08908_;
wire _08909_;
wire _08910_;
wire _08911_;
wire _08912_;
wire _08913_;
wire _08914_;
wire _08915_;
wire _08916_;
wire _08917_;
wire _08918_;
wire _08919_;
wire _08920_;
wire _08921_;
wire _08922_;
wire _08923_;
wire _08924_;
wire _08925_;
wire _08926_;
wire _08927_;
wire _08928_;
wire _08929_;
wire _08930_;
wire _08931_;
wire _08932_;
wire _08933_;
wire _08934_;
wire _08935_;
wire _08936_;
wire _08937_;
wire _08938_;
wire _08939_;
wire _08940_;
wire _08941_;
wire _08942_;
wire _08943_;
wire _08944_;
wire _08945_;
wire _08946_;
wire _08947_;
wire _08948_;
wire _08949_;
wire _08950_;
wire _08951_;
wire _08952_;
wire _08953_;
wire _08954_;
wire _08955_;
wire _08956_;
wire _08957_;
wire _08958_;
wire _08959_;
wire _08960_;
wire _08961_;
wire _08962_;
wire _08963_;
wire _08964_;
wire _08965_;
wire _08966_;
wire _08967_;
wire _08968_;
wire _08969_;
wire _08970_;
wire _08971_;
wire _08972_;
wire _08973_;
wire _08974_;
wire _08975_;
wire _08976_;
wire _08977_;
wire _08978_;
wire _08979_;
wire _08980_;
wire _08981_;
wire _08982_;
wire _08983_;
wire _08984_;
wire _08985_;
wire _08986_;
wire _08987_;
wire _08988_;
wire _08989_;
wire _08990_;
wire _08991_;
wire _08992_;
wire _08993_;
wire _08994_;
wire _08995_;
wire _08996_;
wire _08997_;
wire _08998_;
wire _08999_;
wire _09000_;
wire _09001_;
wire _09002_;
wire _09003_;
wire _09004_;
wire _09005_;
wire _09006_;
wire _09007_;
wire _09008_;
wire _09009_;
wire _09010_;
wire _09011_;
wire _09012_;
wire _09013_;
wire _09014_;
wire _09015_;
wire _09016_;
wire _09017_;
wire _09018_;
wire _09019_;
wire _09020_;
wire _09021_;
wire _09022_;
wire _09023_;
wire _09024_;
wire _09025_;
wire _09026_;
wire _09027_;
wire _09028_;
wire _09029_;
wire _09030_;
wire _09031_;
wire _09032_;
wire _09033_;
wire _09034_;
wire _09035_;
wire _09036_;
wire _09037_;
wire _09038_;
wire _09039_;
wire _09040_;
wire _09041_;
wire _09042_;
wire _09043_;
wire _09044_;
wire _09045_;
wire _09046_;
wire _09047_;
wire _09048_;
wire _09049_;
wire _09050_;
wire _09051_;
wire _09052_;
wire _09053_;
wire _09054_;
wire _09055_;
wire _09056_;
wire _09057_;
wire _09058_;
wire _09059_;
wire _09060_;
wire _09061_;
wire _09062_;
wire _09063_;
wire _09064_;
wire _09065_;
wire _09066_;
wire _09067_;
wire _09068_;
wire _09069_;
wire _09070_;
wire _09071_;
wire _09072_;
wire _09073_;
wire _09074_;
wire _09075_;
wire _09076_;
wire _09077_;
wire _09078_;
wire _09079_;
wire _09080_;
wire _09081_;
wire _09082_;
wire _09083_;
wire _09084_;
wire _09085_;
wire _09086_;
wire _09087_;
wire _09088_;
wire _09089_;
wire _09090_;
wire _09091_;
wire _09092_;
wire _09093_;
wire _09094_;
wire _09095_;
wire _09096_;
wire _09097_;
wire _09098_;
wire _09099_;
wire _09100_;
wire _09101_;
wire _09102_;
wire _09103_;
wire _09104_;
wire _09105_;
wire _09106_;
wire _09107_;
wire _09108_;
wire _09109_;
wire _09110_;
wire _09111_;
wire _09112_;
wire _09113_;
wire _09114_;
wire _09115_;
wire _09116_;
wire _09117_;
wire _09118_;
wire _09119_;
wire _09120_;
wire _09121_;
wire _09122_;
wire _09123_;
wire _09124_;
wire _09125_;
wire _09126_;
wire _09127_;
wire _09128_;
wire _09129_;
wire _09130_;
wire _09131_;
wire _09132_;
wire _09133_;
wire _09134_;
wire _09135_;
wire _09136_;
wire _09137_;
wire _09138_;
wire _09139_;
wire _09140_;
wire _09141_;
wire _09142_;
wire _09143_;
wire _09144_;
wire _09145_;
wire _09146_;
wire _09147_;
wire _09148_;
wire _09149_;
wire _09150_;
wire _09151_;
wire _09152_;
wire _09153_;
wire _09154_;
wire _09155_;
wire _09156_;
wire _09157_;
wire _09158_;
wire _09159_;
wire _09160_;
wire _09161_;
wire _09162_;
wire _09163_;
wire _09164_;
wire _09165_;
wire _09166_;
wire _09167_;
wire _09168_;
wire _09169_;
wire _09170_;
wire _09171_;
wire _09172_;
wire _09173_;
wire _09174_;
wire _09175_;
wire _09176_;
wire _09177_;
wire _09178_;
wire _09179_;
wire _09180_;
wire _09181_;
wire _09182_;
wire _09183_;
wire _09184_;
wire _09185_;
wire _09186_;
wire _09187_;
wire _09188_;
wire _09189_;
wire _09190_;
wire _09191_;
wire _09192_;
wire _09193_;
wire _09194_;
wire _09195_;
wire _09196_;
wire _09197_;
wire _09198_;
wire _09199_;
wire _09200_;
wire _09201_;
wire _09202_;
wire _09203_;
wire _09204_;
wire _09205_;
wire _09206_;
wire _09207_;
wire _09208_;
wire _09209_;
wire _09210_;
wire _09211_;
wire _09212_;
wire _09213_;
wire _09214_;
wire _09215_;
wire _09216_;
wire _09217_;
wire _09218_;
wire _09219_;
wire _09220_;
wire _09221_;
wire _09222_;
wire _09223_;
wire _09224_;
wire _09225_;
wire _09226_;
wire _09227_;
wire _09228_;
wire _09229_;
wire _09230_;
wire _09231_;
wire _09232_;
wire _09233_;
wire _09234_;
wire _09235_;
wire _09236_;
wire _09237_;
wire _09238_;
wire _09239_;
wire _09240_;
wire _09241_;
wire _09242_;
wire _09243_;
wire _09244_;
wire _09245_;
wire _09246_;
wire _09247_;
wire _09248_;
wire _09249_;
wire _09250_;
wire _09251_;
wire _09252_;
wire _09253_;
wire _09254_;
wire _09255_;
wire _09256_;
wire _09257_;
wire _09258_;
wire _09259_;
wire _09260_;
wire _09261_;
wire _09262_;
wire _09263_;
wire _09264_;
wire _09265_;
wire _09266_;
wire _09267_;
wire _09268_;
wire _09269_;
wire _09270_;
wire _09271_;
wire _09272_;
wire _09273_;
wire _09274_;
wire _09275_;
wire _09276_;
wire _09277_;
wire _09278_;
wire _09279_;
wire _09280_;
wire _09281_;
wire _09282_;
wire _09283_;
wire _09284_;
wire _09285_;
wire _09286_;
wire _09287_;
wire _09288_;
wire _09289_;
wire _09290_;
wire _09291_;
wire _09292_;
wire _09293_;
wire _09294_;
wire _09295_;
wire _09296_;
wire _09297_;
wire _09298_;
wire _09299_;
wire _09300_;
wire _09301_;
wire _09302_;
wire _09303_;
wire _09304_;
wire _09305_;
wire _09306_;
wire _09307_;
wire _09308_;
wire _09309_;
wire _09310_;
wire _09311_;
wire _09312_;
wire _09313_;
wire _09314_;
wire _09315_;
wire _09316_;
wire _09317_;
wire _09318_;
wire _09319_;
wire _09320_;
wire _09321_;
wire _09322_;
wire _09323_;
wire _09324_;
wire _09325_;
wire _09326_;
wire _09327_;
wire _09328_;
wire _09329_;
wire _09330_;
wire _09331_;
wire _09332_;
wire _09333_;
wire _09334_;
wire _09335_;
wire _09336_;
wire _09337_;
wire _09338_;
wire _09339_;
wire _09340_;
wire _09341_;
wire _09342_;
wire _09343_;
wire _09344_;
wire _09345_;
wire _09346_;
wire _09347_;
wire _09348_;
wire _09349_;
wire _09350_;
wire _09351_;
wire _09352_;
wire _09353_;
wire _09354_;
wire _09355_;
wire _09356_;
wire _09357_;
wire _09358_;
wire _09359_;
wire _09360_;
wire _09361_;
wire _09362_;
wire _09363_;
wire _09364_;
wire _09365_;
wire _09366_;
wire _09367_;
wire _09368_;
wire _09369_;
wire _09370_;
wire _09371_;
wire _09372_;
wire _09373_;
wire _09374_;
wire _09375_;
wire _09376_;
wire _09377_;
wire _09378_;
wire _09379_;
wire _09380_;
wire _09381_;
wire _09382_;
wire _09383_;
wire _09384_;
wire _09385_;
wire _09386_;
wire _09387_;
wire _09388_;
wire _09389_;
wire _09390_;
wire _09391_;
wire _09392_;
wire _09393_;
wire _09394_;
wire _09395_;
wire _09396_;
wire _09397_;
wire _09398_;
wire _09399_;
wire _09400_;
wire _09401_;
wire _09402_;
wire _09403_;
wire _09404_;
wire _09405_;
wire _09406_;
wire _09407_;
wire _09408_;
wire _09409_;
wire _09410_;
wire _09411_;
wire _09412_;
wire _09413_;
wire _09414_;
wire _09415_;
wire _09416_;
wire _09417_;
wire _09418_;
wire _09419_;
wire _09420_;
wire _09421_;
wire _09422_;
wire _09423_;
wire _09424_;
wire _09425_;
wire _09426_;
wire _09427_;
wire _09428_;
wire _09429_;
wire _09430_;
wire _09431_;
wire _09432_;
wire _09433_;
wire _09434_;
wire _09435_;
wire _09436_;
wire _09437_;
wire _09438_;
wire _09439_;
wire _09440_;
wire _09441_;
wire _09442_;
wire _09443_;
wire _09444_;
wire _09445_;
wire _09446_;
wire _09447_;
wire _09448_;
wire _09449_;
wire _09450_;
wire _09451_;
wire _09452_;
wire _09453_;
wire _09454_;
wire _09455_;
wire _09456_;
wire _09457_;
wire _09458_;
wire _09459_;
wire _09460_;
wire _09461_;
wire _09462_;
wire _09463_;
wire _09464_;
wire _09465_;
wire _09466_;
wire _09467_;
wire _09468_;
wire _09469_;
wire _09470_;
wire _09471_;
wire _09472_;
wire _09473_;
wire _09474_;
wire _09475_;
wire _09476_;
wire _09477_;
wire _09478_;
wire _09479_;
wire _09480_;
wire _09481_;
wire _09482_;
wire _09483_;
wire _09484_;
wire _09485_;
wire _09486_;
wire _09487_;
wire _09488_;
wire _09489_;
wire _09490_;
wire _09491_;
wire _09492_;
wire _09493_;
wire _09494_;
wire _09495_;
wire _09496_;
wire _09497_;
wire _09498_;
wire _09499_;
wire _09500_;
wire _09501_;
wire _09502_;
wire _09503_;
wire _09504_;
wire _09505_;
wire _09506_;
wire _09507_;
wire _09508_;
wire _09509_;
wire _09510_;
wire _09511_;
wire _09512_;
wire _09513_;
wire _09514_;
wire _09515_;
wire _09516_;
wire _09517_;
wire _09518_;
wire _09519_;
wire _09520_;
wire _09521_;
wire _09522_;
wire _09523_;
wire _09524_;
wire _09525_;
wire _09526_;
wire _09527_;
wire _09528_;
wire _09529_;
wire _09530_;
wire _09531_;
wire _09532_;
wire _09533_;
wire _09534_;
wire _09535_;
wire _09536_;
wire _09537_;
wire _09538_;
wire _09539_;
wire _09540_;
wire _09541_;
wire _09542_;
wire _09543_;
wire _09544_;
wire _09545_;
wire _09546_;
wire _09547_;
wire _09548_;
wire _09549_;
wire _09550_;
wire _09551_;
wire _09552_;
wire _09553_;
wire _09554_;
wire _09555_;
wire _09556_;
wire _09557_;
wire _09558_;
wire _09559_;
wire _09560_;
wire _09561_;
wire _09562_;
wire _09563_;
wire _09564_;
wire _09565_;
wire _09566_;
wire _09567_;
wire _09568_;
wire _09569_;
wire _09570_;
wire _09571_;
wire _09572_;
wire _09573_;
wire _09574_;
wire _09575_;
wire _09576_;
wire _09577_;
wire _09578_;
wire _09579_;
wire _09580_;
wire _09581_;
wire _09582_;
wire _09583_;
wire _09584_;
wire _09585_;
wire _09586_;
wire _09587_;
wire _09588_;
wire _09589_;
wire _09590_;
wire _09591_;
wire _09592_;
wire _09593_;
wire _09594_;
wire _09595_;
wire _09596_;
wire _09597_;
wire _09598_;
wire _09599_;
wire _09600_;
wire _09601_;
wire _09602_;
wire _09603_;
wire _09604_;
wire _09605_;
wire _09606_;
wire _09607_;
wire _09608_;
wire _09609_;
wire _09610_;
wire _09611_;
wire _09612_;
wire _09613_;
wire _09614_;
wire _09615_;
wire _09616_;
wire _09617_;
wire _09618_;
wire _09619_;
wire _09620_;
wire _09621_;
wire _09622_;
wire _09623_;
wire _09624_;
wire _09625_;
wire _09626_;
wire _09627_;
wire _09628_;
wire _09629_;
wire _09630_;
wire _09631_;
wire _09632_;
wire _09633_;
wire _09634_;
wire _09635_;
wire _09636_;
wire _09637_;
wire _09638_;
wire _09639_;
wire _09640_;
wire _09641_;
wire _09642_;
wire _09643_;
wire _09644_;
wire _09645_;
wire _09646_;
wire _09647_;
wire _09648_;
wire _09649_;
wire _09650_;
wire _09651_;
wire _09652_;
wire _09653_;
wire _09654_;
wire _09655_;
wire _09656_;
wire _09657_;
wire _09658_;
wire _09659_;
wire _09660_;
wire _09661_;
wire _09662_;
wire _09663_;
wire _09664_;
wire _09665_;
wire _09666_;
wire _09667_;
wire _09668_;
wire _09669_;
wire _09670_;
wire _09671_;
wire _09672_;
wire _09673_;
wire _09674_;
wire _09675_;
wire _09676_;
wire _09677_;
wire _09678_;
wire _09679_;
wire _09680_;
wire _09681_;
wire _09682_;
wire _09683_;
wire _09684_;
wire _09685_;
wire _09686_;
wire _09687_;
wire _09688_;
wire _09689_;
wire _09690_;
wire _09691_;
wire _09692_;
wire _09693_;
wire _09694_;
wire _09695_;
wire _09696_;
wire _09697_;
wire _09698_;
wire _09699_;
wire _09700_;
wire _09701_;
wire _09702_;
wire _09703_;
wire _09704_;
wire _09705_;
wire _09706_;
wire _09707_;
wire _09708_;
wire _09709_;
wire _09710_;
wire _09711_;
wire _09712_;
wire _09713_;
wire _09714_;
wire _09715_;
wire _09716_;
wire _09717_;
wire _09718_;
wire _09719_;
wire _09720_;
wire _09721_;
wire _09722_;
wire _09723_;
wire _09724_;
wire _09725_;
wire _09726_;
wire _09727_;
wire _09728_;
wire _09729_;
wire _09730_;
wire _09731_;
wire _09732_;
wire _09733_;
wire _09734_;
wire _09735_;
wire _09736_;
wire _09737_;
wire _09738_;
wire _09739_;
wire _09740_;
wire _09741_;
wire _09742_;
wire _09743_;
wire _09744_;
wire _09745_;
wire _09746_;
wire _09747_;
wire _09748_;
wire _09749_;
wire _09750_;
wire _09751_;
wire _09752_;
wire _09753_;
wire _09754_;
wire _09755_;
wire _09756_;
wire _09757_;
wire _09758_;
wire _09759_;
wire _09760_;
wire _09761_;
wire _09762_;
wire _09763_;
wire _09764_;
wire _09765_;
wire _09766_;
wire _09767_;
wire _09768_;
wire _09769_;
wire _09770_;
wire _09771_;
wire _09772_;
wire _09773_;
wire _09774_;
wire _09775_;
wire _09776_;
wire _09777_;
wire _09778_;
wire _09779_;
wire _09780_;
wire _09781_;
wire _09782_;
wire _09783_;
wire _09784_;
wire _09785_;
wire _09786_;
wire _09787_;
wire _09788_;
wire _09789_;
wire _09790_;
wire _09791_;
wire _09792_;
wire _09793_;
wire _09794_;
wire _09795_;
wire _09796_;
wire _09797_;
wire _09798_;
wire _09799_;
wire _09800_;
wire _09801_;
wire _09802_;
wire _09803_;
wire _09804_;
wire _09805_;
wire _09806_;
wire _09807_;
wire _09808_;
wire _09809_;
wire _09810_;
wire _09811_;
wire _09812_;
wire _09813_;
wire _09814_;
wire _09815_;
wire _09816_;
wire _09817_;
wire _09818_;
wire _09819_;
wire _09820_;
wire _09821_;
wire _09822_;
wire _09823_;
wire _09824_;
wire _09825_;
wire _09826_;
wire _09827_;
wire _09828_;
wire _09829_;
wire _09830_;
wire _09831_;
wire _09832_;
wire _09833_;
wire _09834_;
wire _09835_;
wire _09836_;
wire _09837_;
wire _09838_;
wire _09839_;
wire _09840_;
wire _09841_;
wire _09842_;
wire _09843_;
wire _09844_;
wire _09845_;
wire _09846_;
wire _09847_;
wire _09848_;
wire _09849_;
wire _09850_;
wire _09851_;
wire _09852_;
wire _09853_;
wire _09854_;
wire _09855_;
wire _09856_;
wire _09857_;
wire _09858_;
wire _09859_;
wire _09860_;
wire _09861_;
wire _09862_;
wire _09863_;
wire _09864_;
wire _09865_;
wire _09866_;
wire _09867_;
wire _09868_;
wire _09869_;
wire _09870_;
wire _09871_;
wire _09872_;
wire _09873_;
wire _09874_;
wire _09875_;
wire _09876_;
wire _09877_;
wire _09878_;
wire _09879_;
wire _09880_;
wire _09881_;
wire _09882_;
wire _09883_;
wire _09884_;
wire _09885_;
wire _09886_;
wire _09887_;
wire _09888_;
wire _09889_;
wire _09890_;
wire _09891_;
wire _09892_;
wire _09893_;
wire _09894_;
wire _09895_;
wire _09896_;
wire _09897_;
wire _09898_;
wire _09899_;
wire _09900_;
wire _09901_;
wire _09902_;
wire _09903_;
wire _09904_;
wire _09905_;
wire _09906_;
wire _09907_;
wire _09908_;
wire _09909_;
wire _09910_;
wire _09911_;
wire _09912_;
wire _09913_;
wire _09914_;
wire _09915_;
wire _09916_;
wire _09917_;
wire _09918_;
wire _09919_;
wire _09920_;
wire _09921_;
wire _09922_;
wire _09923_;
wire _09924_;
wire _09925_;
wire _09926_;
wire _09927_;
wire _09928_;
wire _09929_;
wire _09930_;
wire _09931_;
wire _09932_;
wire _09933_;
wire _09934_;
wire _09935_;
wire _09936_;
wire _09937_;
wire _09938_;
wire _09939_;
wire _09940_;
wire _09941_;
wire _09942_;
wire _09943_;
wire _09944_;
wire _09945_;
wire _09946_;
wire _09947_;
wire _09948_;
wire _09949_;
wire _09950_;
wire _09951_;
wire _09952_;
wire _09953_;
wire _09954_;
wire _09955_;
wire _09956_;
wire _09957_;
wire _09958_;
wire _09959_;
wire _09960_;
wire _09961_;
wire _09962_;
wire _09963_;
wire _09964_;
wire _09965_;
wire _09966_;
wire _09967_;
wire _09968_;
wire _09969_;
wire _09970_;
wire _09971_;
wire _09972_;
wire _09973_;
wire _09974_;
wire _09975_;
wire _09976_;
wire _09977_;
wire _09978_;
wire _09979_;
wire _09980_;
wire _09981_;
wire _09982_;
wire _09983_;
wire _09984_;
wire _09985_;
wire _09986_;
wire _09987_;
wire _09988_;
wire _09989_;
wire _09990_;
wire _09991_;
wire _09992_;
wire _09993_;
wire _09994_;
wire _09995_;
wire _09996_;
wire _09997_;
wire _09998_;
wire _09999_;
wire _10000_;
wire _10001_;
wire _10002_;
wire _10003_;
wire _10004_;
wire _10005_;
wire _10006_;
wire _10007_;
wire _10008_;
wire _10009_;
wire _10010_;
wire _10011_;
wire _10012_;
wire _10013_;
wire _10014_;
wire _10015_;
wire _10016_;
wire _10017_;
wire _10018_;
wire _10019_;
wire _10020_;
wire _10021_;
wire _10022_;
wire _10023_;
wire _10024_;
wire _10025_;
wire _10026_;
wire _10027_;
wire _10028_;
wire _10029_;
wire _10030_;
wire _10031_;
wire _10032_;
wire _10033_;
wire _10034_;
wire _10035_;
wire _10036_;
wire _10037_;
wire _10038_;
wire _10039_;
wire _10040_;
wire _10041_;
wire _10042_;
wire _10043_;
wire _10044_;
wire _10045_;
wire _10046_;
wire _10047_;
wire _10048_;
wire _10049_;
wire _10050_;
wire _10051_;
wire _10052_;
wire _10053_;
wire _10054_;
wire _10055_;
wire _10056_;
wire _10057_;
wire _10058_;
wire _10059_;
wire _10060_;
wire _10061_;
wire _10062_;
wire _10063_;
wire _10064_;
wire _10065_;
wire _10066_;
wire _10067_;
wire _10068_;
wire _10069_;
wire _10070_;
wire _10071_;
wire _10072_;
wire _10073_;
wire _10074_;
wire _10075_;
wire _10076_;
wire _10077_;
wire _10078_;
wire _10079_;
wire _10080_;
wire _10081_;
wire _10082_;
wire _10083_;
wire _10084_;
wire _10085_;
wire _10086_;
wire _10087_;
wire _10088_;
wire _10089_;
wire _10090_;
wire _10091_;
wire _10092_;
wire _10093_;
wire _10094_;
wire _10095_;
wire _10096_;
wire _10097_;
wire _10098_;
wire _10099_;
wire _10100_;
wire _10101_;
wire _10102_;
wire _10103_;
wire _10104_;
wire _10105_;
wire _10106_;
wire _10107_;
wire _10108_;
wire _10109_;
wire _10110_;
wire _10111_;
wire _10112_;
wire _10113_;
wire _10114_;
wire _10115_;
wire _10116_;
wire _10117_;
wire _10118_;
wire _10119_;
wire _10120_;
wire _10121_;
wire _10122_;
wire _10123_;
wire _10124_;
wire _10125_;
wire _10126_;
wire _10127_;
wire _10128_;
wire _10129_;
wire _10130_;
wire _10131_;
wire _10132_;
wire _10133_;
wire _10134_;
wire _10135_;
wire _10136_;
wire _10137_;
wire _10138_;
wire _10139_;
wire _10140_;
wire _10141_;
wire _10142_;
wire _10143_;
wire _10144_;
wire _10145_;
wire _10146_;
wire _10147_;
wire _10148_;
wire _10149_;
wire _10150_;
wire _10151_;
wire _10152_;
wire _10153_;
wire _10154_;
wire _10155_;
wire _10156_;
wire _10157_;
wire _10158_;
wire _10159_;
wire _10160_;
wire _10161_;
wire _10162_;
wire _10163_;
wire _10164_;
wire _10165_;
wire _10166_;
wire _10167_;
wire _10168_;
wire _10169_;
wire _10170_;
wire _10171_;
wire _10172_;
wire _10173_;
wire _10174_;
wire _10175_;
wire _10176_;
wire _10177_;
wire _10178_;
wire _10179_;
wire _10180_;
wire _10181_;
wire _10182_;
wire _10183_;
wire _10184_;
wire _10185_;
wire _10186_;
wire _10187_;
wire _10188_;
wire _10189_;
wire _10190_;
wire _10191_;
wire _10192_;
wire _10193_;
wire _10194_;
wire _10195_;
wire _10196_;
wire _10197_;
wire _10198_;
wire _10199_;
wire _10200_;
wire _10201_;
wire _10202_;
wire _10203_;
wire _10204_;
wire _10205_;
wire _10206_;
wire _10207_;
wire _10208_;
wire _10209_;
wire _10210_;
wire _10211_;
wire _10212_;
wire _10213_;
wire _10214_;
wire _10215_;
wire _10216_;
wire _10217_;
wire _10218_;
wire _10219_;
wire _10220_;
wire _10221_;
wire _10222_;
wire _10223_;
wire _10224_;
wire _10225_;
wire _10226_;
wire _10227_;
wire _10228_;
wire _10229_;
wire _10230_;
wire _10231_;
wire _10232_;
wire _10233_;
wire _10234_;
wire _10235_;
wire _10236_;
wire _10237_;
wire _10238_;
wire _10239_;
wire _10240_;
wire _10241_;
wire _10242_;
wire _10243_;
wire _10244_;
wire _10245_;
wire _10246_;
wire _10247_;
wire _10248_;
wire _10249_;
wire _10250_;
wire _10251_;
wire _10252_;
wire _10253_;
wire _10254_;
wire _10255_;
wire _10256_;
wire _10257_;
wire _10258_;
wire _10259_;
wire _10260_;
wire _10261_;
wire _10262_;
wire _10263_;
wire _10264_;
wire _10265_;
wire _10266_;
wire _10267_;
wire _10268_;
wire _10269_;
wire _10270_;
wire _10271_;
wire _10272_;
wire _10273_;
wire _10274_;
wire _10275_;
wire _10276_;
wire _10277_;
wire _10278_;
wire _10279_;
wire _10280_;
wire _10281_;
wire _10282_;
wire _10283_;
wire _10284_;
wire _10285_;
wire _10286_;
wire _10287_;
wire _10288_;
wire _10289_;
wire _10290_;
wire _10291_;
wire _10292_;
wire _10293_;
wire _10294_;
wire _10295_;
wire _10296_;
wire _10297_;
wire _10298_;
wire _10299_;
wire _10300_;
wire _10301_;
wire _10302_;
wire _10303_;
wire _10304_;
wire _10305_;
wire _10306_;
wire _10307_;
wire _10308_;
wire _10309_;
wire _10310_;
wire _10311_;
wire _10312_;
wire _10313_;
wire _10314_;
wire _10315_;
wire _10316_;
wire _10317_;
wire _10318_;
wire _10319_;
wire _10320_;
wire _10321_;
wire _10322_;
wire _10323_;
wire _10324_;
wire _10325_;
wire _10326_;
wire _10327_;
wire _10328_;
wire _10329_;
wire _10330_;
wire _10331_;
wire _10332_;
wire _10333_;
wire _10334_;
wire _10335_;
wire _10336_;
wire _10337_;
wire _10338_;
wire _10339_;
wire _10340_;
wire _10341_;
wire _10342_;
wire _10343_;
wire _10344_;
wire _10345_;
wire _10346_;
wire _10347_;
wire _10348_;
wire _10349_;
wire _10350_;
wire _10351_;
wire _10352_;
wire _10353_;
wire _10354_;
wire _10355_;
wire _10356_;
wire _10357_;
wire _10358_;
wire _10359_;
wire _10360_;
wire _10361_;
wire _10362_;
wire _10363_;
wire _10364_;
wire _10365_;
wire _10366_;
wire _10367_;
wire _10368_;
wire _10369_;
wire _10370_;
wire _10371_;
wire _10372_;
wire _10373_;
wire _10374_;
wire _10375_;
wire _10376_;
wire _10377_;
wire _10378_;
wire _10379_;
wire _10380_;
wire _10381_;
wire _10382_;
wire _10383_;
wire _10384_;
wire _10385_;
wire _10386_;
wire _10387_;
wire _10388_;
wire _10389_;
wire _10390_;
wire _10391_;
wire _10392_;
wire _10393_;
wire _10394_;
wire _10395_;
wire _10396_;
wire _10397_;
wire _10398_;
wire _10399_;
wire _10400_;
wire _10401_;
wire _10402_;
wire _10403_;
wire _10404_;
wire _10405_;
wire _10406_;
wire _10407_;
wire _10408_;
wire _10409_;
wire _10410_;
wire _10411_;
wire _10412_;
wire _10413_;
wire _10414_;
wire _10415_;
wire _10416_;
wire _10417_;
wire _10418_;
wire _10419_;
wire _10420_;
wire _10421_;
wire _10422_;
wire _10423_;
wire _10424_;
wire _10425_;
wire _10426_;
wire _10427_;
wire _10428_;
wire _10429_;
wire _10430_;
wire _10431_;
wire _10432_;
wire _10433_;
wire _10434_;
wire _10435_;
wire _10436_;
wire _10437_;
wire _10438_;
wire _10439_;
wire _10440_;
wire _10441_;
wire _10442_;
wire _10443_;
wire _10444_;
wire _10445_;
wire _10446_;
wire _10447_;
wire _10448_;
wire _10449_;
wire _10450_;
wire _10451_;
wire _10452_;
wire _10453_;
wire _10454_;
wire _10455_;
wire _10456_;
wire _10457_;
wire _10458_;
wire _10459_;
wire _10460_;
wire _10461_;
wire _10462_;
wire _10463_;
wire _10464_;
wire _10465_;
wire _10466_;
wire _10467_;
wire _10468_;
wire _10469_;
wire _10470_;
wire _10471_;
wire _10472_;
wire _10473_;
wire _10474_;
wire _10475_;
wire _10476_;
wire _10477_;
wire _10478_;
wire _10479_;
wire _10480_;
wire _10481_;
wire _10482_;
wire _10483_;
wire _10484_;
wire _10485_;
wire _10486_;
wire _10487_;
wire _10488_;
wire _10489_;
wire _10490_;
wire _10491_;
wire _10492_;
wire _10493_;
wire _10494_;
wire _10495_;
wire _10496_;
wire _10497_;
wire _10498_;
wire _10499_;
wire _10500_;
wire _10501_;
wire _10502_;
wire _10503_;
wire _10504_;
wire _10505_;
wire _10506_;
wire _10507_;
wire _10508_;
wire _10509_;
wire _10510_;
wire _10511_;
wire _10512_;
wire _10513_;
wire _10514_;
wire _10515_;
wire _10516_;
wire _10517_;
wire _10518_;
wire _10519_;
wire _10520_;
wire _10521_;
wire _10522_;
wire _10523_;
wire _10524_;
wire _10525_;
wire _10526_;
wire _10527_;
wire _10528_;
wire _10529_;
wire _10530_;
wire _10531_;
wire _10532_;
wire _10533_;
wire _10534_;
wire _10535_;
wire _10536_;
wire _10537_;
wire _10538_;
wire _10539_;
wire _10540_;
wire _10541_;
wire _10542_;
wire _10543_;
wire _10544_;
wire _10545_;
wire _10546_;
wire _10547_;
wire _10548_;
wire _10549_;
wire _10550_;
wire _10551_;
wire _10552_;
wire _10553_;
wire _10554_;
wire _10555_;
wire _10556_;
wire _10557_;
wire _10558_;
wire _10559_;
wire _10560_;
wire _10561_;
wire _10562_;
wire _10563_;
wire _10564_;
wire _10565_;
wire _10566_;
wire _10567_;
wire _10568_;
wire _10569_;
wire _10570_;
wire _10571_;
wire _10572_;
wire _10573_;
wire _10574_;
wire _10575_;
wire _10576_;
wire _10577_;
wire _10578_;
wire _10579_;
wire _10580_;
wire _10581_;
wire _10582_;
wire _10583_;
wire _10584_;
wire _10585_;
wire _10586_;
wire _10587_;
wire _10588_;
wire _10589_;
wire _10590_;
wire _10591_;
wire _10592_;
wire _10593_;
wire _10594_;
wire _10595_;
wire _10596_;
wire _10597_;
wire _10598_;
wire _10599_;
wire _10600_;
wire _10601_;
wire _10602_;
wire _10603_;
wire _10604_;
wire _10605_;
wire _10606_;
wire _10607_;
wire _10608_;
wire _10609_;
wire _10610_;
wire _10611_;
wire _10612_;
wire _10613_;
wire _10614_;
wire _10615_;
wire _10616_;
wire _10617_;
wire _10618_;
wire _10619_;
wire _10620_;
wire _10621_;
wire _10622_;
wire _10623_;
wire _10624_;
wire _10625_;
wire _10626_;
wire _10627_;
wire _10628_;
wire _10629_;
wire _10630_;
wire _10631_;
wire _10632_;
wire _10633_;
wire _10634_;
wire _10635_;
wire _10636_;
wire _10637_;
wire _10638_;
wire _10639_;
wire _10640_;
wire _10641_;
wire _10642_;
wire _10643_;
wire _10644_;
wire _10645_;
wire _10646_;
wire _10647_;
wire _10648_;
wire _10649_;
wire _10650_;
wire _10651_;
wire _10652_;
wire _10653_;
wire _10654_;
wire _10655_;
wire _10656_;
wire _10657_;
wire _10658_;
wire _10659_;
wire _10660_;
wire _10661_;
wire _10662_;
wire _10663_;
wire _10664_;
wire _10665_;
wire _10666_;
wire _10667_;
wire _10668_;
wire _10669_;
wire _10670_;
wire _10671_;
wire _10672_;
wire _10673_;
wire _10674_;
wire _10675_;
wire _10676_;
wire _10677_;
wire _10678_;
wire _10679_;
wire _10680_;
wire _10681_;
wire _10682_;
wire _10683_;
wire _10684_;
wire _10685_;
wire _10686_;
wire _10687_;
wire _10688_;
wire _10689_;
wire _10690_;
wire _10691_;
wire _10692_;
wire _10693_;
wire _10694_;
wire _10695_;
wire _10696_;
wire _10697_;
wire _10698_;
wire _10699_;
wire _10700_;
wire _10701_;
wire _10702_;
wire _10703_;
wire _10704_;
wire _10705_;
wire _10706_;
wire _10707_;
wire _10708_;
wire _10709_;
wire _10710_;
wire _10711_;
wire _10712_;
wire _10713_;
wire _10714_;
wire _10715_;
wire _10716_;
wire _10717_;
wire _10718_;
wire _10719_;
wire _10720_;
wire _10721_;
wire _10722_;
wire _10723_;
wire _10724_;
wire _10725_;
wire _10726_;
wire _10727_;
wire _10728_;
wire _10729_;
wire _10730_;
wire _10731_;
wire _10732_;
wire _10733_;
wire _10734_;
wire _10735_;
wire _10736_;
wire _10737_;
wire _10738_;
wire _10739_;
wire _10740_;
wire _10741_;
wire _10742_;
wire _10743_;
wire _10744_;
wire _10745_;
wire _10746_;
wire _10747_;
wire _10748_;
wire _10749_;
wire _10750_;
wire _10751_;
wire _10752_;
wire _10753_;
wire _10754_;
wire _10755_;
wire _10756_;
wire _10757_;
wire _10758_;
wire _10759_;
wire _10760_;
wire _10761_;
wire _10762_;
wire _10763_;
wire _10764_;
wire _10765_;
wire _10766_;
wire _10767_;
wire _10768_;
wire _10769_;
wire _10770_;
wire _10771_;
wire _10772_;
wire _10773_;
wire _10774_;
wire _10775_;
wire _10776_;
wire _10777_;
wire _10778_;
wire _10779_;
wire _10780_;
wire _10781_;
wire _10782_;
wire _10783_;
wire _10784_;
wire _10785_;
wire _10786_;
wire _10787_;
wire _10788_;
wire _10789_;
wire _10790_;
wire _10791_;
wire _10792_;
wire _10793_;
wire _10794_;
wire _10795_;
wire _10796_;
wire _10797_;
wire _10798_;
wire _10799_;
wire _10800_;
wire _10801_;
wire _10802_;
wire _10803_;
wire _10804_;
wire _10805_;
wire _10806_;
wire _10807_;
wire _10808_;
wire _10809_;
wire _10810_;
wire _10811_;
wire _10812_;
wire _10813_;
wire _10814_;
wire _10815_;
wire _10816_;
wire _10817_;
wire _10818_;
wire _10819_;
wire _10820_;
wire _10821_;
wire _10822_;
wire _10823_;
wire _10824_;
wire _10825_;
wire _10826_;
wire _10827_;
wire _10828_;
wire _10829_;
wire _10830_;
wire _10831_;
wire _10832_;
wire _10833_;
wire _10834_;
wire _10835_;
wire _10836_;
wire _10837_;
wire _10838_;
wire _10839_;
wire _10840_;
wire _10841_;
wire _10842_;
wire _10843_;
wire _10844_;
wire _10845_;
wire _10846_;
wire _10847_;
wire _10848_;
wire _10849_;
wire _10850_;
wire _10851_;
wire _10852_;
wire _10853_;
wire _10854_;
wire _10855_;
wire _10856_;
wire _10857_;
wire _10858_;
wire _10859_;
wire _10860_;
wire _10861_;
wire _10862_;
wire _10863_;
wire _10864_;
wire _10865_;
wire _10866_;
wire _10867_;
wire _10868_;
wire _10869_;
wire _10870_;
wire _10871_;
wire _10872_;
wire _10873_;
wire _10874_;
wire _10875_;
wire _10876_;
wire _10877_;
wire _10878_;
wire _10879_;
wire _10880_;
wire _10881_;
wire _10882_;
wire _10883_;
wire _10884_;
wire _10885_;
wire _10886_;
wire _10887_;
wire _10888_;
wire _10889_;
wire _10890_;
wire _10891_;
wire _10892_;
wire _10893_;
wire _10894_;
wire _10895_;
wire _10896_;
wire _10897_;
wire _10898_;
wire _10899_;
wire _10900_;
wire _10901_;
wire _10902_;
wire _10903_;
wire _10904_;
wire _10905_;
wire _10906_;
wire _10907_;
wire _10908_;
wire _10909_;
wire _10910_;
wire _10911_;
wire _10912_;
wire _10913_;
wire _10914_;
wire _10915_;
wire _10916_;
wire _10917_;
wire _10918_;
wire _10919_;
wire _10920_;
wire _10921_;
wire _10922_;
wire _10923_;
wire _10924_;
wire _10925_;
wire _10926_;
wire _10927_;
wire _10928_;
wire _10929_;
wire _10930_;
wire _10931_;
wire _10932_;
wire _10933_;
wire _10934_;
wire _10935_;
wire _10936_;
wire _10937_;
wire _10938_;
wire _10939_;
wire _10940_;
wire _10941_;
wire _10942_;
wire _10943_;
wire _10944_;
wire _10945_;
wire _10946_;
wire _10947_;
wire _10948_;
wire _10949_;
wire _10950_;
wire _10951_;
wire _10952_;
wire _10953_;
wire _10954_;
wire _10955_;
wire _10956_;
wire _10957_;
wire _10958_;
wire _10959_;
wire _10960_;
wire _10961_;
wire _10962_;
wire _10963_;
wire _10964_;
wire _10965_;
wire _10966_;
wire _10967_;
wire _10968_;
wire _10969_;
wire _10970_;
wire _10971_;
wire _10972_;
wire _10973_;
wire _10974_;
wire _10975_;
wire _10976_;
wire _10977_;
wire _10978_;
wire _10979_;
wire _10980_;
wire _10981_;
wire _10982_;
wire _10983_;
wire _10984_;
wire _10985_;
wire _10986_;
wire _10987_;
wire _10988_;
wire _10989_;
wire _10990_;
wire _10991_;
wire _10992_;
wire _10993_;
wire _10994_;
wire _10995_;
wire _10996_;
wire _10997_;
wire _10998_;
wire _10999_;
wire _11000_;
wire _11001_;
wire _11002_;
wire _11003_;
wire _11004_;
wire _11005_;
wire _11006_;
wire _11007_;
wire _11008_;
wire _11009_;
wire _11010_;
wire _11011_;
wire _11012_;
wire _11013_;
wire _11014_;
wire _11015_;
wire _11016_;
wire _11017_;
wire _11018_;
wire _11019_;
wire _11020_;
wire _11021_;
wire _11022_;
wire _11023_;
wire _11024_;
wire _11025_;
wire _11026_;
wire _11027_;
wire _11028_;
wire _11029_;
wire _11030_;
wire _11031_;
wire _11032_;
wire _11033_;
wire _11034_;
wire _11035_;
wire _11036_;
wire _11037_;
wire _11038_;
wire _11039_;
wire _11040_;
wire _11041_;
wire _11042_;
wire _11043_;
wire _11044_;
wire _11045_;
wire _11046_;
wire _11047_;
wire _11048_;
wire _11049_;
wire _11050_;
wire _11051_;
wire _11052_;
wire _11053_;
wire _11054_;
wire _11055_;
wire _11056_;
wire _11057_;
wire _11058_;
wire _11059_;
wire _11060_;
wire _11061_;
wire _11062_;
wire _11063_;
wire _11064_;
wire _11065_;
wire _11066_;
wire _11067_;
wire _11068_;
wire _11069_;
wire _11070_;
wire _11071_;
wire _11072_;
wire _11073_;
wire _11074_;
wire _11075_;
wire _11076_;
wire _11077_;
wire _11078_;
wire _11079_;
wire _11080_;
wire _11081_;
wire _11082_;
wire _11083_;
wire _11084_;
wire _11085_;
wire _11086_;
wire _11087_;
wire _11088_;
wire _11089_;
wire _11090_;
wire _11091_;
wire _11092_;
wire _11093_;
wire _11094_;
wire _11095_;
wire _11096_;
wire _11097_;
wire _11098_;
wire _11099_;
wire _11100_;
wire _11101_;
wire _11102_;
wire _11103_;
wire _11104_;
wire _11105_;
wire _11106_;
wire _11107_;
wire _11108_;
wire _11109_;
wire _11110_;
wire _11111_;
wire _11112_;
wire _11113_;
wire _11114_;
wire _11115_;
wire _11116_;
wire _11117_;
wire _11118_;
wire _11119_;
wire _11120_;
wire _11121_;
wire _11122_;
wire _11123_;
wire _11124_;
wire _11125_;
wire _11126_;
wire _11127_;
wire _11128_;
wire _11129_;
wire _11130_;
wire _11131_;
wire _11132_;
wire _11133_;
wire _11134_;
wire _11135_;
wire _11136_;
wire _11137_;
wire _11138_;
wire _11139_;
wire _11140_;
wire _11141_;
wire _11142_;
wire _11143_;
wire _11144_;
wire _11145_;
wire _11146_;
wire _11147_;
wire _11148_;
wire _11149_;
wire _11150_;
wire _11151_;
wire _11152_;
wire _11153_;
wire _11154_;
wire _11155_;
wire _11156_;
wire _11157_;
wire _11158_;
wire _11159_;
wire _11160_;
wire _11161_;
wire _11162_;
wire _11163_;
wire _11164_;
wire _11165_;
wire _11166_;
wire _11167_;
wire _11168_;
wire _11169_;
wire _11170_;
wire _11171_;
wire _11172_;
wire _11173_;
wire _11174_;
wire _11175_;
wire _11176_;
wire _11177_;
wire _11178_;
wire _11179_;
wire _11180_;
wire _11181_;
wire _11182_;
wire _11183_;
wire _11184_;
wire _11185_;
wire _11186_;
wire _11187_;
wire _11188_;
wire _11189_;
wire _11190_;
wire _11191_;
wire _11192_;
wire _11193_;
wire _11194_;
wire _11195_;
wire _11196_;
wire _11197_;
wire _11198_;
wire _11199_;
wire _11200_;
wire _11201_;
wire _11202_;
wire _11203_;
wire _11204_;
wire _11205_;
wire _11206_;
wire _11207_;
wire _11208_;
wire _11209_;
wire _11210_;
wire _11211_;
wire _11212_;
wire _11213_;
wire _11214_;
wire _11215_;
wire _11216_;
wire _11217_;
wire _11218_;
wire _11219_;
wire _11220_;
wire _11221_;
wire _11222_;
wire _11223_;
wire _11224_;
wire _11225_;
wire _11226_;
wire _11227_;
wire _11228_;
wire _11229_;
wire _11230_;
wire _11231_;
wire _11232_;
wire _11233_;
wire _11234_;
wire _11235_;
wire _11236_;
wire _11237_;
wire _11238_;
wire _11239_;
wire _11240_;
wire _11241_;
wire _11242_;
wire _11243_;
wire _11244_;
wire _11245_;
wire _11246_;
wire _11247_;
wire _11248_;
wire _11249_;
wire _11250_;
wire _11251_;
wire _11252_;
wire _11253_;
wire _11254_;
wire _11255_;
wire _11256_;
wire _11257_;
wire _11258_;
wire _11259_;
wire _11260_;
wire _11261_;
wire _11262_;
wire _11263_;
wire _11264_;
wire _11265_;
wire _11266_;
wire _11267_;
wire _11268_;
wire _11269_;
wire _11270_;
wire _11271_;
wire _11272_;
wire _11273_;
wire _11274_;
wire _11275_;
wire _11276_;
wire _11277_;
wire _11278_;
wire _11279_;
wire _11280_;
wire _11281_;
wire _11282_;
wire _11283_;
wire _11284_;
wire _11285_;
wire _11286_;
wire _11287_;
wire _11288_;
wire _11289_;
wire _11290_;
wire _11291_;
wire _11292_;
wire _11293_;
wire _11294_;
wire _11295_;
wire _11296_;
wire _11297_;
wire _11298_;
wire _11299_;
wire _11300_;
wire _11301_;
wire _11302_;
wire _11303_;
wire _11304_;
wire _11305_;
wire _11306_;
wire _11307_;
wire _11308_;
wire _11309_;
wire _11310_;
wire _11311_;
wire _11312_;
wire _11313_;
wire _11314_;
wire _11315_;
wire _11316_;
wire _11317_;
wire _11318_;
wire _11319_;
wire _11320_;
wire _11321_;
wire _11322_;
wire _11323_;
wire _11324_;
wire _11325_;
wire _11326_;
wire _11327_;
wire _11328_;
wire _11329_;
wire _11330_;
wire _11331_;
wire _11332_;
wire _11333_;
wire _11334_;
wire _11335_;
wire _11336_;
wire _11337_;
wire _11338_;
wire _11339_;
wire _11340_;
wire _11341_;
wire _11342_;
wire _11343_;
wire _11344_;
wire _11345_;
wire _11346_;
wire _11347_;
wire _11348_;
wire _11349_;
wire _11350_;
wire _11351_;
wire _11352_;
wire _11353_;
wire _11354_;
wire _11355_;
wire _11356_;
wire _11357_;
wire _11358_;
wire _11359_;
wire _11360_;
wire _11361_;
wire _11362_;
wire _11363_;
wire _11364_;
wire _11365_;
wire _11366_;
wire _11367_;
wire _11368_;
wire _11369_;
wire _11370_;
wire _11371_;
wire _11372_;
wire _11373_;
wire _11374_;
wire _11375_;
wire _11376_;
wire _11377_;
wire _11378_;
wire _11379_;
wire _11380_;
wire _11381_;
wire _11382_;
wire _11383_;
wire _11384_;
wire _11385_;
wire _11386_;
wire _11387_;
wire _11388_;
wire _11389_;
wire _11390_;
wire _11391_;
wire _11392_;
wire _11393_;
wire _11394_;
wire _11395_;
wire _11396_;
wire _11397_;
wire _11398_;
wire _11399_;
wire _11400_;
wire _11401_;
wire _11402_;
wire _11403_;
wire _11404_;
wire _11405_;
wire _11406_;
wire _11407_;
wire _11408_;
wire _11409_;
wire _11410_;
wire _11411_;
wire _11412_;
wire _11413_;
wire _11414_;
wire _11415_;
wire _11416_;
wire _11417_;
wire _11418_;
wire _11419_;
wire _11420_;
wire _11421_;
wire _11422_;
wire _11423_;
wire _11424_;
wire _11425_;
wire _11426_;
wire _11427_;
wire _11428_;
wire _11429_;
wire _11430_;
wire _11431_;
wire _11432_;
wire _11433_;
wire _11434_;
wire _11435_;
wire _11436_;
wire _11437_;
wire _11438_;
wire _11439_;
wire _11440_;
wire _11441_;
wire _11442_;
wire _11443_;
wire _11444_;
wire _11445_;
wire _11446_;
wire _11447_;
wire _11448_;
wire _11449_;
wire _11450_;
wire _11451_;
wire _11452_;
wire _11453_;
wire _11454_;
wire _11455_;
wire _11456_;
wire _11457_;
wire _11458_;
wire _11459_;
wire _11460_;
wire _11461_;
wire _11462_;
wire _11463_;
wire _11464_;
wire _11465_;
wire _11466_;
wire _11467_;
wire _11468_;
wire _11469_;
wire _11470_;
wire _11471_;
wire _11472_;
wire _11473_;
wire _11474_;
wire _11475_;
wire _11476_;
wire _11477_;
wire _11478_;
wire _11479_;
wire _11480_;
wire _11481_;
wire _11482_;
wire _11483_;
wire _11484_;
wire _11485_;
wire _11486_;
wire _11487_;
wire _11488_;
wire _11489_;
wire _11490_;
wire _11491_;
wire _11492_;
wire _11493_;
wire _11494_;
wire _11495_;
wire _11496_;
wire _11497_;
wire _11498_;
wire _11499_;
wire _11500_;
wire _11501_;
wire _11502_;
wire _11503_;
wire _11504_;
wire _11505_;
wire _11506_;
wire _11507_;
wire _11508_;
wire _11509_;
wire _11510_;
wire _11511_;
wire _11512_;
wire _11513_;
wire _11514_;
wire _11515_;
wire _11516_;
wire _11517_;
wire _11518_;
wire _11519_;
wire _11520_;
wire _11521_;
wire _11522_;
wire _11523_;
wire _11524_;
wire _11525_;
wire _11526_;
wire _11527_;
wire _11528_;
wire _11529_;
wire _11530_;
wire _11531_;
wire _11532_;
wire _11533_;
wire _11534_;
wire _11535_;
wire _11536_;
wire _11537_;
wire _11538_;
wire _11539_;
wire _11540_;
wire _11541_;
wire _11542_;
wire _11543_;
wire _11544_;
wire _11545_;
wire _11546_;
wire _11547_;
wire _11548_;
wire _11549_;
wire _11550_;
wire _11551_;
wire _11552_;
wire _11553_;
wire _11554_;
wire _11555_;
wire _11556_;
wire _11557_;
wire _11558_;
wire _11559_;
wire _11560_;
wire _11561_;
wire _11562_;
wire _11563_;
wire _11564_;
wire _11565_;
wire _11566_;
wire _11567_;
wire _11568_;
wire _11569_;
wire _11570_;
wire _11571_;
wire _11572_;
wire _11573_;
wire _11574_;
wire _11575_;
wire _11576_;
wire _11577_;
wire _11578_;
wire _11579_;
wire _11580_;
wire _11581_;
wire _11582_;
wire _11583_;
wire _11584_;
wire _11585_;
wire _11586_;
wire _11587_;
wire _11588_;
wire _11589_;
wire _11590_;
wire _11591_;
wire _11592_;
wire _11593_;
wire _11594_;
wire _11595_;
wire _11596_;
wire _11597_;
wire _11598_;
wire _11599_;
wire _11600_;
wire _11601_;
wire _11602_;
wire _11603_;
wire _11604_;
wire _11605_;
wire _11606_;
wire _11607_;
wire _11608_;
wire _11609_;
wire _11610_;
wire _11611_;
wire _11612_;
wire _11613_;
wire _11614_;
wire _11615_;
wire _11616_;
wire _11617_;
wire _11618_;
wire _11619_;
wire _11620_;
wire _11621_;
wire _11622_;
wire _11623_;
wire _11624_;
wire _11625_;
wire _11626_;
wire _11627_;
wire _11628_;
wire _11629_;
wire _11630_;
wire _11631_;
wire _11632_;
wire _11633_;
wire _11634_;
wire _11635_;
wire _11636_;
wire _11637_;
wire _11638_;
wire _11639_;
wire _11640_;
wire _11641_;
wire _11642_;
wire _11643_;
wire _11644_;
wire _11645_;
wire _11646_;
wire _11647_;
wire _11648_;
wire _11649_;
wire _11650_;
wire _11651_;
wire _11652_;
wire _11653_;
wire _11654_;
wire _11655_;
wire _11656_;
wire _11657_;
wire _11658_;
wire _11659_;
wire _11660_;
wire _11661_;
wire _11662_;
wire _11663_;
wire _11664_;
wire _11665_;
wire _11666_;
wire _11667_;
wire _11668_;
wire _11669_;
wire _11670_;
wire _11671_;
wire _11672_;
wire _11673_;
wire _11674_;
wire _11675_;
wire _11676_;
wire _11677_;
wire _11678_;
wire _11679_;
wire _11680_;
wire _11681_;
wire _11682_;
wire _11683_;
wire _11684_;
wire _11685_;
wire _11686_;
wire _11687_;
wire _11688_;
wire _11689_;
wire _11690_;
wire _11691_;
wire _11692_;
wire _11693_;
wire _11694_;
wire _11695_;
wire _11696_;
wire _11697_;
wire _11698_;
wire _11699_;
wire _11700_;
wire _11701_;
wire _11702_;
wire _11703_;
wire _11704_;
wire _11705_;
wire _11706_;
wire _11707_;
wire _11708_;
wire _11709_;
wire _11710_;
wire _11711_;
wire _11712_;
wire _11713_;
wire _11714_;
wire _11715_;
wire _11716_;
wire _11717_;
wire _11718_;
wire _11719_;
wire _11720_;
wire _11721_;
wire _11722_;
wire _11723_;
wire _11724_;
wire _11725_;
wire _11726_;
wire _11727_;
wire _11728_;
wire _11729_;
wire _11730_;
wire _11731_;
wire _11732_;
wire _11733_;
wire _11734_;
wire _11735_;
wire _11736_;
wire _11737_;
wire _11738_;
wire _11739_;
wire _11740_;
wire _11741_;
wire _11742_;
wire _11743_;
wire _11744_;
wire _11745_;
wire _11746_;
wire _11747_;
wire _11748_;
wire _11749_;
wire _11750_;
wire _11751_;
wire _11752_;
wire _11753_;
wire _11754_;
wire _11755_;
wire _11756_;
wire _11757_;
wire _11758_;
wire _11759_;
wire _11760_;
wire _11761_;
wire _11762_;
wire _11763_;
wire _11764_;
wire _11765_;
wire _11766_;
wire _11767_;
wire _11768_;
wire _11769_;
wire _11770_;
wire _11771_;
wire _11772_;
wire _11773_;
wire _11774_;
wire _11775_;
wire _11776_;
wire _11777_;
wire _11778_;
wire _11779_;
wire _11780_;
wire _11781_;
wire _11782_;
wire _11783_;
wire _11784_;
wire _11785_;
wire _11786_;
wire _11787_;
wire _11788_;
wire _11789_;
wire _11790_;
wire _11791_;
wire _11792_;
wire _11793_;
wire _11794_;
wire _11795_;
wire _11796_;
wire _11797_;
wire _11798_;
wire _11799_;
wire _11800_;
wire _11801_;
wire _11802_;
wire _11803_;
wire _11804_;
wire _11805_;
wire _11806_;
wire _11807_;
wire _11808_;
wire _11809_;
wire _11810_;
wire _11811_;
wire _11812_;
wire _11813_;
wire _11814_;
wire _11815_;
wire _11816_;
wire _11817_;
wire _11818_;
wire _11819_;
wire _11820_;
wire _11821_;
wire _11822_;
wire _11823_;
wire _11824_;
wire _11825_;
wire _11826_;
wire _11827_;
wire _11828_;
wire _11829_;
wire _11830_;
wire _11831_;
wire _11832_;
wire _11833_;
wire _11834_;
wire _11835_;
wire _11836_;
wire _11837_;
wire _11838_;
wire _11839_;
wire _11840_;
wire _11841_;
wire _11842_;
wire _11843_;
wire _11844_;
wire _11845_;
wire _11846_;
wire _11847_;
wire _11848_;
wire _11849_;
wire _11850_;
wire _11851_;
wire _11852_;
wire _11853_;
wire _11854_;
wire _11855_;
wire _11856_;
wire _11857_;
wire _11858_;
wire _11859_;
wire _11860_;
wire _11861_;
wire _11862_;
wire _11863_;
wire _11864_;
wire _11865_;
wire _11866_;
wire _11867_;
wire _11868_;
wire _11869_;
wire _11870_;
wire _11871_;
wire _11872_;
wire _11873_;
wire _11874_;
wire _11875_;
wire _11876_;
wire _11877_;
wire _11878_;
wire _11879_;
wire _11880_;
wire _11881_;
wire _11882_;
wire _11883_;
wire _11884_;
wire _11885_;
wire _11886_;
wire _11887_;
wire _11888_;
wire _11889_;
wire _11890_;
wire _11891_;
wire _11892_;
wire _11893_;
wire _11894_;
wire _11895_;
wire _11896_;
wire _11897_;
wire _11898_;
wire _11899_;
wire _11900_;
wire _11901_;
wire _11902_;
wire _11903_;
wire _11904_;
wire _11905_;
wire _11906_;
wire _11907_;
wire _11908_;
wire _11909_;
wire _11910_;
wire _11911_;
wire _11912_;
wire _11913_;
wire _11914_;
wire _11915_;
wire _11916_;
wire _11917_;
wire _11918_;
wire _11919_;
wire _11920_;
wire _11921_;
wire _11922_;
wire _11923_;
wire _11924_;
wire _11925_;
wire _11926_;
wire _11927_;
wire _11928_;
wire _11929_;
wire _11930_;
wire _11931_;
wire _11932_;
wire _11933_;
wire _11934_;
wire _11935_;
wire _11936_;
wire _11937_;
wire _11938_;
wire _11939_;
wire _11940_;
wire _11941_;
wire _11942_;
wire _11943_;
wire _11944_;
wire _11945_;
wire _11946_;
wire _11947_;
wire _11948_;
wire _11949_;
wire _11950_;
wire _11951_;
wire _11952_;
wire _11953_;
wire _11954_;
wire _11955_;
wire _11956_;
wire _11957_;
wire _11958_;
wire _11959_;
wire _11960_;
wire _11961_;
wire _11962_;
wire _11963_;
wire _11964_;
wire _11965_;
wire _11966_;
wire _11967_;
wire _11968_;
wire _11969_;
wire _11970_;
wire _11971_;
wire _11972_;
wire _11973_;
wire _11974_;
wire _11975_;
wire _11976_;
wire _11977_;
wire _11978_;
wire _11979_;
wire _11980_;
wire _11981_;
wire _11982_;
wire _11983_;
wire _11984_;
wire _11985_;
wire _11986_;
wire _11987_;
wire _11988_;
wire _11989_;
wire _11990_;
wire _11991_;
wire _11992_;
wire _11993_;
wire _11994_;
wire _11995_;
wire _11996_;
wire _11997_;
wire _11998_;
wire _11999_;
wire _12000_;
wire _12001_;
wire _12002_;
wire _12003_;
wire _12004_;
wire _12005_;
wire _12006_;
wire _12007_;
wire _12008_;
wire _12009_;
wire _12010_;
wire _12011_;
wire _12012_;
wire _12013_;
wire _12014_;
wire _12015_;
wire _12016_;
wire _12017_;
wire _12018_;
wire _12019_;
wire _12020_;
wire _12021_;
wire _12022_;
wire _12023_;
wire _12024_;
wire _12025_;
wire _12026_;
wire _12027_;
wire _12028_;
wire _12029_;
wire _12030_;
wire _12031_;
wire _12032_;
wire _12033_;
wire _12034_;
wire _12035_;
wire _12036_;
wire _12037_;
wire _12038_;
wire _12039_;
wire _12040_;
wire _12041_;
wire _12042_;
wire _12043_;
wire _12044_;
wire _12045_;
wire _12046_;
wire _12047_;
wire _12048_;
wire _12049_;
wire _12050_;
wire _12051_;
wire _12052_;
wire _12053_;
wire _12054_;
wire _12055_;
wire _12056_;
wire _12057_;
wire _12058_;
wire _12059_;
wire _12060_;
wire _12061_;
wire _12062_;
wire _12063_;
wire _12064_;
wire _12065_;
wire _12066_;
wire _12067_;
wire _12068_;
wire _12069_;
wire _12070_;
wire _12071_;
wire _12072_;
wire _12073_;
wire _12074_;
wire _12075_;
wire _12076_;
wire _12077_;
wire _12078_;
wire _12079_;
wire _12080_;
wire _12081_;
wire _12082_;
wire _12083_;
wire _12084_;
wire _12085_;
wire _12086_;
wire _12087_;
wire _12088_;
wire _12089_;
wire _12090_;
wire _12091_;
wire _12092_;
wire _12093_;
wire _12094_;
wire _12095_;
wire _12096_;
wire _12097_;
wire _12098_;
wire _12099_;
wire _12100_;
wire _12101_;
wire _12102_;
wire _12103_;
wire _12104_;
wire _12105_;
wire _12106_;
wire _12107_;
wire _12108_;
wire _12109_;
wire _12110_;
wire _12111_;
wire _12112_;
wire _12113_;
wire _12114_;
wire _12115_;
wire _12116_;
wire _12117_;
wire _12118_;
wire _12119_;
wire _12120_;
wire _12121_;
wire _12122_;
wire _12123_;
wire _12124_;
wire _12125_;
wire _12126_;
wire _12127_;
wire _12128_;
wire _12129_;
wire _12130_;
wire _12131_;
wire _12132_;
wire _12133_;
wire _12134_;
wire _12135_;
wire _12136_;
wire _12137_;
wire _12138_;
wire _12139_;
wire _12140_;
wire _12141_;
wire _12142_;
wire _12143_;
wire _12144_;
wire _12145_;
wire _12146_;
wire _12147_;
wire _12148_;
wire _12149_;
wire _12150_;
wire _12151_;
wire _12152_;
wire _12153_;
wire _12154_;
wire _12155_;
wire _12156_;
wire _12157_;
wire _12158_;
wire _12159_;
wire _12160_;
wire _12161_;
wire _12162_;
wire _12163_;
wire _12164_;
wire _12165_;
wire _12166_;
wire _12167_;
wire _12168_;
wire _12169_;
wire _12170_;
wire _12171_;
wire _12172_;
wire _12173_;
wire _12174_;
wire _12175_;
wire _12176_;
wire _12177_;
wire _12178_;
wire _12179_;
wire _12180_;
wire _12181_;
wire _12182_;
wire _12183_;
wire _12184_;
wire _12185_;
wire _12186_;
wire _12187_;
wire _12188_;
wire _12189_;
wire _12190_;
wire _12191_;
wire _12192_;
wire _12193_;
wire _12194_;
wire _12195_;
wire _12196_;
wire _12197_;
wire _12198_;
wire _12199_;
wire _12200_;
wire _12201_;
wire _12202_;
wire _12203_;
wire _12204_;
wire _12205_;
wire _12206_;
wire _12207_;
wire _12208_;
wire _12209_;
wire _12210_;
wire _12211_;
wire _12212_;
wire _12213_;
wire _12214_;
wire _12215_;
wire _12216_;
wire _12217_;
wire _12218_;
wire _12219_;
wire _12220_;
wire _12221_;
wire _12222_;
wire _12223_;
wire _12224_;
wire _12225_;
wire _12226_;
wire _12227_;
wire _12228_;
wire _12229_;
wire _12230_;
wire _12231_;
wire _12232_;
wire _12233_;
wire _12234_;
wire _12235_;
wire _12236_;
wire _12237_;
wire _12238_;
wire _12239_;
wire _12240_;
wire _12241_;
wire _12242_;
wire _12243_;
wire _12244_;
wire _12245_;
wire _12246_;
wire _12247_;
wire _12248_;
wire _12249_;
wire _12250_;
wire _12251_;
wire _12252_;
wire _12253_;
wire _12254_;
wire _12255_;
wire _12256_;
wire _12257_;
wire _12258_;
wire _12259_;
wire _12260_;
wire _12261_;
wire _12262_;
wire _12263_;
wire _12264_;
wire _12265_;
wire _12266_;
wire _12267_;
wire _12268_;
wire _12269_;
wire _12270_;
wire _12271_;
wire _12272_;
wire _12273_;
wire _12274_;
wire _12275_;
wire _12276_;
wire _12277_;
wire _12278_;
wire _12279_;
wire _12280_;
wire _12281_;
wire _12282_;
wire _12283_;
wire _12284_;
wire _12285_;
wire _12286_;
wire _12287_;
wire _12288_;
wire _12289_;
wire _12290_;
wire _12291_;
wire _12292_;
wire _12293_;
wire _12294_;
wire _12295_;
wire _12296_;
wire _12297_;
wire _12298_;
wire _12299_;
wire _12300_;
wire _12301_;
wire _12302_;
wire _12303_;
wire _12304_;
wire _12305_;
wire _12306_;
wire _12307_;
wire _12308_;
wire _12309_;
wire _12310_;
wire _12311_;
wire _12312_;
wire _12313_;
wire _12314_;
wire _12315_;
wire _12316_;
wire _12317_;
wire _12318_;
wire _12319_;
wire _12320_;
wire _12321_;
wire _12322_;
wire _12323_;
wire _12324_;
wire _12325_;
wire _12326_;
wire _12327_;
wire _12328_;
wire _12329_;
wire _12330_;
wire _12331_;
wire _12332_;
wire _12333_;
wire _12334_;
wire _12335_;
wire _12336_;
wire _12337_;
wire _12338_;
wire _12339_;
wire _12340_;
wire _12341_;
wire _12342_;
wire _12343_;
wire _12344_;
wire _12345_;
wire _12346_;
wire _12347_;
wire _12348_;
wire _12349_;
wire _12350_;
wire _12351_;
wire _12352_;
wire _12353_;
wire _12354_;
wire _12355_;
wire _12356_;
wire _12357_;
wire _12358_;
wire _12359_;
wire _12360_;
wire _12361_;
wire _12362_;
wire _12363_;
wire _12364_;
wire _12365_;
wire _12366_;
wire _12367_;
wire _12368_;
wire _12369_;
wire _12370_;
wire _12371_;
wire _12372_;
wire _12373_;
wire _12374_;
wire _12375_;
wire _12376_;
wire _12377_;
wire _12378_;
wire _12379_;
wire _12380_;
wire _12381_;
wire _12382_;
wire _12383_;
wire _12384_;
wire _12385_;
wire _12386_;
wire _12387_;
wire _12388_;
wire _12389_;
wire _12390_;
wire _12391_;
wire _12392_;
wire _12393_;
wire _12394_;
wire _12395_;
wire _12396_;
wire _12397_;
wire _12398_;
wire _12399_;
wire _12400_;
wire _12401_;
wire _12402_;
wire _12403_;
wire _12404_;
wire _12405_;
wire _12406_;
wire _12407_;
wire _12408_;
wire _12409_;
wire _12410_;
wire _12411_;
wire _12412_;
wire _12413_;
wire _12414_;
wire _12415_;
wire _12416_;
wire _12417_;
wire _12418_;
wire _12419_;
wire _12420_;
wire _12421_;
wire _12422_;
wire _12423_;
wire _12424_;
wire _12425_;
wire _12426_;
wire _12427_;
wire _12428_;
wire _12429_;
wire _12430_;
wire _12431_;
wire _12432_;
wire _12433_;
wire _12434_;
wire _12435_;
wire _12436_;
wire _12437_;
wire _12438_;
wire _12439_;
wire _12440_;
wire _12441_;
wire _12442_;
wire _12443_;
wire _12444_;
wire _12445_;
wire _12446_;
wire _12447_;
wire _12448_;
wire _12449_;
wire _12450_;
wire _12451_;
wire _12452_;
wire _12453_;
wire _12454_;
wire _12455_;
wire _12456_;
wire _12457_;
wire _12458_;
wire _12459_;
wire _12460_;
wire _12461_;
wire _12462_;
wire _12463_;
wire _12464_;
wire _12465_;
wire _12466_;
wire _12467_;
wire _12468_;
wire _12469_;
wire _12470_;
wire _12471_;
wire _12472_;
wire _12473_;
wire _12474_;
wire _12475_;
wire _12476_;
wire _12477_;
wire _12478_;
wire _12479_;
wire _12480_;
wire _12481_;
wire _12482_;
wire _12483_;
wire _12484_;
wire _12485_;
wire _12486_;
wire _12487_;
wire _12488_;
wire _12489_;
wire _12490_;
wire _12491_;
wire _12492_;
wire _12493_;
wire _12494_;
wire _12495_;
wire _12496_;
wire _12497_;
wire _12498_;
wire _12499_;
wire _12500_;
wire _12501_;
wire _12502_;
wire _12503_;
wire _12504_;
wire _12505_;
wire _12506_;
wire _12507_;
wire _12508_;
wire _12509_;
wire _12510_;
wire _12511_;
wire _12512_;
wire _12513_;
wire _12514_;
wire _12515_;
wire _12516_;
wire _12517_;
wire _12518_;
wire _12519_;
wire _12520_;
wire _12521_;
wire _12522_;
wire _12523_;
wire _12524_;
wire _12525_;
wire _12526_;
wire _12527_;
wire _12528_;
wire _12529_;
wire _12530_;
wire _12531_;
wire _12532_;
wire _12533_;
wire _12534_;
wire _12535_;
wire _12536_;
wire _12537_;
wire _12538_;
wire _12539_;
wire _12540_;
wire _12541_;
wire _12542_;
wire _12543_;
wire _12544_;
wire _12545_;
wire _12546_;
wire _12547_;
wire _12548_;
wire _12549_;
wire _12550_;
wire _12551_;
wire _12552_;
wire _12553_;
wire _12554_;
wire _12555_;
wire _12556_;
wire _12557_;
wire _12558_;
wire _12559_;
wire _12560_;
wire _12561_;
wire _12562_;
wire _12563_;
wire _12564_;
wire _12565_;
wire _12566_;
wire _12567_;
wire _12568_;
wire _12569_;
wire _12570_;
wire _12571_;
wire _12572_;
wire _12573_;
wire _12574_;
wire _12575_;
wire _12576_;
wire _12577_;
wire _12578_;
wire _12579_;
wire _12580_;
wire _12581_;
wire _12582_;
wire _12583_;
wire _12584_;
wire _12585_;
wire _12586_;
wire _12587_;
wire _12588_;
wire _12589_;
wire _12590_;
wire _12591_;
wire _12592_;
wire _12593_;
wire _12594_;
wire _12595_;
wire _12596_;
wire _12597_;
wire _12598_;
wire _12599_;
wire _12600_;
wire _12601_;
wire _12602_;
wire _12603_;
wire _12604_;
wire _12605_;
wire _12606_;
wire _12607_;
wire _12608_;
wire _12609_;
wire _12610_;
wire _12611_;
wire _12612_;
wire _12613_;
wire _12614_;
wire _12615_;
wire _12616_;
wire _12617_;
wire _12618_;
wire _12619_;
wire _12620_;
wire _12621_;
wire _12622_;
wire _12623_;
wire _12624_;
wire _12625_;
wire _12626_;
wire _12627_;
wire _12628_;
wire _12629_;
wire _12630_;
wire _12631_;
wire _12632_;
wire _12633_;
wire _12634_;
wire _12635_;
wire _12636_;
wire _12637_;
wire _12638_;
wire _12639_;
wire _12640_;
wire _12641_;
wire _12642_;
wire _12643_;
wire _12644_;
wire _12645_;
wire _12646_;
wire _12647_;
wire _12648_;
wire _12649_;
wire _12650_;
wire _12651_;
wire _12652_;
wire _12653_;
wire _12654_;
wire _12655_;
wire _12656_;
wire _12657_;
wire _12658_;
wire _12659_;
wire _12660_;
wire _12661_;
wire _12662_;
wire _12663_;
wire _12664_;
wire _12665_;
wire _12666_;
wire _12667_;
wire _12668_;
wire _12669_;
wire _12670_;
wire _12671_;
wire _12672_;
wire _12673_;
wire _12674_;
wire _12675_;
wire _12676_;
wire _12677_;
wire _12678_;
wire _12679_;
wire _12680_;
wire _12681_;
wire _12682_;
wire _12683_;
wire _12684_;
wire _12685_;
wire _12686_;
wire _12687_;
wire _12688_;
wire _12689_;
wire _12690_;
wire _12691_;
wire _12692_;
wire _12693_;
wire _12694_;
wire _12695_;
wire _12696_;
wire _12697_;
wire _12698_;
wire _12699_;
wire _12700_;
wire _12701_;
wire _12702_;
wire _12703_;
wire _12704_;
wire _12705_;
wire _12706_;
wire _12707_;
wire _12708_;
wire _12709_;
wire _12710_;
wire _12711_;
wire _12712_;
wire _12713_;
wire _12714_;
wire _12715_;
wire _12716_;
wire _12717_;
wire _12718_;
wire _12719_;
wire _12720_;
wire _12721_;
wire _12722_;
wire _12723_;
wire _12724_;
wire _12725_;
wire _12726_;
wire _12727_;
wire _12728_;
wire _12729_;
wire _12730_;
wire _12731_;
wire _12732_;
wire _12733_;
wire _12734_;
wire _12735_;
wire _12736_;
wire _12737_;
wire _12738_;
wire _12739_;
wire _12740_;
wire _12741_;
wire _12742_;
wire _12743_;
wire _12744_;
wire _12745_;
wire _12746_;
wire _12747_;
wire _12748_;
wire _12749_;
wire _12750_;
wire _12751_;
wire _12752_;
wire _12753_;
wire _12754_;
wire _12755_;
wire _12756_;
wire _12757_;
wire _12758_;
wire _12759_;
wire _12760_;
wire _12761_;
wire _12762_;
wire _12763_;
wire _12764_;
wire _12765_;
wire _12766_;
wire _12767_;
wire _12768_;
wire _12769_;
wire _12770_;
wire _12771_;
wire _12772_;
wire _12773_;
wire _12774_;
wire _12775_;
wire _12776_;
wire _12777_;
wire _12778_;
wire _12779_;
wire _12780_;
wire _12781_;
wire _12782_;
wire _12783_;
wire _12784_;
wire _12785_;
wire _12786_;
wire _12787_;
wire _12788_;
wire _12789_;
wire _12790_;
wire _12791_;
wire _12792_;
wire _12793_;
wire _12794_;
wire _12795_;
wire _12796_;
wire _12797_;
wire _12798_;
wire _12799_;
wire _12800_;
wire _12801_;
wire _12802_;
wire _12803_;
wire _12804_;
wire _12805_;
wire _12806_;
wire _12807_;
wire _12808_;
wire _12809_;
wire _12810_;
wire _12811_;
wire _12812_;
wire _12813_;
wire _12814_;
wire _12815_;
wire _12816_;
wire _12817_;
wire _12818_;
wire _12819_;
wire _12820_;
wire _12821_;
wire _12822_;
wire _12823_;
wire _12824_;
wire _12825_;
wire _12826_;
wire _12827_;
wire _12828_;
wire _12829_;
wire _12830_;
wire _12831_;
wire _12832_;
wire _12833_;
wire _12834_;
wire _12835_;
wire _12836_;
wire _12837_;
wire _12838_;
wire _12839_;
wire _12840_;
wire _12841_;
wire _12842_;
wire _12843_;
wire _12844_;
wire _12845_;
wire _12846_;
wire _12847_;
wire _12848_;
wire _12849_;
wire _12850_;
wire _12851_;
wire _12852_;
wire _12853_;
wire _12854_;
wire _12855_;
wire _12856_;
wire _12857_;
wire _12858_;
wire _12859_;
wire _12860_;
wire _12861_;
wire _12862_;
wire _12863_;
wire _12864_;
wire _12865_;
wire _12866_;
wire _12867_;
wire _12868_;
wire _12869_;
wire _12870_;
wire _12871_;
wire _12872_;
wire _12873_;
wire _12874_;
wire _12875_;
wire _12876_;
wire _12877_;
wire _12878_;
wire _12879_;
wire _12880_;
wire _12881_;
wire _12882_;
wire _12883_;
wire _12884_;
wire _12885_;
wire _12886_;
wire _12887_;
wire _12888_;
wire _12889_;
wire _12890_;
wire _12891_;
wire _12892_;
wire _12893_;
wire _12894_;
wire _12895_;
wire _12896_;
wire _12897_;
wire _12898_;
wire _12899_;
wire _12900_;
wire _12901_;
wire _12902_;
wire _12903_;
wire _12904_;
wire _12905_;
wire _12906_;
wire _12907_;
wire _12908_;
wire _12909_;
wire _12910_;
wire _12911_;
wire _12912_;
wire _12913_;
wire _12914_;
wire _12915_;
wire _12916_;
wire _12917_;
wire _12918_;
wire _12919_;
wire _12920_;
wire _12921_;
wire _12922_;
wire _12923_;
wire _12924_;
wire _12925_;
wire _12926_;
wire _12927_;
wire _12928_;
wire _12929_;
wire _12930_;
wire _12931_;
wire _12932_;
wire _12933_;
wire _12934_;
wire _12935_;
wire _12936_;
wire _12937_;
wire _12938_;
wire _12939_;
wire _12940_;
wire _12941_;
wire _12942_;
wire _12943_;
wire _12944_;
wire _12945_;
wire _12946_;
wire _12947_;
wire _12948_;
wire _12949_;
wire _12950_;
wire _12951_;
wire _12952_;
wire _12953_;
wire _12954_;
wire _12955_;
wire _12956_;
wire _12957_;
wire _12958_;
wire _12959_;
wire _12960_;
wire _12961_;
wire _12962_;
wire _12963_;
wire _12964_;
wire _12965_;
wire _12966_;
wire _12967_;
wire _12968_;
wire _12969_;
wire _12970_;
wire _12971_;
wire _12972_;
wire _12973_;
wire _12974_;
wire _12975_;
wire _12976_;
wire _12977_;
wire _12978_;
wire _12979_;
wire _12980_;
wire _12981_;
wire _12982_;
wire _12983_;
wire _12984_;
wire _12985_;
wire _12986_;
wire _12987_;
wire _12988_;
wire _12989_;
wire _12990_;
wire _12991_;
wire _12992_;
wire _12993_;
wire _12994_;
wire _12995_;
wire _12996_;
wire _12997_;
wire _12998_;
wire _12999_;
wire _13000_;
wire _13001_;
wire _13002_;
wire _13003_;
wire _13004_;
wire _13005_;
wire _13006_;
wire _13007_;
wire _13008_;
wire _13009_;
wire _13010_;
wire _13011_;
wire _13012_;
wire _13013_;
wire _13014_;
wire _13015_;
wire _13016_;
wire _13017_;
wire _13018_;
wire _13019_;
wire _13020_;
wire _13021_;
wire _13022_;
wire _13023_;
wire _13024_;
wire _13025_;
wire _13026_;
wire _13027_;
wire _13028_;
wire _13029_;
wire _13030_;
wire _13031_;
wire _13032_;
wire _13033_;
wire _13034_;
wire _13035_;
wire _13036_;
wire _13037_;
wire _13038_;
wire _13039_;
wire _13040_;
wire _13041_;
wire _13042_;
wire _13043_;
wire _13044_;
wire _13045_;
wire _13046_;
wire _13047_;
wire _13048_;
wire _13049_;
wire _13050_;
wire _13051_;
wire _13052_;
wire _13053_;
wire _13054_;
wire _13055_;
wire _13056_;
wire _13057_;
wire _13058_;
wire _13059_;
wire _13060_;
wire _13061_;
wire _13062_;
wire _13063_;
wire _13064_;
wire _13065_;
wire _13066_;
wire _13067_;
wire _13068_;
wire _13069_;
wire _13070_;
wire _13071_;
wire _13072_;
wire _13073_;
wire _13074_;
wire _13075_;
wire _13076_;
wire _13077_;
wire _13078_;
wire _13079_;
wire _13080_;
wire _13081_;
wire _13082_;
wire _13083_;
wire _13084_;
wire _13085_;
wire _13086_;
wire _13087_;
wire _13088_;
wire _13089_;
wire _13090_;
wire _13091_;
wire _13092_;
wire _13093_;
wire _13094_;
wire _13095_;
wire _13096_;
wire _13097_;
wire _13098_;
wire _13099_;
wire _13100_;
wire _13101_;
wire _13102_;
wire _13103_;
wire _13104_;
wire _13105_;
wire _13106_;
wire _13107_;
wire _13108_;
wire _13109_;
wire _13110_;
wire _13111_;
wire _13112_;
wire _13113_;
wire _13114_;
wire _13115_;
wire _13116_;
wire _13117_;
wire _13118_;
wire _13119_;
wire _13120_;
wire _13121_;
wire _13122_;
wire _13123_;
wire _13124_;
wire _13125_;
wire _13126_;
wire _13127_;
wire _13128_;
wire _13129_;
wire _13130_;
wire _13131_;
wire _13132_;
wire _13133_;
wire _13134_;
wire _13135_;
wire _13136_;
wire _13137_;
wire _13138_;
wire _13139_;
wire _13140_;
wire _13141_;
wire _13142_;
wire _13143_;
wire _13144_;
wire _13145_;
wire _13146_;
wire _13147_;
wire _13148_;
wire _13149_;
wire _13150_;
wire _13151_;
wire _13152_;
wire _13153_;
wire _13154_;
wire _13155_;
wire _13156_;
wire _13157_;
wire _13158_;
wire _13159_;
wire _13160_;
wire _13161_;
wire _13162_;
wire _13163_;
wire _13164_;
wire _13165_;
wire _13166_;
wire _13167_;
wire _13168_;
wire _13169_;
wire _13170_;
wire _13171_;
wire _13172_;
wire _13173_;
wire _13174_;
wire _13175_;
wire _13176_;
wire _13177_;
wire _13178_;
wire _13179_;
wire _13180_;
wire _13181_;
wire _13182_;
wire _13183_;
wire _13184_;
wire _13185_;
wire _13186_;
wire _13187_;
wire _13188_;
wire _13189_;
wire _13190_;
wire _13191_;
wire _13192_;
wire _13193_;
wire _13194_;
wire _13195_;
wire _13196_;
wire _13197_;
wire _13198_;
wire _13199_;
wire _13200_;
wire _13201_;
wire _13202_;
wire _13203_;
wire _13204_;
wire _13205_;
wire _13206_;
wire _13207_;
wire _13208_;
wire _13209_;
wire _13210_;
wire _13211_;
wire _13212_;
wire _13213_;
wire _13214_;
wire _13215_;
wire _13216_;
wire _13217_;
wire _13218_;
wire _13219_;
wire _13220_;
wire _13221_;
wire _13222_;
wire _13223_;
wire _13224_;
wire _13225_;
wire _13226_;
wire _13227_;
wire _13228_;
wire _13229_;
wire _13230_;
wire _13231_;
wire _13232_;
wire _13233_;
wire _13234_;
wire _13235_;
wire _13236_;
wire _13237_;
wire _13238_;
wire _13239_;
wire _13240_;
wire _13241_;
wire _13242_;
wire _13243_;
wire _13244_;
wire _13245_;
wire _13246_;
wire _13247_;
wire _13248_;
wire _13249_;
wire _13250_;
wire _13251_;
wire _13252_;
wire _13253_;
wire _13254_;
wire _13255_;
wire _13256_;
wire _13257_;
wire _13258_;
wire _13259_;
wire _13260_;
wire _13261_;
wire _13262_;
wire _13263_;
wire _13264_;
wire _13265_;
wire _13266_;
wire _13267_;
wire _13268_;
wire _13269_;
wire _13270_;
wire _13271_;
wire _13272_;
wire _13273_;
wire _13274_;
wire _13275_;
wire _13276_;
wire _13277_;
wire _13278_;
wire _13279_;
wire _13280_;
wire _13281_;
wire _13282_;
wire _13283_;
wire _13284_;
wire _13285_;
wire _13286_;
wire _13287_;
wire _13288_;
wire _13289_;
wire _13290_;
wire _13291_;
wire _13292_;
wire _13293_;
wire _13294_;
wire _13295_;
wire _13296_;
wire _13297_;
wire _13298_;
wire _13299_;
wire _13300_;
wire _13301_;
wire _13302_;
wire _13303_;
wire _13304_;
wire _13305_;
wire _13306_;
wire _13307_;
wire _13308_;
wire _13309_;
wire _13310_;
wire _13311_;
wire _13312_;
wire _13313_;
wire _13314_;
wire _13315_;
wire _13316_;
wire _13317_;
wire _13318_;
wire _13319_;
wire _13320_;
wire _13321_;
wire _13322_;
wire _13323_;
wire _13324_;
wire _13325_;
wire _13326_;
wire _13327_;
wire _13328_;
wire _13329_;
wire _13330_;
wire _13331_;
wire _13332_;
wire _13333_;
wire _13334_;
wire _13335_;
wire _13336_;
wire _13337_;
wire _13338_;
wire _13339_;
wire _13340_;
wire _13341_;
wire _13342_;
wire _13343_;
wire _13344_;
wire _13345_;
wire _13346_;
wire _13347_;
wire _13348_;
wire _13349_;
wire _13350_;
wire _13351_;
wire _13352_;
wire _13353_;
wire _13354_;
wire _13355_;
wire _13356_;
wire _13357_;
wire _13358_;
wire _13359_;
wire _13360_;
wire _13361_;
wire _13362_;
wire _13363_;
wire _13364_;
wire _13365_;
wire _13366_;
wire _13367_;
wire _13368_;
wire _13369_;
wire _13370_;
wire _13371_;
wire _13372_;
wire _13373_;
wire _13374_;
wire _13375_;
wire _13376_;
wire _13377_;
wire _13378_;
wire _13379_;
wire _13380_;
wire _13381_;
wire _13382_;
wire _13383_;
wire _13384_;
wire _13385_;
wire _13386_;
wire _13387_;
wire _13388_;
wire _13389_;
wire _13390_;
wire _13391_;
wire _13392_;
wire _13393_;
wire _13394_;
wire _13395_;
wire _13396_;
wire _13397_;
wire _13398_;
wire _13399_;
wire _13400_;
wire _13401_;
wire _13402_;
wire _13403_;
wire _13404_;
wire _13405_;
wire _13406_;
wire _13407_;
wire _13408_;
wire _13409_;
wire _13410_;
wire _13411_;
wire _13412_;
wire _13413_;
wire _13414_;
wire _13415_;
wire _13416_;
wire _13417_;
wire _13418_;
wire _13419_;
wire _13420_;
wire _13421_;
wire _13422_;
wire _13423_;
wire _13424_;
wire _13425_;
wire _13426_;
wire _13427_;
wire _13428_;
wire _13429_;
wire _13430_;
wire _13431_;
wire _13432_;
wire _13433_;
wire _13434_;
wire _13435_;
wire _13436_;
wire _13437_;
wire _13438_;
wire _13439_;
wire _13440_;
wire _13441_;
wire _13442_;
wire _13443_;
wire _13444_;
wire _13445_;
wire _13446_;
wire _13447_;
wire _13448_;
wire _13449_;
wire _13450_;
wire _13451_;
wire _13452_;
wire _13453_;
wire _13454_;
wire _13455_;
wire _13456_;
wire _13457_;
wire _13458_;
wire _13459_;
wire _13460_;
wire _13461_;
wire _13462_;
wire _13463_;
wire _13464_;
wire _13465_;
wire _13466_;
wire _13467_;
wire _13468_;
wire _13469_;
wire _13470_;
wire _13471_;
wire _13472_;
wire _13473_;
wire _13474_;
wire _13475_;
wire _13476_;
wire _13477_;
wire _13478_;
wire _13479_;
wire _13480_;
wire _13481_;
wire _13482_;
wire _13483_;
wire _13484_;
wire _13485_;
wire _13486_;
wire _13487_;
wire _13488_;
wire _13489_;
wire _13490_;
wire _13491_;
wire _13492_;
wire _13493_;
wire _13494_;
wire _13495_;
wire _13496_;
wire _13497_;
wire _13498_;
wire _13499_;
wire _13500_;
wire _13501_;
wire _13502_;
wire _13503_;
wire _13504_;
wire _13505_;
wire _13506_;
wire _13507_;
wire _13508_;
wire _13509_;
wire _13510_;
wire _13511_;
wire _13512_;
wire _13513_;
wire _13514_;
wire _13515_;
wire _13516_;
wire _13517_;
wire _13518_;
wire _13519_;
wire _13520_;
wire _13521_;
wire _13522_;
wire _13523_;
wire _13524_;
wire _13525_;
wire _13526_;
wire _13527_;
wire _13528_;
wire _13529_;
wire _13530_;
wire _13531_;
wire _13532_;
wire _13533_;
wire _13534_;
wire _13535_;
wire _13536_;
wire _13537_;
wire _13538_;
wire _13539_;
wire _13540_;
wire _13541_;
wire _13542_;
wire _13543_;
wire _13544_;
wire _13545_;
wire _13546_;
wire _13547_;
wire _13548_;
wire _13549_;
wire _13550_;
wire _13551_;
wire _13552_;
wire _13553_;
wire _13554_;
wire _13555_;
wire _13556_;
wire _13557_;
wire _13558_;
wire _13559_;
wire _13560_;
wire _13561_;
wire _13562_;
wire _13563_;
wire _13564_;
wire _13565_;
wire _13566_;
wire _13567_;
wire _13568_;
wire _13569_;
wire _13570_;
wire _13571_;
wire _13572_;
wire _13573_;
wire _13574_;
wire _13575_;
wire _13576_;
wire _13577_;
wire _13578_;
wire _13579_;
wire _13580_;
wire _13581_;
wire _13582_;
wire _13583_;
wire _13584_;
wire _13585_;
wire _13586_;
wire _13587_;
wire _13588_;
wire _13589_;
wire _13590_;
wire _13591_;
wire _13592_;
wire _13593_;
wire _13594_;
wire _13595_;
wire _13596_;
wire _13597_;
wire _13598_;
wire _13599_;
wire _13600_;
wire _13601_;
wire _13602_;
wire _13603_;
wire _13604_;
wire _13605_;
wire _13606_;
wire _13607_;
wire _13608_;
wire _13609_;
wire _13610_;
wire _13611_;
wire _13612_;
wire _13613_;
wire _13614_;
wire _13615_;
wire _13616_;
wire _13617_;
wire _13618_;
wire _13619_;
wire _13620_;
wire _13621_;
wire _13622_;
wire _13623_;
wire _13624_;
wire _13625_;
wire _13626_;
wire _13627_;
wire _13628_;
wire _13629_;
wire _13630_;
wire _13631_;
wire _13632_;
wire _13633_;
wire _13634_;
wire _13635_;
wire _13636_;
wire _13637_;
wire _13638_;
wire _13639_;
wire _13640_;
wire _13641_;
wire _13642_;
wire _13643_;
wire _13644_;
wire _13645_;
wire _13646_;
wire _13647_;
wire _13648_;
wire _13649_;
wire _13650_;
wire _13651_;
wire _13652_;
wire _13653_;
wire _13654_;
wire _13655_;
wire _13656_;
wire _13657_;
wire _13658_;
wire _13659_;
wire _13660_;
wire _13661_;
wire _13662_;
wire _13663_;
wire _13664_;
wire _13665_;
wire _13666_;
wire _13667_;
wire _13668_;
wire _13669_;
wire _13670_;
wire _13671_;
wire _13672_;
wire _13673_;
wire _13674_;
wire _13675_;
wire _13676_;
wire _13677_;
wire _13678_;
wire _13679_;
wire _13680_;
wire _13681_;
wire _13682_;
wire _13683_;
wire _13684_;
wire _13685_;
wire _13686_;
wire _13687_;
wire _13688_;
wire _13689_;
wire _13690_;
wire _13691_;
wire _13692_;
wire _13693_;
wire _13694_;
wire _13695_;
wire _13696_;
wire _13697_;
wire _13698_;
wire _13699_;
wire _13700_;
wire _13701_;
wire _13702_;
wire _13703_;
wire _13704_;
wire _13705_;
wire _13706_;
wire _13707_;
wire _13708_;
wire _13709_;
wire _13710_;
wire _13711_;
wire _13712_;
wire _13713_;
wire _13714_;
wire _13715_;
wire _13716_;
wire _13717_;
wire _13718_;
wire _13719_;
wire _13720_;
wire _13721_;
wire _13722_;
wire _13723_;
wire _13724_;
wire _13725_;
wire _13726_;
wire _13727_;
wire _13728_;
wire _13729_;
wire _13730_;
wire _13731_;
wire _13732_;
wire _13733_;
wire _13734_;
wire _13735_;
wire _13736_;
wire _13737_;
wire _13738_;
wire _13739_;
wire _13740_;
wire _13741_;
wire _13742_;
wire _13743_;
wire _13744_;
wire _13745_;
wire _13746_;
wire _13747_;
wire _13748_;
wire _13749_;
wire _13750_;
wire _13751_;
wire _13752_;
wire _13753_;
wire _13754_;
wire _13755_;
wire _13756_;
wire _13757_;
wire _13758_;
wire _13759_;
wire _13760_;
wire _13761_;
wire _13762_;
wire _13763_;
wire _13764_;
wire _13765_;
wire _13766_;
wire _13767_;
wire _13768_;
wire _13769_;
wire _13770_;
wire _13771_;
wire _13772_;
wire _13773_;
wire _13774_;
wire _13775_;
wire _13776_;
wire _13777_;
wire _13778_;
wire _13779_;
wire _13780_;
wire _13781_;
wire _13782_;
wire _13783_;
wire _13784_;
wire _13785_;
wire _13786_;
wire _13787_;
wire _13788_;
wire _13789_;
wire _13790_;
wire _13791_;
wire _13792_;
wire _13793_;
wire _13794_;
wire _13795_;
wire _13796_;
wire _13797_;
wire _13798_;
wire _13799_;
wire _13800_;
wire _13801_;
wire _13802_;
wire _13803_;
wire _13804_;
wire _13805_;
wire _13806_;
wire _13807_;
wire _13808_;
wire _13809_;
wire _13810_;
wire _13811_;
wire _13812_;
wire _13813_;
wire _13814_;
wire _13815_;
wire _13816_;
wire _13817_;
wire _13818_;
wire _13819_;
wire _13820_;
wire _13821_;
wire _13822_;
wire _13823_;
wire _13824_;
wire _13825_;
wire _13826_;
wire _13827_;
wire _13828_;
wire _13829_;
wire _13830_;
wire _13831_;
wire _13832_;
wire _13833_;
wire _13834_;
wire _13835_;
wire _13836_;
wire _13837_;
wire _13838_;
wire _13839_;
wire _13840_;
wire _13841_;
wire _13842_;
wire _13843_;
wire _13844_;
wire _13845_;
wire _13846_;
wire _13847_;
wire _13848_;
wire _13849_;
wire _13850_;
wire _13851_;
wire _13852_;
wire _13853_;
wire _13854_;
wire _13855_;
wire _13856_;
wire _13857_;
wire _13858_;
wire _13859_;
wire _13860_;
wire _13861_;
wire _13862_;
wire _13863_;
wire _13864_;
wire _13865_;
wire _13866_;
wire _13867_;
wire _13868_;
wire _13869_;
wire _13870_;
wire _13871_;
wire _13872_;
wire _13873_;
wire _13874_;
wire _13875_;
wire _13876_;
wire _13877_;
wire _13878_;
wire _13879_;
wire _13880_;
wire _13881_;
wire _13882_;
wire _13883_;
wire _13884_;
wire _13885_;
wire _13886_;
wire _13887_;
wire _13888_;
wire _13889_;
wire _13890_;
wire _13891_;
wire _13892_;
wire _13893_;
wire _13894_;
wire _13895_;
wire _13896_;
wire _13897_;
wire _13898_;
wire _13899_;
wire _13900_;
wire _13901_;
wire _13902_;
wire _13903_;
wire _13904_;
wire _13905_;
wire _13906_;
wire _13907_;
wire _13908_;
wire _13909_;
wire _13910_;
wire _13911_;
wire _13912_;
wire _13913_;
wire _13914_;
wire _13915_;
wire _13916_;
wire _13917_;
wire _13918_;
wire _13919_;
wire _13920_;
wire _13921_;
wire _13922_;
wire _13923_;
wire _13924_;
wire _13925_;
wire _13926_;
wire _13927_;
wire _13928_;
wire _13929_;
wire _13930_;
wire _13931_;
wire _13932_;
wire _13933_;
wire _13934_;
wire _13935_;
wire _13936_;
wire _13937_;
wire _13938_;
wire _13939_;
wire _13940_;
wire _13941_;
wire _13942_;
wire _13943_;
wire _13944_;
wire _13945_;
wire _13946_;
wire _13947_;
wire _13948_;
wire _13949_;
wire _13950_;
wire _13951_;
wire _13952_;
wire _13953_;
wire _13954_;
wire _13955_;
wire _13956_;
wire _13957_;
wire _13958_;
wire _13959_;
wire _13960_;
wire _13961_;
wire _13962_;
wire _13963_;
wire _13964_;
wire _13965_;
wire _13966_;
wire _13967_;
wire _13968_;
wire _13969_;
wire _13970_;
wire _13971_;
wire _13972_;
wire _13973_;
wire _13974_;
wire _13975_;
wire _13976_;
wire _13977_;
wire _13978_;
wire _13979_;
wire _13980_;
wire _13981_;
wire _13982_;
wire _13983_;
wire _13984_;
wire _13985_;
wire _13986_;
wire _13987_;
wire _13988_;
wire _13989_;
wire _13990_;
wire _13991_;
wire _13992_;
wire _13993_;
wire _13994_;
wire _13995_;
wire _13996_;
wire _13997_;
wire _13998_;
wire _13999_;
wire _14000_;
wire _14001_;
wire _14002_;
wire _14003_;
wire _14004_;
wire _14005_;
wire _14006_;
wire _14007_;
wire _14008_;
wire _14009_;
wire _14010_;
wire _14011_;
wire _14012_;
wire _14013_;
wire _14014_;
wire _14015_;
wire _14016_;
wire _14017_;
wire _14018_;
wire _14019_;
wire _14020_;
wire _14021_;
wire _14022_;
wire _14023_;
wire _14024_;
wire _14025_;
wire _14026_;
wire _14027_;
wire _14028_;
wire _14029_;
wire _14030_;
wire _14031_;
wire _14032_;
wire _14033_;
wire _14034_;
wire _14035_;
wire _14036_;
wire _14037_;
wire _14038_;
wire _14039_;
wire _14040_;
wire _14041_;
wire _14042_;
wire _14043_;
wire _14044_;
wire _14045_;
wire _14046_;
wire _14047_;
wire _14048_;
wire _14049_;
wire _14050_;
wire _14051_;
wire _14052_;
wire _14053_;
wire _14054_;
wire _14055_;
wire _14056_;
wire _14057_;
wire _14058_;
wire _14059_;
wire _14060_;
wire _14061_;
wire _14062_;
wire _14063_;
wire _14064_;
wire _14065_;
wire _14066_;
wire _14067_;
wire _14068_;
wire _14069_;
wire _14070_;
wire _14071_;
wire _14072_;
wire _14073_;
wire _14074_;
wire _14075_;
wire _14076_;
wire _14077_;
wire _14078_;
wire _14079_;
wire _14080_;
wire _14081_;
wire _14082_;
wire _14083_;
wire _14084_;
wire _14085_;
wire _14086_;
wire _14087_;
wire _14088_;
wire _14089_;
wire _14090_;
wire _14091_;
wire _14092_;
wire _14093_;
wire _14094_;
wire _14095_;
wire _14096_;
wire _14097_;
wire _14098_;
wire _14099_;
wire _14100_;
wire _14101_;
wire _14102_;
wire _14103_;
wire _14104_;
wire _14105_;
wire _14106_;
wire _14107_;
wire _14108_;
wire _14109_;
wire _14110_;
wire _14111_;
wire _14112_;
wire _14113_;
wire _14114_;
wire _14115_;
wire _14116_;
wire _14117_;
wire _14118_;
wire _14119_;
wire _14120_;
wire _14121_;
wire _14122_;
wire _14123_;
wire _14124_;
wire _14125_;
wire _14126_;
wire _14127_;
wire _14128_;
wire _14129_;
wire _14130_;
wire _14131_;
wire _14132_;
wire _14133_;
wire _14134_;
wire _14135_;
wire _14136_;
wire _14137_;
wire _14138_;
wire _14139_;
wire _14140_;
wire _14141_;
wire _14142_;
wire _14143_;
wire _14144_;
wire _14145_;
wire _14146_;
wire _14147_;
wire _14148_;
wire _14149_;
wire _14150_;
wire _14151_;
wire _14152_;
wire _14153_;
wire _14154_;
wire _14155_;
wire _14156_;
wire _14157_;
wire _14158_;
wire _14159_;
wire _14160_;
wire _14161_;
wire _14162_;
wire _14163_;
wire _14164_;
wire _14165_;
wire _14166_;
wire _14167_;
wire _14168_;
wire _14169_;
wire _14170_;
wire _14171_;
wire _14172_;
wire _14173_;
wire _14174_;
wire _14175_;
wire _14176_;
wire _14177_;
wire _14178_;
wire _14179_;
wire _14180_;
wire _14181_;
wire _14182_;
wire _14183_;
wire _14184_;
wire _14185_;
wire _14186_;
wire _14187_;
wire _14188_;
wire _14189_;
wire _14190_;
wire _14191_;
wire _14192_;
wire _14193_;
wire _14194_;
wire _14195_;
wire _14196_;
wire _14197_;
wire _14198_;
wire _14199_;
wire _14200_;
wire _14201_;
wire _14202_;
wire _14203_;
wire _14204_;
wire _14205_;
wire _14206_;
wire _14207_;
wire _14208_;
wire _14209_;
wire _14210_;
wire _14211_;
wire _14212_;
wire _14213_;
wire _14214_;
wire _14215_;
wire _14216_;
wire _14217_;
wire _14218_;
wire _14219_;
wire _14220_;
wire _14221_;
wire _14222_;
wire _14223_;
wire _14224_;
wire _14225_;
wire _14226_;
wire _14227_;
wire _14228_;
wire _14229_;
wire _14230_;
wire _14231_;
wire _14232_;
wire _14233_;
wire _14234_;
wire _14235_;
wire _14236_;
wire _14237_;
wire _14238_;
wire _14239_;
wire _14240_;
wire _14241_;
wire _14242_;
wire _14243_;
wire _14244_;
wire _14245_;
wire _14246_;
wire _14247_;
wire _14248_;
wire _14249_;
wire _14250_;
wire _14251_;
wire _14252_;
wire _14253_;
wire _14254_;
wire _14255_;
wire _14256_;
wire _14257_;
wire _14258_;
wire _14259_;
wire _14260_;
wire _14261_;
wire _14262_;
wire _14263_;
wire _14264_;
wire _14265_;
wire _14266_;
wire _14267_;
wire _14268_;
wire _14269_;
wire _14270_;
wire _14271_;
wire _14272_;
wire _14273_;
wire _14274_;
wire _14275_;
wire _14276_;
wire _14277_;
wire _14278_;
wire _14279_;
wire _14280_;
wire _14281_;
wire _14282_;
wire _14283_;
wire _14284_;
wire _14285_;
wire _14286_;
wire _14287_;
wire _14288_;
wire _14289_;
wire _14290_;
wire _14291_;
wire _14292_;
wire _14293_;
wire _14294_;
wire _14295_;
wire _14296_;
wire _14297_;
wire _14298_;
wire _14299_;
wire _14300_;
wire _14301_;
wire _14302_;
wire _14303_;
wire _14304_;
wire _14305_;
wire _14306_;
wire _14307_;
wire _14308_;
wire _14309_;
wire _14310_;
wire _14311_;
wire _14312_;
wire _14313_;
wire _14314_;
wire _14315_;
wire _14316_;
wire _14317_;
wire _14318_;
wire _14319_;
wire _14320_;
wire _14321_;
wire _14322_;
wire _14323_;
wire _14324_;
wire _14325_;
wire _14326_;
wire _14327_;
wire _14328_;
wire _14329_;
wire _14330_;
wire _14331_;
wire _14332_;
wire _14333_;
wire _14334_;
wire _14335_;
wire _14336_;
wire _14337_;
wire _14338_;
wire _14339_;
wire _14340_;
wire _14341_;
wire _14342_;
wire _14343_;
wire _14344_;
wire _14345_;
wire _14346_;
wire _14347_;
wire _14348_;
wire _14349_;
wire _14350_;
wire _14351_;
wire _14352_;
wire _14353_;
wire _14354_;
wire _14355_;
wire _14356_;
wire _14357_;
wire _14358_;
wire _14359_;
wire _14360_;
wire _14361_;
wire _14362_;
wire _14363_;
wire _14364_;
wire _14365_;
wire _14366_;
wire _14367_;
wire _14368_;
wire _14369_;
wire _14370_;
wire _14371_;
wire _14372_;
wire _14373_;
wire _14374_;
wire _14375_;
wire _14376_;
wire _14377_;
wire _14378_;
wire _14379_;
wire _14380_;
wire _14381_;
wire _14382_;
wire _14383_;
wire _14384_;
wire _14385_;
wire _14386_;
wire _14387_;
wire _14388_;
wire _14389_;
wire _14390_;
wire _14391_;
wire _14392_;
wire _14393_;
wire _14394_;
wire _14395_;
wire _14396_;
wire _14397_;
wire _14398_;
wire _14399_;
wire _14400_;
wire _14401_;
wire _14402_;
wire _14403_;
wire _14404_;
wire _14405_;
wire _14406_;
wire _14407_;
wire _14408_;
wire _14409_;
wire _14410_;
wire _14411_;
wire _14412_;
wire _14413_;
wire _14414_;
wire _14415_;
wire _14416_;
wire _14417_;
wire _14418_;
wire _14419_;
wire _14420_;
wire _14421_;
wire _14422_;
wire _14423_;
wire _14424_;
wire _14425_;
wire _14426_;
wire _14427_;
wire _14428_;
wire _14429_;
wire _14430_;
wire _14431_;
wire _14432_;
wire _14433_;
wire _14434_;
wire _14435_;
wire _14436_;
wire _14437_;
wire _14438_;
wire _14439_;
wire _14440_;
wire _14441_;
wire _14442_;
wire _14443_;
wire _14444_;
wire _14445_;
wire _14446_;
wire _14447_;
wire _14448_;
wire _14449_;
wire _14450_;
wire _14451_;
wire _14452_;
wire _14453_;
wire _14454_;
wire _14455_;
wire _14456_;
wire _14457_;
wire _14458_;
wire _14459_;
wire _14460_;
wire _14461_;
wire _14462_;
wire _14463_;
wire _14464_;
wire _14465_;
wire _14466_;
wire _14467_;
wire _14468_;
wire _14469_;
wire _14470_;
wire _14471_;
wire _14472_;
wire _14473_;
wire _14474_;
wire _14475_;
wire _14476_;
wire _14477_;
wire _14478_;
wire _14479_;
wire _14480_;
wire _14481_;
wire _14482_;
wire _14483_;
wire _14484_;
wire _14485_;
wire _14486_;
wire _14487_;
wire _14488_;
wire _14489_;
wire _14490_;
wire _14491_;
wire _14492_;
wire _14493_;
wire _14494_;
wire _14495_;
wire _14496_;
wire _14497_;
wire _14498_;
wire _14499_;
wire _14500_;
wire _14501_;
wire _14502_;
wire _14503_;
wire _14504_;
wire _14505_;
wire _14506_;
wire _14507_;
wire _14508_;
wire _14509_;
wire _14510_;
wire _14511_;
wire _14512_;
wire _14513_;
wire _14514_;
wire _14515_;
wire _14516_;
wire _14517_;
wire _14518_;
wire _14519_;
wire _14520_;
wire _14521_;
wire _14522_;
wire _14523_;
wire _14524_;
wire _14525_;
wire _14526_;
wire _14527_;
wire _14528_;
wire _14529_;
wire _14530_;
wire _14531_;
wire _14532_;
wire _14533_;
wire _14534_;
wire _14535_;
wire _14536_;
wire _14537_;
wire _14538_;
wire _14539_;
wire _14540_;
wire _14541_;
wire _14542_;
wire _14543_;
wire _14544_;
wire _14545_;
wire _14546_;
wire _14547_;
wire _14548_;
wire _14549_;
wire _14550_;
wire _14551_;
wire _14552_;
wire _14553_;
wire _14554_;
wire _14555_;
wire _14556_;
wire _14557_;
wire _14558_;
wire _14559_;
wire _14560_;
wire _14561_;
wire _14562_;
wire _14563_;
wire _14564_;
wire _14565_;
wire _14566_;
wire _14567_;
wire _14568_;
wire _14569_;
wire _14570_;
wire _14571_;
wire _14572_;
wire _14573_;
wire _14574_;
wire _14575_;
wire _14576_;
wire _14577_;
wire _14578_;
wire _14579_;
wire _14580_;
wire _14581_;
wire _14582_;
wire _14583_;
wire _14584_;
wire _14585_;
wire _14586_;
wire _14587_;
wire _14588_;
wire _14589_;
wire _14590_;
wire _14591_;
wire _14592_;
wire _14593_;
wire _14594_;
wire _14595_;
wire _14596_;
wire _14597_;
wire _14598_;
wire _14599_;
wire _14600_;
wire _14601_;
wire _14602_;
wire _14603_;
wire _14604_;
wire _14605_;
wire _14606_;
wire _14607_;
wire _14608_;
wire _14609_;
wire _14610_;
wire _14611_;
wire _14612_;
wire _14613_;
wire _14614_;
wire _14615_;
wire _14616_;
wire _14617_;
wire _14618_;
wire _14619_;
wire _14620_;
wire _14621_;
wire _14622_;
wire _14623_;
wire _14624_;
wire _14625_;
wire _14626_;
wire _14627_;
wire _14628_;
wire _14629_;
wire _14630_;
wire _14631_;
wire _14632_;
wire _14633_;
wire _14634_;
wire _14635_;
wire _14636_;
wire _14637_;
wire _14638_;
wire _14639_;
wire _14640_;
wire _14641_;
wire _14642_;
wire _14643_;
wire _14644_;
wire _14645_;
wire _14646_;
wire _14647_;
wire _14648_;
wire _14649_;
wire _14650_;
wire _14651_;
wire _14652_;
wire _14653_;
wire _14654_;
wire _14655_;
wire _14656_;
wire _14657_;
wire _14658_;
wire _14659_;
wire _14660_;
wire _14661_;
wire _14662_;
wire _14663_;
wire _14664_;
wire _14665_;
wire _14666_;
wire _14667_;
wire _14668_;
wire _14669_;
wire _14670_;
wire _14671_;
wire _14672_;
wire _14673_;
wire _14674_;
wire _14675_;
wire _14676_;
wire _14677_;
wire _14678_;
wire _14679_;
wire _14680_;
wire _14681_;
wire _14682_;
wire _14683_;
wire _14684_;
wire _14685_;
wire _14686_;
wire _14687_;
wire _14688_;
wire _14689_;
wire _14690_;
wire _14691_;
wire _14692_;
wire _14693_;
wire _14694_;
wire _14695_;
wire _14696_;
wire _14697_;
wire _14698_;
wire _14699_;
wire _14700_;
wire _14701_;
wire _14702_;
wire _14703_;
wire _14704_;
wire _14705_;
wire _14706_;
wire _14707_;
wire _14708_;
wire _14709_;
wire _14710_;
wire _14711_;
wire _14712_;
wire _14713_;
wire _14714_;
wire _14715_;
wire _14716_;
wire _14717_;
wire _14718_;
wire _14719_;
wire _14720_;
wire _14721_;
wire _14722_;
wire _14723_;
wire _14724_;
wire _14725_;
wire _14726_;
wire _14727_;
wire _14728_;
wire _14729_;
wire _14730_;
wire _14731_;
wire _14732_;
wire _14733_;
wire _14734_;
wire _14735_;
wire _14736_;
wire _14737_;
wire _14738_;
wire _14739_;
wire _14740_;
wire _14741_;
wire _14742_;
wire _14743_;
wire _14744_;
wire _14745_;
wire _14746_;
wire _14747_;
wire _14748_;
wire _14749_;
wire _14750_;
wire _14751_;
wire _14752_;
wire _14753_;
wire _14754_;
wire _14755_;
wire _14756_;
wire _14757_;
wire _14758_;
wire _14759_;
wire _14760_;
wire _14761_;
wire _14762_;
wire _14763_;
wire _14764_;
wire _14765_;
wire _14766_;
wire _14767_;
wire _14768_;
wire _14769_;
wire _14770_;
wire _14771_;
wire _14772_;
wire _14773_;
wire _14774_;
wire _14775_;
wire _14776_;
wire _14777_;
wire _14778_;
wire _14779_;
wire _14780_;
wire _14781_;
wire _14782_;
wire _14783_;
wire _14784_;
wire _14785_;
wire _14786_;
wire _14787_;
wire _14788_;
wire _14789_;
wire _14790_;
wire _14791_;
wire _14792_;
wire _14793_;
wire _14794_;
wire _14795_;
wire _14796_;
wire _14797_;
wire _14798_;
wire _14799_;
wire _14800_;
wire _14801_;
wire _14802_;
wire _14803_;
wire _14804_;
wire _14805_;
wire _14806_;
wire _14807_;
wire _14808_;
wire _14809_;
wire _14810_;
wire _14811_;
wire _14812_;
wire _14813_;
wire _14814_;
wire _14815_;
wire _14816_;
wire _14817_;
wire _14818_;
wire _14819_;
wire _14820_;
wire _14821_;
wire _14822_;
wire _14823_;
wire _14824_;
wire _14825_;
wire _14826_;
wire _14827_;
wire _14828_;
wire _14829_;
wire _14830_;
wire _14831_;
wire _14832_;
wire _14833_;
wire _14834_;
wire _14835_;
wire _14836_;
wire _14837_;
wire _14838_;
wire _14839_;
wire _14840_;
wire _14841_;
wire _14842_;
wire _14843_;
wire _14844_;
wire _14845_;
wire _14846_;
wire _14847_;
wire _14848_;
wire _14849_;
wire _14850_;
wire _14851_;
wire _14852_;
wire _14853_;
wire _14854_;
wire _14855_;
wire _14856_;
wire _14857_;
wire _14858_;
wire _14859_;
wire _14860_;
wire _14861_;
wire _14862_;
wire _14863_;
wire _14864_;
wire _14865_;
wire _14866_;
wire _14867_;
wire _14868_;
wire _14869_;
wire _14870_;
wire _14871_;
wire _14872_;
wire _14873_;
wire _14874_;
wire _14875_;
wire _14876_;
wire _14877_;
wire _14878_;
wire _14879_;
wire _14880_;
wire _14881_;
wire _14882_;
wire _14883_;
wire _14884_;
wire _14885_;
wire _14886_;
wire _14887_;
wire _14888_;
wire _14889_;
wire _14890_;
wire _14891_;
wire _14892_;
wire _14893_;
wire _14894_;
wire _14895_;
wire _14896_;
wire _14897_;
wire _14898_;
wire _14899_;
wire _14900_;
wire _14901_;
wire _14902_;
wire _14903_;
wire _14904_;
wire _14905_;
wire _14906_;
wire _14907_;
wire _14908_;
wire _14909_;
wire _14910_;
wire _14911_;
wire _14912_;
wire _14913_;
wire _14914_;
wire _14915_;
wire _14916_;
wire _14917_;
wire _14918_;
wire _14919_;
wire _14920_;
wire _14921_;
wire _14922_;
wire _14923_;
wire _14924_;
wire _14925_;
wire _14926_;
wire _14927_;
wire _14928_;
wire _14929_;
wire _14930_;
wire _14931_;
wire _14932_;
wire _14933_;
wire _14934_;
wire _14935_;
wire _14936_;
wire _14937_;
wire _14938_;
wire _14939_;
wire _14940_;
wire _14941_;
wire _14942_;
wire _14943_;
wire _14944_;
wire _14945_;
wire _14946_;
wire _14947_;
wire _14948_;
wire _14949_;
wire _14950_;
wire _14951_;
wire _14952_;
wire _14953_;
wire _14954_;
wire _14955_;
wire _14956_;
wire _14957_;
wire _14958_;
wire _14959_;
wire _14960_;
wire _14961_;
wire _14962_;
wire _14963_;
wire _14964_;
wire _14965_;
wire _14966_;
wire _14967_;
wire _14968_;
wire _14969_;
wire _14970_;
wire _14971_;
wire _14972_;
wire _14973_;
wire _14974_;
wire _14975_;
wire _14976_;
wire _14977_;
wire _14978_;
wire _14979_;
wire _14980_;
wire _14981_;
wire _14982_;
wire _14983_;
wire _14984_;
wire _14985_;
wire _14986_;
wire _14987_;
wire _14988_;
wire _14989_;
wire _14990_;
wire _14991_;
wire _14992_;
wire _14993_;
wire _14994_;
wire _14995_;
wire _14996_;
wire _14997_;
wire _14998_;
wire [31:0] alu_out;
wire [31:0] alu_out_q;
input clk;
wire clk;
wire [63:0] count_cycle;
wire [63:0] count_instr;
wire [7:0] cpu_state;
wire [31:0] cpuregs[0];
wire [31:0] cpuregs[10];
wire [31:0] cpuregs[11];
wire [31:0] cpuregs[12];
wire [31:0] cpuregs[13];
wire [31:0] cpuregs[14];
wire [31:0] cpuregs[15];
wire [31:0] cpuregs[16];
wire [31:0] cpuregs[17];
wire [31:0] cpuregs[18];
wire [31:0] cpuregs[19];
wire [31:0] cpuregs[1];
wire [31:0] cpuregs[20];
wire [31:0] cpuregs[21];
wire [31:0] cpuregs[22];
wire [31:0] cpuregs[23];
wire [31:0] cpuregs[24];
wire [31:0] cpuregs[25];
wire [31:0] cpuregs[26];
wire [31:0] cpuregs[27];
wire [31:0] cpuregs[28];
wire [31:0] cpuregs[29];
wire [31:0] cpuregs[2];
wire [31:0] cpuregs[30];
wire [31:0] cpuregs[31];
wire [31:0] cpuregs[3];
wire [31:0] cpuregs[4];
wire [31:0] cpuregs[5];
wire [31:0] cpuregs[6];
wire [31:0] cpuregs[7];
wire [31:0] cpuregs[8];
wire [31:0] cpuregs[9];
wire [31:0] decoded_imm;
wire [31:0] decoded_imm_j;
wire [4:0] decoded_rd;
wire decoder_pseudo_trigger;
wire decoder_trigger;
output [31:0] eoi;
wire [31:0] eoi;
wire instr_add;
wire instr_addi;
wire instr_and;
wire instr_andi;
wire instr_auipc;
wire instr_beq;
wire instr_bge;
wire instr_bgeu;
wire instr_blt;
wire instr_bltu;
wire instr_bne;
wire instr_jal;
wire instr_jalr;
wire instr_lb;
wire instr_lbu;
wire instr_lh;
wire instr_lhu;
wire instr_lui;
wire instr_lw;
wire instr_or;
wire instr_ori;
wire instr_rdcycle;
wire instr_rdcycleh;
wire instr_rdinstr;
wire instr_rdinstrh;
wire instr_sb;
wire instr_sh;
wire instr_sll;
wire instr_slli;
wire instr_slt;
wire instr_slti;
wire instr_sltiu;
wire instr_sltu;
wire instr_sra;
wire instr_srai;
wire instr_srl;
wire instr_srli;
wire instr_sub;
wire instr_sw;
wire instr_xor;
wire instr_xori;
input [31:0] irq;
wire [31:0] irq;
wire is_alu_reg_imm;
wire is_alu_reg_reg;
wire is_beq_bne_blt_bge_bltu_bgeu;
wire is_compare;
wire is_jalr_addi_slti_sltiu_xori_ori_andi;
wire is_lb_lh_lw_lbu_lhu;
wire is_lbu_lhu_lw;
wire is_lui_auipc_jal;
wire is_lui_auipc_jal_jalr_addi_add_sub;
wire is_sb_sh_sw;
wire is_sll_srl_sra;
wire is_slli_srli_srai;
wire is_slti_blt_slt;
wire is_sltiu_bltu_sltu;
wire latched_branch;
wire latched_is_lb;
wire latched_is_lh;
wire latched_is_lu;
wire [4:0] latched_rd;
wire latched_stalu;
wire latched_store;
output [31:0] mem_addr;
wire [31:0] mem_addr;
wire mem_do_prefetch;
wire mem_do_rdata;
wire mem_do_rinst;
wire mem_do_wdata;
output mem_instr;
wire mem_instr;
output [31:0] mem_la_addr;
wire [31:0] mem_la_addr;
output mem_la_read;
wire mem_la_read;
output [31:0] mem_la_wdata;
wire [31:0] mem_la_wdata;
output mem_la_write;
wire mem_la_write;
output [3:0] mem_la_wstrb;
wire [3:0] mem_la_wstrb;
input [31:0] mem_rdata;
wire [31:0] mem_rdata;
wire [31:0] mem_rdata_q;
input mem_ready;
wire mem_ready;
wire [1:0] mem_state;
output mem_valid;
wire mem_valid;
output [31:0] mem_wdata;
wire [31:0] mem_wdata;
wire [1:0] mem_wordsize;
output [3:0] mem_wstrb;
wire [3:0] mem_wstrb;
output [31:0] pcpi_insn;
wire [31:0] pcpi_insn;
input [31:0] pcpi_rd;
wire [31:0] pcpi_rd;
input pcpi_ready;
wire pcpi_ready;
output [31:0] pcpi_rs1;
wire [31:0] pcpi_rs1;
output [31:0] pcpi_rs2;
wire [31:0] pcpi_rs2;
output pcpi_valid;
wire pcpi_valid;
input pcpi_wait;
wire pcpi_wait;
input pcpi_wr;
wire pcpi_wr;
wire [31:0] reg_next_pc;
wire [31:0] reg_out;
wire [31:0] reg_pc;
wire [4:0] reg_sh;
input resetn;
wire resetn;
output [35:0] trace_data;
wire [35:0] trace_data;
output trace_valid;
wire trace_valid;
output trap;
wire trap;
NOT_g _14999_ (.A(count_instr[62]), .Y(_08761_));
NOT_g _15000_ (.A(count_instr[60]), .Y(_08762_));
NOT_g _15001_ (.A(count_instr[58]), .Y(_08763_));
NOT_g _15002_ (.A(count_instr[54]), .Y(_08764_));
NOT_g _15003_ (.A(count_instr[52]), .Y(_08765_));
NOT_g _15004_ (.A(count_instr[49]), .Y(_08766_));
NOT_g _15005_ (.A(count_instr[47]), .Y(_08767_));
NOT_g _15006_ (.A(count_instr[46]), .Y(_08768_));
NOT_g _15007_ (.A(count_instr[45]), .Y(_08769_));
NOT_g _15008_ (.A(count_instr[41]), .Y(_08770_));
NOT_g _15009_ (.A(count_instr[39]), .Y(_08771_));
NOT_g _15010_ (.A(count_instr[37]), .Y(_08772_));
NOT_g _15011_ (.A(count_instr[35]), .Y(_08773_));
NOT_g _15012_ (.A(count_instr[30]), .Y(_08774_));
NOT_g _15013_ (.A(count_instr[28]), .Y(_08775_));
NOT_g _15014_ (.A(count_instr[25]), .Y(_08776_));
NOT_g _15015_ (.A(count_instr[22]), .Y(_08777_));
NOT_g _15016_ (.A(count_instr[19]), .Y(_08778_));
NOT_g _15017_ (.A(count_instr[17]), .Y(_08779_));
NOT_g _15018_ (.A(count_instr[15]), .Y(_08780_));
NOT_g _15019_ (.A(count_instr[14]), .Y(_08781_));
NOT_g _15020_ (.A(count_instr[13]), .Y(_08782_));
NOT_g _15021_ (.A(count_instr[12]), .Y(_08783_));
NOT_g _15022_ (.A(count_instr[11]), .Y(_08784_));
NOT_g _15023_ (.A(count_instr[8]), .Y(_08785_));
NOT_g _15024_ (.A(count_instr[5]), .Y(_08786_));
NOT_g _15025_ (.A(count_instr[3]), .Y(_08787_));
NOT_g _15026_ (.A(count_instr[1]), .Y(_08788_));
NOT_g _15027_ (.A(mem_do_wdata), .Y(_08789_));
NOT_g _15028_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .Y(_08790_));
NOT_g _15029_ (.A(instr_sra), .Y(_08791_));
NOT_g _15030_ (.A(instr_xor), .Y(_08792_));
NOT_g _15031_ (.A(instr_sll), .Y(_08793_));
NOT_g _15032_ (.A(instr_sub), .Y(_08794_));
NOT_g _15033_ (.A(instr_xori), .Y(_08795_));
NOT_g _15034_ (.A(instr_addi), .Y(_08796_));
NOT_g _15035_ (.A(instr_bltu), .Y(_08797_));
NOT_g _15036_ (.A(instr_blt), .Y(_08798_));
NOT_g _15037_ (.A(latched_is_lh), .Y(_08799_));
NOT_g _15038_ (.A(latched_is_lu), .Y(_08800_));
NOT_g _15039_ (.A(latched_branch), .Y(_08801_));
NOT_g _15040_ (.A(latched_stalu), .Y(_08802_));
NOT_g _15041_ (.A(mem_do_rdata), .Y(_08803_));
NOT_g _15042_ (.A(mem_do_rinst), .Y(_08804_));
NOT_g _15043_ (.A(reg_pc[31]), .Y(_08805_));
NOT_g _15044_ (.A(reg_pc[2]), .Y(_08806_));
NOT_g _15045_ (.A(mem_do_prefetch), .Y(_08807_));
NOT_g _15046_ (.A(cpuregs[15][2]), .Y(_08808_));
NOT_g _15047_ (.A(cpuregs[15][19]), .Y(_08809_));
NOT_g _15048_ (.A(cpuregs[15][20]), .Y(_08810_));
NOT_g _15049_ (.A(resetn), .Y(_08811_));
NOT_g _15050_ (.A(pcpi_rs2[1]), .Y(_08812_));
NOT_g _15051_ (.A(pcpi_rs2[2]), .Y(_08813_));
NOT_g _15052_ (.A(pcpi_rs2[4]), .Y(_08814_));
NOT_g _15053_ (.A(pcpi_rs2[5]), .Y(_08815_));
NOT_g _15054_ (.A(pcpi_rs2[6]), .Y(_08816_));
NOT_g _15055_ (.A(pcpi_rs2[7]), .Y(_08817_));
NOT_g _15056_ (.A(pcpi_rs2[8]), .Y(_08818_));
NOT_g _15057_ (.A(pcpi_rs2[9]), .Y(_08819_));
NOT_g _15058_ (.A(pcpi_rs2[10]), .Y(_08820_));
NOT_g _15059_ (.A(pcpi_rs2[11]), .Y(_08821_));
NOT_g _15060_ (.A(pcpi_rs2[12]), .Y(_08822_));
NOT_g _15061_ (.A(pcpi_rs2[13]), .Y(_08823_));
NOT_g _15062_ (.A(pcpi_rs2[14]), .Y(_08824_));
NOT_g _15063_ (.A(pcpi_rs2[15]), .Y(_08825_));
NOT_g _15064_ (.A(pcpi_rs2[16]), .Y(_08826_));
NOT_g _15065_ (.A(pcpi_rs2[17]), .Y(_08827_));
NOT_g _15066_ (.A(pcpi_rs2[18]), .Y(_08828_));
NOT_g _15067_ (.A(pcpi_rs2[19]), .Y(_08829_));
NOT_g _15068_ (.A(pcpi_rs2[20]), .Y(_08830_));
NOT_g _15069_ (.A(pcpi_rs2[21]), .Y(_08831_));
NOT_g _15070_ (.A(pcpi_rs2[22]), .Y(_08832_));
NOT_g _15071_ (.A(pcpi_rs2[23]), .Y(_08833_));
NOT_g _15072_ (.A(pcpi_rs2[24]), .Y(_08834_));
NOT_g _15073_ (.A(pcpi_rs2[25]), .Y(_08835_));
NOT_g _15074_ (.A(pcpi_rs2[26]), .Y(_08836_));
NOT_g _15075_ (.A(pcpi_rs2[27]), .Y(_08837_));
NOT_g _15076_ (.A(pcpi_rs2[28]), .Y(_08838_));
NOT_g _15077_ (.A(pcpi_rs2[29]), .Y(_08839_));
NOT_g _15078_ (.A(pcpi_rs2[30]), .Y(_08840_));
NOT_g _15079_ (.A(pcpi_rs2[31]), .Y(_08841_));
NOT_g _15080_ (.A(mem_wordsize[0]), .Y(_08842_));
NOT_g _15081_ (.A(mem_wordsize[1]), .Y(_08843_));
NOT_g _15082_ (.A(cpuregs[20][6]), .Y(_08844_));
NOT_g _15083_ (.A(cpuregs[20][11]), .Y(_08845_));
NOT_g _15084_ (.A(cpuregs[20][12]), .Y(_08846_));
NOT_g _15085_ (.A(cpuregs[20][14]), .Y(_08847_));
NOT_g _15086_ (.A(cpuregs[20][15]), .Y(_08848_));
NOT_g _15087_ (.A(cpuregs[20][16]), .Y(_08849_));
NOT_g _15088_ (.A(cpuregs[20][23]), .Y(_08850_));
NOT_g _15089_ (.A(cpuregs[20][25]), .Y(_08851_));
NOT_g _15090_ (.A(latched_rd[1]), .Y(_08852_));
NOT_g _15091_ (.A(latched_rd[2]), .Y(_08853_));
NOT_g _15092_ (.A(latched_rd[3]), .Y(_08854_));
NOT_g _15093_ (.A(instr_lui), .Y(_08855_));
NOT_g _15094_ (.A(instr_auipc), .Y(_08856_));
NOT_g _15095_ (.A(instr_jal), .Y(_08857_));
NOT_g _15096_ (.A(instr_lhu), .Y(_08858_));
NOT_g _15097_ (.A(instr_slli), .Y(_08859_));
NOT_g _15098_ (.A(instr_srai), .Y(_08860_));
NOT_g _15099_ (.A(is_slli_srli_srai), .Y(_08861_));
NOT_g _15100_ (.A(is_sll_srl_sra), .Y(_08862_));
NOT_g _15101_ (.A(is_alu_reg_imm), .Y(_08863_));
NOT_g _15102_ (.A(is_sb_sh_sw), .Y(_08864_));
NOT_g _15103_ (.A(mem_rdata_q[12]), .Y(_08865_));
NOT_g _15104_ (.A(mem_rdata_q[13]), .Y(_08866_));
NOT_g _15105_ (.A(mem_rdata_q[14]), .Y(_08867_));
NOT_g _15106_ (.A(mem_rdata_q[20]), .Y(_08868_));
NOT_g _15107_ (.A(mem_rdata_q[27]), .Y(_08869_));
NOT_g _15108_ (.A(mem_rdata_q[29]), .Y(_08870_));
NOT_g _15109_ (.A(mem_rdata_q[30]), .Y(_08871_));
NOT_g _15110_ (.A(mem_rdata_q[31]), .Y(_08872_));
NOT_g _15111_ (.A(mem_state[1]), .Y(_08873_));
NOT_g _15112_ (.A(mem_rdata_q[2]), .Y(_08874_));
NOT_g _15113_ (.A(mem_rdata_q[3]), .Y(_08875_));
NOT_g _15114_ (.A(cpuregs[29][2]), .Y(_08876_));
NOT_g _15115_ (.A(cpuregs[29][4]), .Y(_08877_));
NOT_g _15116_ (.A(cpuregs[29][18]), .Y(_08878_));
NOT_g _15117_ (.A(decoded_imm_j[4]), .Y(_08879_));
NOT_g _15118_ (.A(cpuregs[12][6]), .Y(_08880_));
NOT_g _15119_ (.A(cpuregs[12][10]), .Y(_08881_));
NOT_g _15120_ (.A(cpuregs[12][23]), .Y(_08882_));
NOT_g _15121_ (.A(cpuregs[12][25]), .Y(_08883_));
NOT_g _15122_ (.A(cpuregs[12][30]), .Y(_08884_));
NOT_g _15123_ (.A(cpuregs[23][1]), .Y(_08885_));
NOT_g _15124_ (.A(cpuregs[23][6]), .Y(_08886_));
NOT_g _15125_ (.A(cpuregs[23][8]), .Y(_08887_));
NOT_g _15126_ (.A(cpuregs[23][9]), .Y(_08888_));
NOT_g _15127_ (.A(cpuregs[23][10]), .Y(_08889_));
NOT_g _15128_ (.A(cpuregs[23][11]), .Y(_08890_));
NOT_g _15129_ (.A(cpuregs[23][12]), .Y(_08891_));
NOT_g _15130_ (.A(cpuregs[23][14]), .Y(_08892_));
NOT_g _15131_ (.A(cpuregs[23][15]), .Y(_08893_));
NOT_g _15132_ (.A(cpuregs[23][16]), .Y(_08894_));
NOT_g _15133_ (.A(cpuregs[23][19]), .Y(_08895_));
NOT_g _15134_ (.A(cpuregs[23][20]), .Y(_08896_));
NOT_g _15135_ (.A(cpuregs[23][21]), .Y(_08897_));
NOT_g _15136_ (.A(cpuregs[23][22]), .Y(_08898_));
NOT_g _15137_ (.A(cpuregs[23][23]), .Y(_08899_));
NOT_g _15138_ (.A(cpuregs[23][25]), .Y(_08900_));
NOT_g _15139_ (.A(cpuregs[23][27]), .Y(_08901_));
NOT_g _15140_ (.A(cpuregs[23][28]), .Y(_08902_));
NOT_g _15141_ (.A(cpuregs[23][30]), .Y(_08903_));
NOT_g _15142_ (.A(cpuregs[4][0]), .Y(_08904_));
NOT_g _15143_ (.A(cpuregs[4][6]), .Y(_08905_));
NOT_g _15144_ (.A(cpuregs[4][8]), .Y(_08906_));
NOT_g _15145_ (.A(cpuregs[4][9]), .Y(_08907_));
NOT_g _15146_ (.A(cpuregs[4][11]), .Y(_08908_));
NOT_g _15147_ (.A(cpuregs[4][12]), .Y(_08909_));
NOT_g _15148_ (.A(cpuregs[4][14]), .Y(_08910_));
NOT_g _15149_ (.A(cpuregs[4][15]), .Y(_08911_));
NOT_g _15150_ (.A(cpuregs[4][16]), .Y(_08912_));
NOT_g _15151_ (.A(cpuregs[4][18]), .Y(_08913_));
NOT_g _15152_ (.A(cpuregs[4][19]), .Y(_08914_));
NOT_g _15153_ (.A(cpuregs[4][20]), .Y(_08915_));
NOT_g _15154_ (.A(cpuregs[4][21]), .Y(_08916_));
NOT_g _15155_ (.A(cpuregs[4][28]), .Y(_08917_));
NOT_g _15156_ (.A(cpuregs[22][6]), .Y(_08918_));
NOT_g _15157_ (.A(cpuregs[22][11]), .Y(_08919_));
NOT_g _15158_ (.A(cpuregs[22][12]), .Y(_08920_));
NOT_g _15159_ (.A(cpuregs[22][14]), .Y(_08921_));
NOT_g _15160_ (.A(cpuregs[22][15]), .Y(_08922_));
NOT_g _15161_ (.A(cpuregs[22][16]), .Y(_08923_));
NOT_g _15162_ (.A(cpuregs[22][23]), .Y(_08924_));
NOT_g _15163_ (.A(cpuregs[22][25]), .Y(_08925_));
NOT_g _15164_ (.A(cpuregs[13][2]), .Y(_08926_));
NOT_g _15165_ (.A(cpuregs[13][4]), .Y(_08927_));
NOT_g _15166_ (.A(cpuregs[13][6]), .Y(_08928_));
NOT_g _15167_ (.A(cpuregs[13][10]), .Y(_08929_));
NOT_g _15168_ (.A(cpuregs[13][19]), .Y(_08930_));
NOT_g _15169_ (.A(cpuregs[13][20]), .Y(_08931_));
NOT_g _15170_ (.A(cpuregs[13][23]), .Y(_08932_));
NOT_g _15171_ (.A(cpuregs[13][25]), .Y(_08933_));
NOT_g _15172_ (.A(cpuregs[13][26]), .Y(_08934_));
NOT_g _15173_ (.A(cpuregs[13][30]), .Y(_08935_));
NOT_g _15174_ (.A(cpuregs[18][10]), .Y(_08936_));
NOT_g _15175_ (.A(cpuregs[18][22]), .Y(_08937_));
NOT_g _15176_ (.A(cpuregs[18][27]), .Y(_08938_));
NOT_g _15177_ (.A(cpuregs[14][19]), .Y(_08939_));
NOT_g _15178_ (.A(cpuregs[14][20]), .Y(_08940_));
NOT_g _15179_ (.A(cpuregs[17][6]), .Y(_08941_));
NOT_g _15180_ (.A(cpuregs[17][12]), .Y(_08942_));
NOT_g _15181_ (.A(cpuregs[17][14]), .Y(_08943_));
NOT_g _15182_ (.A(cpuregs[17][16]), .Y(_08944_));
NOT_g _15183_ (.A(decoded_imm_j[19]), .Y(_08945_));
NOT_g _15184_ (.A(cpuregs[5][0]), .Y(_08946_));
NOT_g _15185_ (.A(cpuregs[5][6]), .Y(_08947_));
NOT_g _15186_ (.A(cpuregs[5][8]), .Y(_08948_));
NOT_g _15187_ (.A(cpuregs[5][9]), .Y(_08949_));
NOT_g _15188_ (.A(cpuregs[5][11]), .Y(_08950_));
NOT_g _15189_ (.A(cpuregs[5][12]), .Y(_08951_));
NOT_g _15190_ (.A(cpuregs[5][14]), .Y(_08952_));
NOT_g _15191_ (.A(cpuregs[5][15]), .Y(_08953_));
NOT_g _15192_ (.A(cpuregs[5][16]), .Y(_08954_));
NOT_g _15193_ (.A(cpuregs[5][18]), .Y(_08955_));
NOT_g _15194_ (.A(cpuregs[5][19]), .Y(_08956_));
NOT_g _15195_ (.A(cpuregs[5][20]), .Y(_08957_));
NOT_g _15196_ (.A(cpuregs[5][21]), .Y(_08958_));
NOT_g _15197_ (.A(cpuregs[5][24]), .Y(_08959_));
NOT_g _15198_ (.A(cpuregs[5][28]), .Y(_08960_));
NOT_g _15199_ (.A(pcpi_rs1[0]), .Y(_08961_));
NOT_g _15200_ (.A(pcpi_rs1[7]), .Y(_08962_));
NOT_g _15201_ (.A(cpuregs[7][0]), .Y(_08963_));
NOT_g _15202_ (.A(cpuregs[7][6]), .Y(_08964_));
NOT_g _15203_ (.A(cpuregs[7][8]), .Y(_08965_));
NOT_g _15204_ (.A(cpuregs[7][9]), .Y(_08966_));
NOT_g _15205_ (.A(cpuregs[7][11]), .Y(_08967_));
NOT_g _15206_ (.A(cpuregs[7][12]), .Y(_08968_));
NOT_g _15207_ (.A(cpuregs[7][14]), .Y(_08969_));
NOT_g _15208_ (.A(cpuregs[7][15]), .Y(_08970_));
NOT_g _15209_ (.A(cpuregs[7][16]), .Y(_08971_));
NOT_g _15210_ (.A(cpuregs[7][18]), .Y(_08972_));
NOT_g _15211_ (.A(cpuregs[7][19]), .Y(_08973_));
NOT_g _15212_ (.A(cpuregs[7][20]), .Y(_08974_));
NOT_g _15213_ (.A(cpuregs[7][21]), .Y(_08975_));
NOT_g _15214_ (.A(cpuregs[7][22]), .Y(_08976_));
NOT_g _15215_ (.A(cpuregs[7][24]), .Y(_08977_));
NOT_g _15216_ (.A(cpuregs[7][27]), .Y(_08978_));
NOT_g _15217_ (.A(cpuregs[7][28]), .Y(_08979_));
NOT_g _15218_ (.A(cpuregs[9][10]), .Y(_08980_));
NOT_g _15219_ (.A(cpuregs[9][25]), .Y(_08981_));
NOT_g _15220_ (.A(cpuregs[21][1]), .Y(_08982_));
NOT_g _15221_ (.A(cpuregs[21][2]), .Y(_08983_));
NOT_g _15222_ (.A(cpuregs[21][4]), .Y(_08984_));
NOT_g _15223_ (.A(cpuregs[21][6]), .Y(_08985_));
NOT_g _15224_ (.A(cpuregs[21][8]), .Y(_08986_));
NOT_g _15225_ (.A(cpuregs[21][9]), .Y(_08987_));
NOT_g _15226_ (.A(cpuregs[21][10]), .Y(_08988_));
NOT_g _15227_ (.A(cpuregs[21][11]), .Y(_08989_));
NOT_g _15228_ (.A(cpuregs[21][12]), .Y(_08990_));
NOT_g _15229_ (.A(cpuregs[21][14]), .Y(_08991_));
NOT_g _15230_ (.A(cpuregs[21][15]), .Y(_08992_));
NOT_g _15231_ (.A(cpuregs[21][16]), .Y(_08993_));
NOT_g _15232_ (.A(cpuregs[21][19]), .Y(_08994_));
NOT_g _15233_ (.A(cpuregs[21][20]), .Y(_08995_));
NOT_g _15234_ (.A(cpuregs[21][21]), .Y(_08996_));
NOT_g _15235_ (.A(cpuregs[21][22]), .Y(_08997_));
NOT_g _15236_ (.A(cpuregs[21][23]), .Y(_08998_));
NOT_g _15237_ (.A(cpuregs[21][25]), .Y(_08999_));
NOT_g _15238_ (.A(cpuregs[21][27]), .Y(_09000_));
NOT_g _15239_ (.A(cpuregs[21][28]), .Y(_09001_));
NOT_g _15240_ (.A(cpuregs[21][30]), .Y(_09002_));
NOT_g _15241_ (.A(cpuregs[6][0]), .Y(_09003_));
NOT_g _15242_ (.A(cpuregs[6][6]), .Y(_09004_));
NOT_g _15243_ (.A(cpuregs[6][8]), .Y(_09005_));
NOT_g _15244_ (.A(cpuregs[6][9]), .Y(_09006_));
NOT_g _15245_ (.A(cpuregs[6][11]), .Y(_09007_));
NOT_g _15246_ (.A(cpuregs[6][12]), .Y(_09008_));
NOT_g _15247_ (.A(cpuregs[6][14]), .Y(_09009_));
NOT_g _15248_ (.A(cpuregs[6][15]), .Y(_09010_));
NOT_g _15249_ (.A(cpuregs[6][16]), .Y(_09011_));
NOT_g _15250_ (.A(cpuregs[6][18]), .Y(_09012_));
NOT_g _15251_ (.A(cpuregs[6][19]), .Y(_09013_));
NOT_g _15252_ (.A(cpuregs[6][20]), .Y(_09014_));
NOT_g _15253_ (.A(cpuregs[6][21]), .Y(_09015_));
NOT_g _15254_ (.A(cpuregs[6][28]), .Y(_09016_));
NOT_g _15255_ (.A(decoded_imm_j[31]), .Y(_09017_));
NOT_g _15256_ (.A(cpu_state[6]), .Y(_09018_));
NOT_g _15257_ (.A(cpu_state[2]), .Y(_09019_));
NOT_g _15258_ (.A(cpu_state[4]), .Y(_09020_));
NOT_g _15259_ (.A(reg_sh[0]), .Y(_09021_));
NOT_g _15260_ (.A(reg_sh[4]), .Y(_09022_));
NOT_g _15261_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(_09023_));
NOT_g _15262_ (.A(decoder_pseudo_trigger), .Y(_09024_));
NOT_g _15263_ (.A(_00007_[0]), .Y(_09025_));
NOT_g _15264_ (.A(_00007_[1]), .Y(_09026_));
NOT_g _15265_ (.A(_00007_[2]), .Y(_09027_));
NOT_g _15266_ (.A(_00007_[3]), .Y(_09028_));
NOT_g _15267_ (.A(_00007_[4]), .Y(_09029_));
NOT_g _15268_ (.A(_00008_[0]), .Y(_09030_));
NOT_g _15269_ (.A(_00008_[1]), .Y(_09031_));
NOT_g _15270_ (.A(_00008_[2]), .Y(_09032_));
NOT_g _15271_ (.A(_00008_[3]), .Y(_09033_));
NOT_g _15272_ (.A(count_cycle[2]), .Y(_09034_));
NOT_g _15273_ (.A(count_cycle[4]), .Y(_09035_));
NOT_g _15274_ (.A(count_cycle[6]), .Y(_09036_));
NOT_g _15275_ (.A(count_cycle[8]), .Y(_09037_));
NOT_g _15276_ (.A(count_cycle[10]), .Y(_09038_));
NOT_g _15277_ (.A(count_cycle[12]), .Y(_09039_));
NOT_g _15278_ (.A(count_cycle[14]), .Y(_09040_));
NOT_g _15279_ (.A(count_cycle[16]), .Y(_09041_));
NOT_g _15280_ (.A(count_cycle[18]), .Y(_09042_));
NOT_g _15281_ (.A(count_cycle[20]), .Y(_09043_));
NOT_g _15282_ (.A(count_cycle[22]), .Y(_09044_));
NOT_g _15283_ (.A(count_cycle[24]), .Y(_09045_));
NOT_g _15284_ (.A(count_cycle[26]), .Y(_09046_));
NOT_g _15285_ (.A(count_cycle[28]), .Y(_09047_));
NOT_g _15286_ (.A(count_cycle[30]), .Y(_09048_));
NOT_g _15287_ (.A(count_cycle[32]), .Y(_09049_));
NOT_g _15288_ (.A(count_cycle[34]), .Y(_09050_));
NOT_g _15289_ (.A(count_cycle[36]), .Y(_09051_));
NOT_g _15290_ (.A(count_cycle[38]), .Y(_09052_));
NOT_g _15291_ (.A(count_cycle[40]), .Y(_09053_));
NOT_g _15292_ (.A(count_cycle[42]), .Y(_09054_));
NOT_g _15293_ (.A(count_cycle[44]), .Y(_09055_));
NOT_g _15294_ (.A(count_cycle[46]), .Y(_09056_));
NOT_g _15295_ (.A(count_cycle[48]), .Y(_09057_));
NOT_g _15296_ (.A(count_cycle[50]), .Y(_09058_));
NOT_g _15297_ (.A(count_cycle[52]), .Y(_09059_));
NOT_g _15298_ (.A(count_cycle[54]), .Y(_09060_));
NOT_g _15299_ (.A(count_cycle[56]), .Y(_09061_));
NOT_g _15300_ (.A(count_cycle[58]), .Y(_09062_));
NOT_g _15301_ (.A(count_cycle[60]), .Y(_09063_));
NOT_g _15302_ (.A(count_cycle[62]), .Y(_09064_));
NOR_g _15303_ (.A(latched_branch), .B(latched_store), .Y(_09065_));
NOT_g _15304_ (.A(_09065_), .Y(_09066_));
NOR_g _15305_ (.A(cpu_state[0]), .B(cpu_state[1]), .Y(_09067_));
NOR_g _15306_ (.A(cpu_state[2]), .B(cpu_state[3]), .Y(_09068_));
AND_g _15307_ (.A(_09067_), .B(_09068_), .Y(_09069_));
NOR_g _15308_ (.A(cpu_state[5]), .B(cpu_state[4]), .Y(_09070_));
NOR_g _15309_ (.A(_09018_), .B(cpu_state[7]), .Y(_09071_));
AND_g _15310_ (.A(_09070_), .B(_09071_), .Y(_09072_));
AND_g _15311_ (.A(_09069_), .B(_09072_), .Y(_09073_));
NAND_g _15312_ (.A(_09069_), .B(_09072_), .Y(_09074_));
AND_g _15313_ (.A(resetn), .B(_09073_), .Y(_09075_));
AND_g _15314_ (.A(_09066_), .B(_09075_), .Y(_09076_));
AND_g _15315_ (.A(latched_rd[3]), .B(_09076_), .Y(_09077_));
NOR_g _15316_ (.A(latched_rd[2]), .B(latched_rd[4]), .Y(_09078_));
NOR_g _15317_ (.A(latched_rd[0]), .B(latched_rd[1]), .Y(_09079_));
AND_g _15318_ (.A(_09078_), .B(_09079_), .Y(_09080_));
NAND_g _15319_ (.A(_08854_), .B(_09080_), .Y(_09081_));
AND_g _15320_ (.A(_09076_), .B(_09081_), .Y(_09082_));
NAND_g _15321_ (.A(latched_rd[0]), .B(_09076_), .Y(_09083_));
NAND_g _15322_ (.A(latched_rd[1]), .B(_09082_), .Y(_09084_));
NOR_g _15323_ (.A(_08852_), .B(_09083_), .Y(_09085_));
NOR_g _15324_ (.A(_08853_), .B(latched_rd[4]), .Y(_09086_));
AND_g _15325_ (.A(_09077_), .B(_09086_), .Y(_09087_));
AND_g _15326_ (.A(_09085_), .B(_09087_), .Y(_09088_));
NAND_g _15327_ (.A(_09085_), .B(_09087_), .Y(_09089_));
NAND_g _15328_ (.A(cpuregs[15][0]), .B(_09089_), .Y(_09090_));
NAND_g _15329_ (.A(reg_next_pc[0]), .B(latched_branch), .Y(_09091_));
NOR_g _15330_ (.A(latched_stalu), .B(reg_out[0]), .Y(_09092_));
NOR_g _15331_ (.A(_08802_), .B(alu_out_q[0]), .Y(_09093_));
AND_g _15332_ (.A(_08801_), .B(latched_store), .Y(_09094_));
NOR_g _15333_ (.A(_09092_), .B(_09093_), .Y(_09095_));
NAND_g _15334_ (.A(_09094_), .B(_09095_), .Y(_09096_));
NAND_g _15335_ (.A(_09091_), .B(_09096_), .Y(_09097_));
AND_g _15336_ (.A(_09082_), .B(_09097_), .Y(_09098_));
NAND_g _15337_ (.A(_09088_), .B(_09098_), .Y(_09099_));
AND_g _15338_ (.A(latched_rd[2]), .B(_09082_), .Y(_09100_));
NAND_g _15339_ (.A(latched_rd[2]), .B(_09082_), .Y(_09101_));
NAND_g _15340_ (.A(_09090_), .B(_09099_), .Y(_00019_));
NAND_g _15341_ (.A(cpuregs[15][1]), .B(_09089_), .Y(_09102_));
NAND_g _15342_ (.A(latched_stalu), .B(alu_out_q[1]), .Y(_09103_));
NAND_g _15343_ (.A(_08802_), .B(reg_out[1]), .Y(_09104_));
NAND_g _15344_ (.A(_09103_), .B(_09104_), .Y(_09105_));
NAND_g _15345_ (.A(_09094_), .B(_09105_), .Y(_09106_));
NAND_g _15346_ (.A(latched_branch), .B(reg_pc[1]), .Y(_09107_));
NAND_g _15347_ (.A(_09106_), .B(_09107_), .Y(_09108_));
AND_g _15348_ (.A(_09082_), .B(_09108_), .Y(_09109_));
NAND_g _15349_ (.A(_09088_), .B(_09109_), .Y(_09110_));
NAND_g _15350_ (.A(_09102_), .B(_09110_), .Y(_00020_));
NAND_g _15351_ (.A(cpuregs[15][2]), .B(_09089_), .Y(_09111_));
NAND_g _15352_ (.A(latched_stalu), .B(alu_out_q[2]), .Y(_09112_));
NAND_g _15353_ (.A(_08802_), .B(reg_out[2]), .Y(_09113_));
NAND_g _15354_ (.A(_09112_), .B(_09113_), .Y(_09114_));
NAND_g _15355_ (.A(_09094_), .B(_09114_), .Y(_09115_));
NAND_g _15356_ (.A(latched_branch), .B(_08806_), .Y(_09116_));
NAND_g _15357_ (.A(_09115_), .B(_09116_), .Y(_09117_));
AND_g _15358_ (.A(_09082_), .B(_09117_), .Y(_09118_));
NAND_g _15359_ (.A(_09088_), .B(_09118_), .Y(_09119_));
NAND_g _15360_ (.A(_09111_), .B(_09119_), .Y(_00021_));
NAND_g _15361_ (.A(cpuregs[15][3]), .B(_09089_), .Y(_09120_));
NAND_g _15362_ (.A(latched_stalu), .B(alu_out_q[3]), .Y(_09121_));
NAND_g _15363_ (.A(_08802_), .B(reg_out[3]), .Y(_09122_));
NAND_g _15364_ (.A(_09121_), .B(_09122_), .Y(_09123_));
NAND_g _15365_ (.A(_09094_), .B(_09123_), .Y(_09124_));
NOR_g _15366_ (.A(reg_pc[3]), .B(reg_pc[2]), .Y(_09125_));
AND_g _15367_ (.A(reg_pc[3]), .B(reg_pc[2]), .Y(_09126_));
NAND_g _15368_ (.A(reg_pc[3]), .B(reg_pc[2]), .Y(_09127_));
NOR_g _15369_ (.A(_08801_), .B(_09125_), .Y(_09128_));
NAND_g _15370_ (.A(_09127_), .B(_09128_), .Y(_09129_));
NAND_g _15371_ (.A(_09124_), .B(_09129_), .Y(_09130_));
AND_g _15372_ (.A(_09082_), .B(_09130_), .Y(_09131_));
NAND_g _15373_ (.A(_09088_), .B(_09131_), .Y(_09132_));
NAND_g _15374_ (.A(_09120_), .B(_09132_), .Y(_00022_));
NAND_g _15375_ (.A(cpuregs[15][4]), .B(_09089_), .Y(_09133_));
NAND_g _15376_ (.A(latched_stalu), .B(alu_out_q[4]), .Y(_09134_));
NAND_g _15377_ (.A(_08802_), .B(reg_out[4]), .Y(_09135_));
NAND_g _15378_ (.A(_09134_), .B(_09135_), .Y(_09136_));
NAND_g _15379_ (.A(_09094_), .B(_09136_), .Y(_09137_));
NOR_g _15380_ (.A(reg_pc[4]), .B(_09126_), .Y(_09138_));
AND_g _15381_ (.A(reg_pc[4]), .B(_09126_), .Y(_09139_));
NAND_g _15382_ (.A(reg_pc[4]), .B(_09126_), .Y(_09140_));
NOR_g _15383_ (.A(_08801_), .B(_09138_), .Y(_09141_));
NAND_g _15384_ (.A(_09140_), .B(_09141_), .Y(_09142_));
NAND_g _15385_ (.A(_09137_), .B(_09142_), .Y(_09143_));
AND_g _15386_ (.A(_09082_), .B(_09143_), .Y(_09144_));
NAND_g _15387_ (.A(_09088_), .B(_09144_), .Y(_09145_));
NAND_g _15388_ (.A(_09133_), .B(_09145_), .Y(_00023_));
NAND_g _15389_ (.A(cpuregs[15][5]), .B(_09089_), .Y(_09146_));
NAND_g _15390_ (.A(latched_stalu), .B(alu_out_q[5]), .Y(_09147_));
NAND_g _15391_ (.A(_08802_), .B(reg_out[5]), .Y(_09148_));
NAND_g _15392_ (.A(_09147_), .B(_09148_), .Y(_09149_));
NAND_g _15393_ (.A(_09094_), .B(_09149_), .Y(_09150_));
NOR_g _15394_ (.A(reg_pc[5]), .B(_09139_), .Y(_09151_));
AND_g _15395_ (.A(reg_pc[5]), .B(_09139_), .Y(_09152_));
NAND_g _15396_ (.A(reg_pc[5]), .B(_09139_), .Y(_09153_));
NOR_g _15397_ (.A(_08801_), .B(_09151_), .Y(_09154_));
NAND_g _15398_ (.A(_09153_), .B(_09154_), .Y(_09155_));
NAND_g _15399_ (.A(_09150_), .B(_09155_), .Y(_09156_));
AND_g _15400_ (.A(_09082_), .B(_09156_), .Y(_09157_));
NAND_g _15401_ (.A(_09088_), .B(_09157_), .Y(_09158_));
NAND_g _15402_ (.A(_09146_), .B(_09158_), .Y(_00024_));
NAND_g _15403_ (.A(cpuregs[15][6]), .B(_09089_), .Y(_09159_));
NAND_g _15404_ (.A(latched_stalu), .B(alu_out_q[6]), .Y(_09160_));
NAND_g _15405_ (.A(_08802_), .B(reg_out[6]), .Y(_09161_));
NAND_g _15406_ (.A(_09160_), .B(_09161_), .Y(_09162_));
NAND_g _15407_ (.A(_09094_), .B(_09162_), .Y(_09163_));
NOR_g _15408_ (.A(reg_pc[6]), .B(_09152_), .Y(_09164_));
AND_g _15409_ (.A(reg_pc[6]), .B(_09152_), .Y(_09165_));
NAND_g _15410_ (.A(reg_pc[6]), .B(_09152_), .Y(_09166_));
NOR_g _15411_ (.A(_08801_), .B(_09164_), .Y(_09167_));
NAND_g _15412_ (.A(_09166_), .B(_09167_), .Y(_09168_));
NAND_g _15413_ (.A(_09163_), .B(_09168_), .Y(_09169_));
AND_g _15414_ (.A(_09082_), .B(_09169_), .Y(_09170_));
NAND_g _15415_ (.A(_09088_), .B(_09170_), .Y(_09171_));
NAND_g _15416_ (.A(_09159_), .B(_09171_), .Y(_00025_));
NAND_g _15417_ (.A(cpuregs[15][7]), .B(_09089_), .Y(_09172_));
NAND_g _15418_ (.A(latched_stalu), .B(alu_out_q[7]), .Y(_09173_));
NAND_g _15419_ (.A(_08802_), .B(reg_out[7]), .Y(_09174_));
NAND_g _15420_ (.A(_09173_), .B(_09174_), .Y(_09175_));
NAND_g _15421_ (.A(_09094_), .B(_09175_), .Y(_09176_));
NOR_g _15422_ (.A(reg_pc[7]), .B(_09165_), .Y(_09177_));
AND_g _15423_ (.A(reg_pc[7]), .B(_09165_), .Y(_09178_));
NAND_g _15424_ (.A(reg_pc[7]), .B(_09165_), .Y(_09179_));
NOR_g _15425_ (.A(_08801_), .B(_09177_), .Y(_09180_));
NAND_g _15426_ (.A(_09179_), .B(_09180_), .Y(_09181_));
NAND_g _15427_ (.A(_09176_), .B(_09181_), .Y(_09182_));
AND_g _15428_ (.A(_09082_), .B(_09182_), .Y(_09183_));
NAND_g _15429_ (.A(_09088_), .B(_09183_), .Y(_09184_));
NAND_g _15430_ (.A(_09172_), .B(_09184_), .Y(_00026_));
NAND_g _15431_ (.A(cpuregs[15][8]), .B(_09089_), .Y(_09185_));
NAND_g _15432_ (.A(latched_stalu), .B(alu_out_q[8]), .Y(_09186_));
NAND_g _15433_ (.A(_08802_), .B(reg_out[8]), .Y(_09187_));
NAND_g _15434_ (.A(_09186_), .B(_09187_), .Y(_09188_));
NAND_g _15435_ (.A(_09094_), .B(_09188_), .Y(_09189_));
NOR_g _15436_ (.A(reg_pc[8]), .B(_09178_), .Y(_09190_));
AND_g _15437_ (.A(reg_pc[8]), .B(_09178_), .Y(_09191_));
NAND_g _15438_ (.A(reg_pc[8]), .B(_09178_), .Y(_09192_));
NOR_g _15439_ (.A(_08801_), .B(_09190_), .Y(_09193_));
NAND_g _15440_ (.A(_09192_), .B(_09193_), .Y(_09194_));
NAND_g _15441_ (.A(_09189_), .B(_09194_), .Y(_09195_));
AND_g _15442_ (.A(_09082_), .B(_09195_), .Y(_09196_));
NAND_g _15443_ (.A(_09088_), .B(_09196_), .Y(_09197_));
NAND_g _15444_ (.A(_09185_), .B(_09197_), .Y(_00027_));
NAND_g _15445_ (.A(cpuregs[15][9]), .B(_09089_), .Y(_09198_));
NAND_g _15446_ (.A(latched_stalu), .B(alu_out_q[9]), .Y(_09199_));
NAND_g _15447_ (.A(_08802_), .B(reg_out[9]), .Y(_09200_));
NAND_g _15448_ (.A(_09199_), .B(_09200_), .Y(_09201_));
NAND_g _15449_ (.A(_09094_), .B(_09201_), .Y(_09202_));
NOR_g _15450_ (.A(reg_pc[9]), .B(_09191_), .Y(_09203_));
AND_g _15451_ (.A(reg_pc[9]), .B(_09191_), .Y(_09204_));
NAND_g _15452_ (.A(reg_pc[9]), .B(_09191_), .Y(_09205_));
NOR_g _15453_ (.A(_08801_), .B(_09203_), .Y(_09206_));
NAND_g _15454_ (.A(_09205_), .B(_09206_), .Y(_09207_));
NAND_g _15455_ (.A(_09202_), .B(_09207_), .Y(_09208_));
AND_g _15456_ (.A(_09082_), .B(_09208_), .Y(_09209_));
NAND_g _15457_ (.A(_09088_), .B(_09209_), .Y(_09210_));
NAND_g _15458_ (.A(_09198_), .B(_09210_), .Y(_00028_));
NAND_g _15459_ (.A(cpuregs[15][10]), .B(_09089_), .Y(_09211_));
NAND_g _15460_ (.A(latched_stalu), .B(alu_out_q[10]), .Y(_09212_));
NAND_g _15461_ (.A(_08802_), .B(reg_out[10]), .Y(_09213_));
NAND_g _15462_ (.A(_09212_), .B(_09213_), .Y(_09214_));
NAND_g _15463_ (.A(_09094_), .B(_09214_), .Y(_09215_));
NOR_g _15464_ (.A(reg_pc[10]), .B(_09204_), .Y(_09216_));
AND_g _15465_ (.A(reg_pc[10]), .B(_09204_), .Y(_09217_));
NAND_g _15466_ (.A(reg_pc[10]), .B(_09204_), .Y(_09218_));
NOR_g _15467_ (.A(_08801_), .B(_09216_), .Y(_09219_));
NAND_g _15468_ (.A(_09218_), .B(_09219_), .Y(_09220_));
NAND_g _15469_ (.A(_09215_), .B(_09220_), .Y(_09221_));
AND_g _15470_ (.A(_09082_), .B(_09221_), .Y(_09222_));
NAND_g _15471_ (.A(_09088_), .B(_09222_), .Y(_09223_));
NAND_g _15472_ (.A(_09211_), .B(_09223_), .Y(_00029_));
NAND_g _15473_ (.A(cpuregs[15][11]), .B(_09089_), .Y(_09224_));
NAND_g _15474_ (.A(latched_stalu), .B(alu_out_q[11]), .Y(_09225_));
NAND_g _15475_ (.A(_08802_), .B(reg_out[11]), .Y(_09226_));
NAND_g _15476_ (.A(_09225_), .B(_09226_), .Y(_09227_));
NAND_g _15477_ (.A(_09094_), .B(_09227_), .Y(_09228_));
NOR_g _15478_ (.A(reg_pc[11]), .B(_09217_), .Y(_09229_));
AND_g _15479_ (.A(reg_pc[11]), .B(_09217_), .Y(_09230_));
NAND_g _15480_ (.A(reg_pc[11]), .B(_09217_), .Y(_09231_));
NOR_g _15481_ (.A(_08801_), .B(_09229_), .Y(_09232_));
NAND_g _15482_ (.A(_09231_), .B(_09232_), .Y(_09233_));
NAND_g _15483_ (.A(_09228_), .B(_09233_), .Y(_09234_));
AND_g _15484_ (.A(_09082_), .B(_09234_), .Y(_09235_));
NAND_g _15485_ (.A(_09088_), .B(_09235_), .Y(_09236_));
NAND_g _15486_ (.A(_09224_), .B(_09236_), .Y(_00030_));
NAND_g _15487_ (.A(cpuregs[15][12]), .B(_09089_), .Y(_09237_));
NAND_g _15488_ (.A(latched_stalu), .B(alu_out_q[12]), .Y(_09238_));
NAND_g _15489_ (.A(_08802_), .B(reg_out[12]), .Y(_09239_));
NAND_g _15490_ (.A(_09238_), .B(_09239_), .Y(_09240_));
NAND_g _15491_ (.A(_09094_), .B(_09240_), .Y(_09241_));
NOR_g _15492_ (.A(reg_pc[12]), .B(_09230_), .Y(_09242_));
AND_g _15493_ (.A(reg_pc[12]), .B(_09230_), .Y(_09243_));
NAND_g _15494_ (.A(reg_pc[12]), .B(_09230_), .Y(_09244_));
NOR_g _15495_ (.A(_08801_), .B(_09242_), .Y(_09245_));
NAND_g _15496_ (.A(_09244_), .B(_09245_), .Y(_09246_));
NAND_g _15497_ (.A(_09241_), .B(_09246_), .Y(_09247_));
AND_g _15498_ (.A(_09082_), .B(_09247_), .Y(_09248_));
NAND_g _15499_ (.A(_09088_), .B(_09248_), .Y(_09249_));
NAND_g _15500_ (.A(_09237_), .B(_09249_), .Y(_00031_));
NAND_g _15501_ (.A(cpuregs[15][13]), .B(_09089_), .Y(_09250_));
NAND_g _15502_ (.A(latched_stalu), .B(alu_out_q[13]), .Y(_09251_));
NAND_g _15503_ (.A(_08802_), .B(reg_out[13]), .Y(_09252_));
NAND_g _15504_ (.A(_09251_), .B(_09252_), .Y(_09253_));
NAND_g _15505_ (.A(_09094_), .B(_09253_), .Y(_09254_));
NOR_g _15506_ (.A(reg_pc[13]), .B(_09243_), .Y(_09255_));
AND_g _15507_ (.A(reg_pc[13]), .B(_09243_), .Y(_09256_));
NAND_g _15508_ (.A(reg_pc[13]), .B(_09243_), .Y(_09257_));
NOR_g _15509_ (.A(_08801_), .B(_09255_), .Y(_09258_));
NAND_g _15510_ (.A(_09257_), .B(_09258_), .Y(_09259_));
NAND_g _15511_ (.A(_09254_), .B(_09259_), .Y(_09260_));
AND_g _15512_ (.A(_09082_), .B(_09260_), .Y(_09261_));
NAND_g _15513_ (.A(_09088_), .B(_09261_), .Y(_09262_));
NAND_g _15514_ (.A(_09250_), .B(_09262_), .Y(_00032_));
NAND_g _15515_ (.A(cpuregs[15][14]), .B(_09089_), .Y(_09263_));
NAND_g _15516_ (.A(latched_stalu), .B(alu_out_q[14]), .Y(_09264_));
NAND_g _15517_ (.A(_08802_), .B(reg_out[14]), .Y(_09265_));
NAND_g _15518_ (.A(_09264_), .B(_09265_), .Y(_09266_));
NAND_g _15519_ (.A(_09094_), .B(_09266_), .Y(_09267_));
NOR_g _15520_ (.A(reg_pc[14]), .B(_09256_), .Y(_09268_));
AND_g _15521_ (.A(reg_pc[14]), .B(_09256_), .Y(_09269_));
NAND_g _15522_ (.A(reg_pc[14]), .B(_09256_), .Y(_09270_));
NOR_g _15523_ (.A(_08801_), .B(_09268_), .Y(_09271_));
NAND_g _15524_ (.A(_09270_), .B(_09271_), .Y(_09272_));
NAND_g _15525_ (.A(_09267_), .B(_09272_), .Y(_09273_));
AND_g _15526_ (.A(_09082_), .B(_09273_), .Y(_09274_));
NAND_g _15527_ (.A(_09088_), .B(_09274_), .Y(_09275_));
NAND_g _15528_ (.A(_09263_), .B(_09275_), .Y(_00033_));
NAND_g _15529_ (.A(cpuregs[15][15]), .B(_09089_), .Y(_09276_));
NAND_g _15530_ (.A(latched_stalu), .B(alu_out_q[15]), .Y(_09277_));
NAND_g _15531_ (.A(_08802_), .B(reg_out[15]), .Y(_09278_));
NAND_g _15532_ (.A(_09277_), .B(_09278_), .Y(_09279_));
NAND_g _15533_ (.A(_09094_), .B(_09279_), .Y(_09280_));
NOR_g _15534_ (.A(reg_pc[15]), .B(_09269_), .Y(_09281_));
AND_g _15535_ (.A(reg_pc[15]), .B(_09269_), .Y(_09282_));
NAND_g _15536_ (.A(reg_pc[15]), .B(_09269_), .Y(_09283_));
NOR_g _15537_ (.A(_08801_), .B(_09281_), .Y(_09284_));
NAND_g _15538_ (.A(_09283_), .B(_09284_), .Y(_09285_));
NAND_g _15539_ (.A(_09280_), .B(_09285_), .Y(_09286_));
AND_g _15540_ (.A(_09082_), .B(_09286_), .Y(_09287_));
NAND_g _15541_ (.A(_09088_), .B(_09287_), .Y(_09288_));
NAND_g _15542_ (.A(_09276_), .B(_09288_), .Y(_00034_));
NOR_g _15543_ (.A(cpuregs[15][16]), .B(_09088_), .Y(_09289_));
NAND_g _15544_ (.A(latched_stalu), .B(alu_out_q[16]), .Y(_09290_));
NAND_g _15545_ (.A(_08802_), .B(reg_out[16]), .Y(_09291_));
NAND_g _15546_ (.A(_09290_), .B(_09291_), .Y(_09292_));
NAND_g _15547_ (.A(_09094_), .B(_09292_), .Y(_09293_));
NOR_g _15548_ (.A(reg_pc[16]), .B(_09282_), .Y(_09294_));
AND_g _15549_ (.A(reg_pc[16]), .B(_09282_), .Y(_09295_));
NAND_g _15550_ (.A(reg_pc[16]), .B(_09282_), .Y(_09296_));
NOR_g _15551_ (.A(_08801_), .B(_09294_), .Y(_09297_));
NAND_g _15552_ (.A(_09296_), .B(_09297_), .Y(_09298_));
NAND_g _15553_ (.A(_09293_), .B(_09298_), .Y(_09299_));
AND_g _15554_ (.A(_09082_), .B(_09299_), .Y(_09300_));
NOR_g _15555_ (.A(_09089_), .B(_09300_), .Y(_09301_));
NOR_g _15556_ (.A(_09289_), .B(_09301_), .Y(_00035_));
NOR_g _15557_ (.A(cpuregs[15][17]), .B(_09088_), .Y(_09302_));
NAND_g _15558_ (.A(latched_stalu), .B(alu_out_q[17]), .Y(_09303_));
NAND_g _15559_ (.A(_08802_), .B(reg_out[17]), .Y(_09304_));
NAND_g _15560_ (.A(_09303_), .B(_09304_), .Y(_09305_));
NAND_g _15561_ (.A(_09094_), .B(_09305_), .Y(_09306_));
NOR_g _15562_ (.A(reg_pc[17]), .B(_09295_), .Y(_09307_));
AND_g _15563_ (.A(reg_pc[17]), .B(_09295_), .Y(_09308_));
NAND_g _15564_ (.A(reg_pc[17]), .B(_09295_), .Y(_09309_));
NOR_g _15565_ (.A(_08801_), .B(_09307_), .Y(_09310_));
NAND_g _15566_ (.A(_09309_), .B(_09310_), .Y(_09311_));
NAND_g _15567_ (.A(_09306_), .B(_09311_), .Y(_09312_));
AND_g _15568_ (.A(_09082_), .B(_09312_), .Y(_09313_));
NOR_g _15569_ (.A(_09089_), .B(_09313_), .Y(_09314_));
NOR_g _15570_ (.A(_09302_), .B(_09314_), .Y(_00036_));
NAND_g _15571_ (.A(latched_stalu), .B(alu_out_q[18]), .Y(_09315_));
NAND_g _15572_ (.A(_08802_), .B(reg_out[18]), .Y(_09316_));
NAND_g _15573_ (.A(_09315_), .B(_09316_), .Y(_09317_));
NAND_g _15574_ (.A(_09094_), .B(_09317_), .Y(_09318_));
NOR_g _15575_ (.A(reg_pc[18]), .B(_09308_), .Y(_09319_));
AND_g _15576_ (.A(reg_pc[18]), .B(_09308_), .Y(_09320_));
NAND_g _15577_ (.A(reg_pc[18]), .B(_09308_), .Y(_09321_));
NOR_g _15578_ (.A(_08801_), .B(_09319_), .Y(_09322_));
NAND_g _15579_ (.A(_09321_), .B(_09322_), .Y(_09323_));
NAND_g _15580_ (.A(_09318_), .B(_09323_), .Y(_09324_));
AND_g _15581_ (.A(_09082_), .B(_09324_), .Y(_09325_));
NOR_g _15582_ (.A(cpuregs[15][18]), .B(_09088_), .Y(_09326_));
NOR_g _15583_ (.A(_09089_), .B(_09325_), .Y(_09327_));
NOR_g _15584_ (.A(_09326_), .B(_09327_), .Y(_00037_));
NAND_g _15585_ (.A(latched_stalu), .B(alu_out_q[19]), .Y(_09328_));
NAND_g _15586_ (.A(_08802_), .B(reg_out[19]), .Y(_09329_));
NAND_g _15587_ (.A(_09328_), .B(_09329_), .Y(_09330_));
NAND_g _15588_ (.A(_09094_), .B(_09330_), .Y(_09331_));
NOR_g _15589_ (.A(reg_pc[19]), .B(_09320_), .Y(_09332_));
AND_g _15590_ (.A(reg_pc[19]), .B(_09320_), .Y(_09333_));
NAND_g _15591_ (.A(reg_pc[19]), .B(_09320_), .Y(_09334_));
NOR_g _15592_ (.A(_08801_), .B(_09332_), .Y(_09335_));
NAND_g _15593_ (.A(_09334_), .B(_09335_), .Y(_09336_));
NAND_g _15594_ (.A(_09331_), .B(_09336_), .Y(_09337_));
AND_g _15595_ (.A(_09082_), .B(_09337_), .Y(_09338_));
NOR_g _15596_ (.A(_09089_), .B(_09338_), .Y(_09339_));
AND_g _15597_ (.A(_08809_), .B(_09089_), .Y(_09340_));
NOR_g _15598_ (.A(_09339_), .B(_09340_), .Y(_00038_));
NAND_g _15599_ (.A(latched_stalu), .B(alu_out_q[20]), .Y(_09341_));
NAND_g _15600_ (.A(_08802_), .B(reg_out[20]), .Y(_09342_));
NAND_g _15601_ (.A(_09341_), .B(_09342_), .Y(_09343_));
NAND_g _15602_ (.A(_09094_), .B(_09343_), .Y(_09344_));
NOR_g _15603_ (.A(reg_pc[20]), .B(_09333_), .Y(_09345_));
AND_g _15604_ (.A(reg_pc[20]), .B(_09333_), .Y(_09346_));
NAND_g _15605_ (.A(reg_pc[20]), .B(_09333_), .Y(_09347_));
NOR_g _15606_ (.A(_08801_), .B(_09345_), .Y(_09348_));
NAND_g _15607_ (.A(_09347_), .B(_09348_), .Y(_09349_));
NAND_g _15608_ (.A(_09344_), .B(_09349_), .Y(_09350_));
AND_g _15609_ (.A(_09082_), .B(_09350_), .Y(_09351_));
AND_g _15610_ (.A(_08810_), .B(_09089_), .Y(_09352_));
NOR_g _15611_ (.A(_09089_), .B(_09351_), .Y(_09353_));
NOR_g _15612_ (.A(_09352_), .B(_09353_), .Y(_00039_));
NAND_g _15613_ (.A(latched_stalu), .B(alu_out_q[21]), .Y(_09354_));
NAND_g _15614_ (.A(_08802_), .B(reg_out[21]), .Y(_09355_));
NAND_g _15615_ (.A(_09354_), .B(_09355_), .Y(_09356_));
NAND_g _15616_ (.A(_09094_), .B(_09356_), .Y(_09357_));
NOR_g _15617_ (.A(reg_pc[21]), .B(_09346_), .Y(_09358_));
AND_g _15618_ (.A(reg_pc[21]), .B(_09346_), .Y(_09359_));
NAND_g _15619_ (.A(reg_pc[21]), .B(_09346_), .Y(_09360_));
NOR_g _15620_ (.A(_08801_), .B(_09358_), .Y(_09361_));
NAND_g _15621_ (.A(_09360_), .B(_09361_), .Y(_09362_));
NAND_g _15622_ (.A(_09357_), .B(_09362_), .Y(_09363_));
AND_g _15623_ (.A(_09082_), .B(_09363_), .Y(_09364_));
NOR_g _15624_ (.A(cpuregs[15][21]), .B(_09088_), .Y(_09365_));
NOR_g _15625_ (.A(_09089_), .B(_09364_), .Y(_09366_));
NOR_g _15626_ (.A(_09365_), .B(_09366_), .Y(_00040_));
NAND_g _15627_ (.A(latched_stalu), .B(alu_out_q[22]), .Y(_09367_));
NAND_g _15628_ (.A(_08802_), .B(reg_out[22]), .Y(_09368_));
NAND_g _15629_ (.A(_09367_), .B(_09368_), .Y(_09369_));
NAND_g _15630_ (.A(_09094_), .B(_09369_), .Y(_09370_));
NOR_g _15631_ (.A(reg_pc[22]), .B(_09359_), .Y(_09371_));
AND_g _15632_ (.A(reg_pc[22]), .B(_09359_), .Y(_09372_));
NAND_g _15633_ (.A(reg_pc[22]), .B(_09359_), .Y(_09373_));
NOR_g _15634_ (.A(_08801_), .B(_09371_), .Y(_09374_));
NAND_g _15635_ (.A(_09373_), .B(_09374_), .Y(_09375_));
NAND_g _15636_ (.A(_09370_), .B(_09375_), .Y(_09376_));
AND_g _15637_ (.A(_09082_), .B(_09376_), .Y(_09377_));
NOR_g _15638_ (.A(_09089_), .B(_09377_), .Y(_09378_));
NOR_g _15639_ (.A(cpuregs[15][22]), .B(_09088_), .Y(_09379_));
NOR_g _15640_ (.A(_09378_), .B(_09379_), .Y(_00041_));
NAND_g _15641_ (.A(latched_stalu), .B(alu_out_q[23]), .Y(_09380_));
NAND_g _15642_ (.A(_08802_), .B(reg_out[23]), .Y(_09381_));
NAND_g _15643_ (.A(_09380_), .B(_09381_), .Y(_09382_));
NAND_g _15644_ (.A(_09094_), .B(_09382_), .Y(_09383_));
NOR_g _15645_ (.A(reg_pc[23]), .B(_09372_), .Y(_09384_));
AND_g _15646_ (.A(reg_pc[23]), .B(_09372_), .Y(_09385_));
NAND_g _15647_ (.A(reg_pc[23]), .B(_09372_), .Y(_09386_));
NOR_g _15648_ (.A(_08801_), .B(_09384_), .Y(_09387_));
NAND_g _15649_ (.A(_09386_), .B(_09387_), .Y(_09388_));
NAND_g _15650_ (.A(_09383_), .B(_09388_), .Y(_09389_));
AND_g _15651_ (.A(_09082_), .B(_09389_), .Y(_09390_));
NOR_g _15652_ (.A(_09089_), .B(_09390_), .Y(_09391_));
NOR_g _15653_ (.A(cpuregs[15][23]), .B(_09088_), .Y(_09392_));
NOR_g _15654_ (.A(_09391_), .B(_09392_), .Y(_00042_));
NAND_g _15655_ (.A(latched_stalu), .B(alu_out_q[24]), .Y(_09393_));
NAND_g _15656_ (.A(_08802_), .B(reg_out[24]), .Y(_09394_));
NAND_g _15657_ (.A(_09393_), .B(_09394_), .Y(_09395_));
NAND_g _15658_ (.A(_09094_), .B(_09395_), .Y(_09396_));
NOR_g _15659_ (.A(reg_pc[24]), .B(_09385_), .Y(_09397_));
AND_g _15660_ (.A(reg_pc[24]), .B(_09385_), .Y(_09398_));
NAND_g _15661_ (.A(reg_pc[24]), .B(_09385_), .Y(_09399_));
NOR_g _15662_ (.A(_08801_), .B(_09397_), .Y(_09400_));
NAND_g _15663_ (.A(_09399_), .B(_09400_), .Y(_09401_));
NAND_g _15664_ (.A(_09396_), .B(_09401_), .Y(_09402_));
AND_g _15665_ (.A(_09082_), .B(_09402_), .Y(_09403_));
NOR_g _15666_ (.A(_09089_), .B(_09403_), .Y(_09404_));
NOR_g _15667_ (.A(cpuregs[15][24]), .B(_09088_), .Y(_09405_));
NOR_g _15668_ (.A(_09404_), .B(_09405_), .Y(_00043_));
NAND_g _15669_ (.A(latched_stalu), .B(alu_out_q[25]), .Y(_09406_));
NAND_g _15670_ (.A(_08802_), .B(reg_out[25]), .Y(_09407_));
NAND_g _15671_ (.A(_09406_), .B(_09407_), .Y(_09408_));
NAND_g _15672_ (.A(_09094_), .B(_09408_), .Y(_09409_));
NOR_g _15673_ (.A(reg_pc[25]), .B(_09398_), .Y(_09410_));
AND_g _15674_ (.A(reg_pc[25]), .B(_09398_), .Y(_09411_));
NAND_g _15675_ (.A(reg_pc[25]), .B(_09398_), .Y(_09412_));
NOR_g _15676_ (.A(_08801_), .B(_09410_), .Y(_09413_));
NAND_g _15677_ (.A(_09412_), .B(_09413_), .Y(_09414_));
NAND_g _15678_ (.A(_09409_), .B(_09414_), .Y(_09415_));
AND_g _15679_ (.A(_09082_), .B(_09415_), .Y(_09416_));
NOR_g _15680_ (.A(cpuregs[15][25]), .B(_09088_), .Y(_09417_));
NOR_g _15681_ (.A(_09089_), .B(_09416_), .Y(_09418_));
NOR_g _15682_ (.A(_09417_), .B(_09418_), .Y(_00044_));
NAND_g _15683_ (.A(latched_stalu), .B(alu_out_q[26]), .Y(_09419_));
NAND_g _15684_ (.A(_08802_), .B(reg_out[26]), .Y(_09420_));
NAND_g _15685_ (.A(_09419_), .B(_09420_), .Y(_09421_));
NAND_g _15686_ (.A(_09094_), .B(_09421_), .Y(_09422_));
NOR_g _15687_ (.A(reg_pc[26]), .B(_09411_), .Y(_09423_));
AND_g _15688_ (.A(reg_pc[26]), .B(_09411_), .Y(_09424_));
NAND_g _15689_ (.A(reg_pc[26]), .B(_09411_), .Y(_09425_));
NOR_g _15690_ (.A(_08801_), .B(_09423_), .Y(_09426_));
NAND_g _15691_ (.A(_09425_), .B(_09426_), .Y(_09427_));
NAND_g _15692_ (.A(_09422_), .B(_09427_), .Y(_09428_));
AND_g _15693_ (.A(_09082_), .B(_09428_), .Y(_09429_));
NOR_g _15694_ (.A(_09089_), .B(_09429_), .Y(_09430_));
NOR_g _15695_ (.A(cpuregs[15][26]), .B(_09088_), .Y(_09431_));
NOR_g _15696_ (.A(_09430_), .B(_09431_), .Y(_00045_));
NAND_g _15697_ (.A(latched_stalu), .B(alu_out_q[27]), .Y(_09432_));
NAND_g _15698_ (.A(_08802_), .B(reg_out[27]), .Y(_09433_));
NAND_g _15699_ (.A(_09432_), .B(_09433_), .Y(_09434_));
NAND_g _15700_ (.A(_09094_), .B(_09434_), .Y(_09435_));
NOR_g _15701_ (.A(reg_pc[27]), .B(_09424_), .Y(_09436_));
AND_g _15702_ (.A(reg_pc[27]), .B(_09424_), .Y(_09437_));
NAND_g _15703_ (.A(reg_pc[27]), .B(_09424_), .Y(_09438_));
NOR_g _15704_ (.A(_08801_), .B(_09436_), .Y(_09439_));
NAND_g _15705_ (.A(_09438_), .B(_09439_), .Y(_09440_));
NAND_g _15706_ (.A(_09435_), .B(_09440_), .Y(_09441_));
AND_g _15707_ (.A(_09082_), .B(_09441_), .Y(_09442_));
NOR_g _15708_ (.A(_09089_), .B(_09442_), .Y(_09443_));
NOR_g _15709_ (.A(cpuregs[15][27]), .B(_09088_), .Y(_09444_));
NOR_g _15710_ (.A(_09443_), .B(_09444_), .Y(_00046_));
NAND_g _15711_ (.A(latched_stalu), .B(alu_out_q[28]), .Y(_09445_));
NAND_g _15712_ (.A(_08802_), .B(reg_out[28]), .Y(_09446_));
NAND_g _15713_ (.A(_09445_), .B(_09446_), .Y(_09447_));
NAND_g _15714_ (.A(_09094_), .B(_09447_), .Y(_09448_));
NOR_g _15715_ (.A(reg_pc[28]), .B(_09437_), .Y(_09449_));
AND_g _15716_ (.A(reg_pc[28]), .B(_09437_), .Y(_09450_));
NAND_g _15717_ (.A(reg_pc[28]), .B(_09437_), .Y(_09451_));
NOR_g _15718_ (.A(_08801_), .B(_09449_), .Y(_09452_));
NAND_g _15719_ (.A(_09451_), .B(_09452_), .Y(_09453_));
NAND_g _15720_ (.A(_09448_), .B(_09453_), .Y(_09454_));
AND_g _15721_ (.A(_09082_), .B(_09454_), .Y(_09455_));
NOR_g _15722_ (.A(_09089_), .B(_09455_), .Y(_09456_));
NOR_g _15723_ (.A(cpuregs[15][28]), .B(_09088_), .Y(_09457_));
NOR_g _15724_ (.A(_09456_), .B(_09457_), .Y(_00047_));
NAND_g _15725_ (.A(latched_stalu), .B(alu_out_q[29]), .Y(_09458_));
NAND_g _15726_ (.A(_08802_), .B(reg_out[29]), .Y(_09459_));
NAND_g _15727_ (.A(_09458_), .B(_09459_), .Y(_09460_));
NAND_g _15728_ (.A(_09094_), .B(_09460_), .Y(_09461_));
NOR_g _15729_ (.A(reg_pc[29]), .B(_09450_), .Y(_09462_));
AND_g _15730_ (.A(reg_pc[29]), .B(_09450_), .Y(_09463_));
NAND_g _15731_ (.A(reg_pc[29]), .B(_09450_), .Y(_09464_));
NOR_g _15732_ (.A(_08801_), .B(_09462_), .Y(_09465_));
NAND_g _15733_ (.A(_09464_), .B(_09465_), .Y(_09466_));
NAND_g _15734_ (.A(_09461_), .B(_09466_), .Y(_09467_));
AND_g _15735_ (.A(_09082_), .B(_09467_), .Y(_09468_));
NOR_g _15736_ (.A(cpuregs[15][29]), .B(_09088_), .Y(_09469_));
NOR_g _15737_ (.A(_09089_), .B(_09468_), .Y(_09470_));
NOR_g _15738_ (.A(_09469_), .B(_09470_), .Y(_00048_));
NAND_g _15739_ (.A(latched_stalu), .B(alu_out_q[30]), .Y(_09471_));
NAND_g _15740_ (.A(_08802_), .B(reg_out[30]), .Y(_09472_));
NAND_g _15741_ (.A(_09471_), .B(_09472_), .Y(_09473_));
NAND_g _15742_ (.A(_09094_), .B(_09473_), .Y(_09474_));
NOR_g _15743_ (.A(reg_pc[30]), .B(_09463_), .Y(_09475_));
NAND_g _15744_ (.A(reg_pc[30]), .B(_09463_), .Y(_09476_));
NOT_g _15745_ (.A(_09476_), .Y(_09477_));
NOR_g _15746_ (.A(_08801_), .B(_09475_), .Y(_09478_));
NAND_g _15747_ (.A(_09476_), .B(_09478_), .Y(_09479_));
NAND_g _15748_ (.A(_09474_), .B(_09479_), .Y(_09480_));
AND_g _15749_ (.A(_09082_), .B(_09480_), .Y(_09481_));
NOR_g _15750_ (.A(_09089_), .B(_09481_), .Y(_09482_));
NOR_g _15751_ (.A(cpuregs[15][30]), .B(_09088_), .Y(_09483_));
NOR_g _15752_ (.A(_09482_), .B(_09483_), .Y(_00049_));
NAND_g _15753_ (.A(latched_stalu), .B(alu_out_q[31]), .Y(_09484_));
NAND_g _15754_ (.A(_08802_), .B(reg_out[31]), .Y(_09485_));
NAND_g _15755_ (.A(_09484_), .B(_09485_), .Y(_09486_));
NAND_g _15756_ (.A(_09094_), .B(_09486_), .Y(_09487_));
NAND_g _15757_ (.A(reg_pc[31]), .B(_09477_), .Y(_09488_));
NAND_g _15758_ (.A(_08805_), .B(_09476_), .Y(_09489_));
AND_g _15759_ (.A(latched_branch), .B(_09489_), .Y(_09490_));
NAND_g _15760_ (.A(_09488_), .B(_09490_), .Y(_09491_));
NAND_g _15761_ (.A(_09487_), .B(_09491_), .Y(_09492_));
AND_g _15762_ (.A(_09082_), .B(_09492_), .Y(_09493_));
NOR_g _15763_ (.A(_09089_), .B(_09493_), .Y(_09494_));
NOR_g _15764_ (.A(cpuregs[15][31]), .B(_09088_), .Y(_09495_));
NOR_g _15765_ (.A(_09494_), .B(_09495_), .Y(_00050_));
NOR_g _15766_ (.A(latched_rd[0]), .B(_09084_), .Y(_09496_));
AND_g _15767_ (.A(latched_rd[4]), .B(_09082_), .Y(_09497_));
NAND_g _15768_ (.A(latched_rd[4]), .B(_09077_), .Y(_09498_));
NOR_g _15769_ (.A(_08853_), .B(_09498_), .Y(_09499_));
AND_g _15770_ (.A(_09496_), .B(_09499_), .Y(_09500_));
NAND_g _15771_ (.A(_09496_), .B(_09499_), .Y(_09501_));
NAND_g _15772_ (.A(_09098_), .B(_09500_), .Y(_09502_));
NAND_g _15773_ (.A(cpuregs[30][0]), .B(_09501_), .Y(_09503_));
NAND_g _15774_ (.A(_09502_), .B(_09503_), .Y(_00051_));
NAND_g _15775_ (.A(_09109_), .B(_09500_), .Y(_09504_));
NAND_g _15776_ (.A(cpuregs[30][1]), .B(_09501_), .Y(_09505_));
NAND_g _15777_ (.A(_09504_), .B(_09505_), .Y(_00052_));
NAND_g _15778_ (.A(_09118_), .B(_09500_), .Y(_09506_));
NAND_g _15779_ (.A(cpuregs[30][2]), .B(_09501_), .Y(_09507_));
NAND_g _15780_ (.A(_09506_), .B(_09507_), .Y(_00053_));
NAND_g _15781_ (.A(_09131_), .B(_09500_), .Y(_09508_));
NAND_g _15782_ (.A(cpuregs[30][3]), .B(_09501_), .Y(_09509_));
NAND_g _15783_ (.A(_09508_), .B(_09509_), .Y(_00054_));
NAND_g _15784_ (.A(_09144_), .B(_09500_), .Y(_09510_));
NAND_g _15785_ (.A(cpuregs[30][4]), .B(_09501_), .Y(_09511_));
NAND_g _15786_ (.A(_09510_), .B(_09511_), .Y(_00055_));
NAND_g _15787_ (.A(_09157_), .B(_09500_), .Y(_09512_));
NAND_g _15788_ (.A(cpuregs[30][5]), .B(_09501_), .Y(_09513_));
NAND_g _15789_ (.A(_09512_), .B(_09513_), .Y(_00056_));
NAND_g _15790_ (.A(_09170_), .B(_09500_), .Y(_09514_));
NAND_g _15791_ (.A(cpuregs[30][6]), .B(_09501_), .Y(_09515_));
NAND_g _15792_ (.A(_09514_), .B(_09515_), .Y(_00057_));
NAND_g _15793_ (.A(_09183_), .B(_09500_), .Y(_09516_));
NAND_g _15794_ (.A(cpuregs[30][7]), .B(_09501_), .Y(_09517_));
NAND_g _15795_ (.A(_09516_), .B(_09517_), .Y(_00058_));
NAND_g _15796_ (.A(_09196_), .B(_09500_), .Y(_09518_));
NAND_g _15797_ (.A(cpuregs[30][8]), .B(_09501_), .Y(_09519_));
NAND_g _15798_ (.A(_09518_), .B(_09519_), .Y(_00059_));
NAND_g _15799_ (.A(_09209_), .B(_09500_), .Y(_09520_));
NAND_g _15800_ (.A(cpuregs[30][9]), .B(_09501_), .Y(_09521_));
NAND_g _15801_ (.A(_09520_), .B(_09521_), .Y(_00060_));
NAND_g _15802_ (.A(_09222_), .B(_09500_), .Y(_09522_));
NAND_g _15803_ (.A(cpuregs[30][10]), .B(_09501_), .Y(_09523_));
NAND_g _15804_ (.A(_09522_), .B(_09523_), .Y(_00061_));
NAND_g _15805_ (.A(_09235_), .B(_09500_), .Y(_09524_));
NAND_g _15806_ (.A(cpuregs[30][11]), .B(_09501_), .Y(_09525_));
NAND_g _15807_ (.A(_09524_), .B(_09525_), .Y(_00062_));
NAND_g _15808_ (.A(_09248_), .B(_09500_), .Y(_09526_));
NAND_g _15809_ (.A(cpuregs[30][12]), .B(_09501_), .Y(_09527_));
NAND_g _15810_ (.A(_09526_), .B(_09527_), .Y(_00063_));
NAND_g _15811_ (.A(_09261_), .B(_09500_), .Y(_09528_));
NAND_g _15812_ (.A(cpuregs[30][13]), .B(_09501_), .Y(_09529_));
NAND_g _15813_ (.A(_09528_), .B(_09529_), .Y(_00064_));
NAND_g _15814_ (.A(_09274_), .B(_09500_), .Y(_09530_));
NAND_g _15815_ (.A(cpuregs[30][14]), .B(_09501_), .Y(_09531_));
NAND_g _15816_ (.A(_09530_), .B(_09531_), .Y(_00065_));
NAND_g _15817_ (.A(_09287_), .B(_09500_), .Y(_09532_));
NAND_g _15818_ (.A(cpuregs[30][15]), .B(_09501_), .Y(_09533_));
NAND_g _15819_ (.A(_09532_), .B(_09533_), .Y(_00066_));
NAND_g _15820_ (.A(_09300_), .B(_09500_), .Y(_09534_));
NAND_g _15821_ (.A(cpuregs[30][16]), .B(_09501_), .Y(_09535_));
NAND_g _15822_ (.A(_09534_), .B(_09535_), .Y(_00067_));
NOR_g _15823_ (.A(cpuregs[30][17]), .B(_09500_), .Y(_09536_));
NOR_g _15824_ (.A(_09313_), .B(_09501_), .Y(_09537_));
NOR_g _15825_ (.A(_09536_), .B(_09537_), .Y(_00068_));
NAND_g _15826_ (.A(_09325_), .B(_09500_), .Y(_09538_));
NAND_g _15827_ (.A(cpuregs[30][18]), .B(_09501_), .Y(_09539_));
NAND_g _15828_ (.A(_09538_), .B(_09539_), .Y(_00069_));
NAND_g _15829_ (.A(_09338_), .B(_09500_), .Y(_09540_));
NAND_g _15830_ (.A(cpuregs[30][19]), .B(_09501_), .Y(_09541_));
NAND_g _15831_ (.A(_09540_), .B(_09541_), .Y(_00070_));
NAND_g _15832_ (.A(_09351_), .B(_09500_), .Y(_09542_));
NAND_g _15833_ (.A(cpuregs[30][20]), .B(_09501_), .Y(_09543_));
NAND_g _15834_ (.A(_09542_), .B(_09543_), .Y(_00071_));
NAND_g _15835_ (.A(_09364_), .B(_09500_), .Y(_09544_));
NAND_g _15836_ (.A(cpuregs[30][21]), .B(_09501_), .Y(_09545_));
NAND_g _15837_ (.A(_09544_), .B(_09545_), .Y(_00072_));
NAND_g _15838_ (.A(_09377_), .B(_09500_), .Y(_09546_));
NAND_g _15839_ (.A(cpuregs[30][22]), .B(_09501_), .Y(_09547_));
NAND_g _15840_ (.A(_09546_), .B(_09547_), .Y(_00073_));
NAND_g _15841_ (.A(_09390_), .B(_09500_), .Y(_09548_));
NAND_g _15842_ (.A(cpuregs[30][23]), .B(_09501_), .Y(_09549_));
NAND_g _15843_ (.A(_09548_), .B(_09549_), .Y(_00074_));
NAND_g _15844_ (.A(_09403_), .B(_09500_), .Y(_09550_));
NAND_g _15845_ (.A(cpuregs[30][24]), .B(_09501_), .Y(_09551_));
NAND_g _15846_ (.A(_09550_), .B(_09551_), .Y(_00075_));
NAND_g _15847_ (.A(_09416_), .B(_09500_), .Y(_09552_));
NAND_g _15848_ (.A(cpuregs[30][25]), .B(_09501_), .Y(_09553_));
NAND_g _15849_ (.A(_09552_), .B(_09553_), .Y(_00076_));
NAND_g _15850_ (.A(_09429_), .B(_09500_), .Y(_09554_));
NAND_g _15851_ (.A(cpuregs[30][26]), .B(_09501_), .Y(_09555_));
NAND_g _15852_ (.A(_09554_), .B(_09555_), .Y(_00077_));
NAND_g _15853_ (.A(_09442_), .B(_09500_), .Y(_09556_));
NAND_g _15854_ (.A(cpuregs[30][27]), .B(_09501_), .Y(_09557_));
NAND_g _15855_ (.A(_09556_), .B(_09557_), .Y(_00078_));
NAND_g _15856_ (.A(_09455_), .B(_09500_), .Y(_09558_));
NAND_g _15857_ (.A(cpuregs[30][28]), .B(_09501_), .Y(_09559_));
NAND_g _15858_ (.A(_09558_), .B(_09559_), .Y(_00079_));
NAND_g _15859_ (.A(_09468_), .B(_09500_), .Y(_09560_));
NAND_g _15860_ (.A(cpuregs[30][29]), .B(_09501_), .Y(_09561_));
NAND_g _15861_ (.A(_09560_), .B(_09561_), .Y(_00080_));
NAND_g _15862_ (.A(_09481_), .B(_09500_), .Y(_09562_));
NAND_g _15863_ (.A(cpuregs[30][30]), .B(_09501_), .Y(_09563_));
NAND_g _15864_ (.A(_09562_), .B(_09563_), .Y(_00081_));
NAND_g _15865_ (.A(_09493_), .B(_09500_), .Y(_09564_));
NAND_g _15866_ (.A(cpuregs[30][31]), .B(_09501_), .Y(_09565_));
NAND_g _15867_ (.A(_09564_), .B(_09565_), .Y(_00082_));
NOR_g _15868_ (.A(_09077_), .B(_09497_), .Y(_09566_));
AND_g _15869_ (.A(_09101_), .B(_09566_), .Y(_09567_));
AND_g _15870_ (.A(_09496_), .B(_09567_), .Y(_09568_));
NAND_g _15871_ (.A(_09496_), .B(_09567_), .Y(_09569_));
NAND_g _15872_ (.A(_09098_), .B(_09568_), .Y(_09570_));
NAND_g _15873_ (.A(cpuregs[2][0]), .B(_09569_), .Y(_09571_));
NAND_g _15874_ (.A(_09570_), .B(_09571_), .Y(_00083_));
NAND_g _15875_ (.A(_09109_), .B(_09568_), .Y(_09572_));
NAND_g _15876_ (.A(cpuregs[2][1]), .B(_09569_), .Y(_09573_));
NAND_g _15877_ (.A(_09572_), .B(_09573_), .Y(_00084_));
NAND_g _15878_ (.A(_09118_), .B(_09568_), .Y(_09574_));
NAND_g _15879_ (.A(cpuregs[2][2]), .B(_09569_), .Y(_09575_));
NAND_g _15880_ (.A(_09574_), .B(_09575_), .Y(_00085_));
NAND_g _15881_ (.A(_09131_), .B(_09568_), .Y(_09576_));
NAND_g _15882_ (.A(cpuregs[2][3]), .B(_09569_), .Y(_09577_));
NAND_g _15883_ (.A(_09576_), .B(_09577_), .Y(_00086_));
NAND_g _15884_ (.A(_09144_), .B(_09568_), .Y(_09578_));
NAND_g _15885_ (.A(cpuregs[2][4]), .B(_09569_), .Y(_09579_));
NAND_g _15886_ (.A(_09578_), .B(_09579_), .Y(_00087_));
NAND_g _15887_ (.A(_09157_), .B(_09568_), .Y(_09580_));
NAND_g _15888_ (.A(cpuregs[2][5]), .B(_09569_), .Y(_09581_));
NAND_g _15889_ (.A(_09580_), .B(_09581_), .Y(_00088_));
NAND_g _15890_ (.A(_09170_), .B(_09568_), .Y(_09582_));
NAND_g _15891_ (.A(cpuregs[2][6]), .B(_09569_), .Y(_09583_));
NAND_g _15892_ (.A(_09582_), .B(_09583_), .Y(_00089_));
NAND_g _15893_ (.A(_09183_), .B(_09568_), .Y(_09584_));
NAND_g _15894_ (.A(cpuregs[2][7]), .B(_09569_), .Y(_09585_));
NAND_g _15895_ (.A(_09584_), .B(_09585_), .Y(_00090_));
NAND_g _15896_ (.A(_09196_), .B(_09568_), .Y(_09586_));
NAND_g _15897_ (.A(cpuregs[2][8]), .B(_09569_), .Y(_09587_));
NAND_g _15898_ (.A(_09586_), .B(_09587_), .Y(_00091_));
NAND_g _15899_ (.A(_09209_), .B(_09568_), .Y(_09588_));
NAND_g _15900_ (.A(cpuregs[2][9]), .B(_09569_), .Y(_09589_));
NAND_g _15901_ (.A(_09588_), .B(_09589_), .Y(_00092_));
NAND_g _15902_ (.A(_09222_), .B(_09568_), .Y(_09590_));
NAND_g _15903_ (.A(cpuregs[2][10]), .B(_09569_), .Y(_09591_));
NAND_g _15904_ (.A(_09590_), .B(_09591_), .Y(_00093_));
NAND_g _15905_ (.A(_09235_), .B(_09568_), .Y(_09592_));
NAND_g _15906_ (.A(cpuregs[2][11]), .B(_09569_), .Y(_09593_));
NAND_g _15907_ (.A(_09592_), .B(_09593_), .Y(_00094_));
NAND_g _15908_ (.A(_09248_), .B(_09568_), .Y(_09594_));
NAND_g _15909_ (.A(cpuregs[2][12]), .B(_09569_), .Y(_09595_));
NAND_g _15910_ (.A(_09594_), .B(_09595_), .Y(_00095_));
NAND_g _15911_ (.A(_09261_), .B(_09568_), .Y(_09596_));
NAND_g _15912_ (.A(cpuregs[2][13]), .B(_09569_), .Y(_09597_));
NAND_g _15913_ (.A(_09596_), .B(_09597_), .Y(_00096_));
NAND_g _15914_ (.A(_09274_), .B(_09568_), .Y(_09598_));
NAND_g _15915_ (.A(cpuregs[2][14]), .B(_09569_), .Y(_09599_));
NAND_g _15916_ (.A(_09598_), .B(_09599_), .Y(_00097_));
NAND_g _15917_ (.A(_09287_), .B(_09568_), .Y(_09600_));
NAND_g _15918_ (.A(cpuregs[2][15]), .B(_09569_), .Y(_09601_));
NAND_g _15919_ (.A(_09600_), .B(_09601_), .Y(_00098_));
NAND_g _15920_ (.A(_09300_), .B(_09568_), .Y(_09602_));
NAND_g _15921_ (.A(cpuregs[2][16]), .B(_09569_), .Y(_09603_));
NAND_g _15922_ (.A(_09602_), .B(_09603_), .Y(_00099_));
NOR_g _15923_ (.A(cpuregs[2][17]), .B(_09568_), .Y(_09604_));
NOR_g _15924_ (.A(_09313_), .B(_09569_), .Y(_09605_));
NOR_g _15925_ (.A(_09604_), .B(_09605_), .Y(_00100_));
NOR_g _15926_ (.A(cpuregs[2][18]), .B(_09568_), .Y(_09606_));
NOR_g _15927_ (.A(_09325_), .B(_09569_), .Y(_09607_));
NOR_g _15928_ (.A(_09606_), .B(_09607_), .Y(_00101_));
NAND_g _15929_ (.A(_09338_), .B(_09568_), .Y(_09608_));
NAND_g _15930_ (.A(cpuregs[2][19]), .B(_09569_), .Y(_09609_));
NAND_g _15931_ (.A(_09608_), .B(_09609_), .Y(_00102_));
NAND_g _15932_ (.A(_09351_), .B(_09568_), .Y(_09610_));
NAND_g _15933_ (.A(cpuregs[2][20]), .B(_09569_), .Y(_09611_));
NAND_g _15934_ (.A(_09610_), .B(_09611_), .Y(_00103_));
NAND_g _15935_ (.A(_09364_), .B(_09568_), .Y(_09612_));
NAND_g _15936_ (.A(cpuregs[2][21]), .B(_09569_), .Y(_09613_));
NAND_g _15937_ (.A(_09612_), .B(_09613_), .Y(_00104_));
NAND_g _15938_ (.A(_09377_), .B(_09568_), .Y(_09614_));
NAND_g _15939_ (.A(cpuregs[2][22]), .B(_09569_), .Y(_09615_));
NAND_g _15940_ (.A(_09614_), .B(_09615_), .Y(_00105_));
NAND_g _15941_ (.A(_09390_), .B(_09568_), .Y(_09616_));
NAND_g _15942_ (.A(cpuregs[2][23]), .B(_09569_), .Y(_09617_));
NAND_g _15943_ (.A(_09616_), .B(_09617_), .Y(_00106_));
NAND_g _15944_ (.A(_09403_), .B(_09568_), .Y(_09618_));
NAND_g _15945_ (.A(cpuregs[2][24]), .B(_09569_), .Y(_09619_));
NAND_g _15946_ (.A(_09618_), .B(_09619_), .Y(_00107_));
NAND_g _15947_ (.A(_09416_), .B(_09568_), .Y(_09620_));
NAND_g _15948_ (.A(cpuregs[2][25]), .B(_09569_), .Y(_09621_));
NAND_g _15949_ (.A(_09620_), .B(_09621_), .Y(_00108_));
NAND_g _15950_ (.A(_09429_), .B(_09568_), .Y(_09622_));
NAND_g _15951_ (.A(cpuregs[2][26]), .B(_09569_), .Y(_09623_));
NAND_g _15952_ (.A(_09622_), .B(_09623_), .Y(_00109_));
NAND_g _15953_ (.A(_09442_), .B(_09568_), .Y(_09624_));
NAND_g _15954_ (.A(cpuregs[2][27]), .B(_09569_), .Y(_09625_));
NAND_g _15955_ (.A(_09624_), .B(_09625_), .Y(_00110_));
NAND_g _15956_ (.A(_09455_), .B(_09568_), .Y(_09626_));
NAND_g _15957_ (.A(cpuregs[2][28]), .B(_09569_), .Y(_09627_));
NAND_g _15958_ (.A(_09626_), .B(_09627_), .Y(_00111_));
NAND_g _15959_ (.A(_09468_), .B(_09568_), .Y(_09628_));
NAND_g _15960_ (.A(cpuregs[2][29]), .B(_09569_), .Y(_09629_));
NAND_g _15961_ (.A(_09628_), .B(_09629_), .Y(_00112_));
NAND_g _15962_ (.A(_09481_), .B(_09568_), .Y(_09630_));
NAND_g _15963_ (.A(cpuregs[2][30]), .B(_09569_), .Y(_09631_));
NAND_g _15964_ (.A(_09630_), .B(_09631_), .Y(_00113_));
NAND_g _15965_ (.A(_09493_), .B(_09568_), .Y(_09632_));
NAND_g _15966_ (.A(cpuregs[2][31]), .B(_09569_), .Y(_09633_));
NAND_g _15967_ (.A(_09632_), .B(_09633_), .Y(_00114_));
NOR_g _15968_ (.A(_08811_), .B(count_cycle[0]), .Y(_00115_));
NAND_g _15969_ (.A(count_cycle[0]), .B(count_cycle[1]), .Y(_09634_));
NOR_g _15970_ (.A(count_cycle[0]), .B(count_cycle[1]), .Y(_09635_));
NOR_g _15971_ (.A(_08811_), .B(_09635_), .Y(_09636_));
AND_g _15972_ (.A(_09634_), .B(_09636_), .Y(_00116_));
NOR_g _15973_ (.A(_09034_), .B(_09634_), .Y(_09637_));
NAND_g _15974_ (.A(_09034_), .B(_09634_), .Y(_09638_));
NAND_g _15975_ (.A(resetn), .B(_09638_), .Y(_09639_));
NOR_g _15976_ (.A(_09637_), .B(_09639_), .Y(_00117_));
NAND_g _15977_ (.A(count_cycle[3]), .B(_09637_), .Y(_09640_));
NOR_g _15978_ (.A(count_cycle[3]), .B(_09637_), .Y(_09641_));
NOR_g _15979_ (.A(_08811_), .B(_09641_), .Y(_09642_));
AND_g _15980_ (.A(_09640_), .B(_09642_), .Y(_00118_));
NOR_g _15981_ (.A(_09035_), .B(_09640_), .Y(_09643_));
NAND_g _15982_ (.A(_09035_), .B(_09640_), .Y(_09644_));
NAND_g _15983_ (.A(resetn), .B(_09644_), .Y(_09645_));
NOR_g _15984_ (.A(_09643_), .B(_09645_), .Y(_00119_));
NAND_g _15985_ (.A(count_cycle[5]), .B(_09643_), .Y(_09646_));
NOR_g _15986_ (.A(count_cycle[5]), .B(_09643_), .Y(_09647_));
NOR_g _15987_ (.A(_08811_), .B(_09647_), .Y(_09648_));
AND_g _15988_ (.A(_09646_), .B(_09648_), .Y(_00120_));
NOR_g _15989_ (.A(_09036_), .B(_09646_), .Y(_09649_));
NAND_g _15990_ (.A(_09036_), .B(_09646_), .Y(_09650_));
NAND_g _15991_ (.A(resetn), .B(_09650_), .Y(_09651_));
NOR_g _15992_ (.A(_09649_), .B(_09651_), .Y(_00121_));
NAND_g _15993_ (.A(count_cycle[7]), .B(_09649_), .Y(_09652_));
NOR_g _15994_ (.A(count_cycle[7]), .B(_09649_), .Y(_09653_));
NOR_g _15995_ (.A(_08811_), .B(_09653_), .Y(_09654_));
AND_g _15996_ (.A(_09652_), .B(_09654_), .Y(_00122_));
NOR_g _15997_ (.A(_09037_), .B(_09652_), .Y(_09655_));
NAND_g _15998_ (.A(_09037_), .B(_09652_), .Y(_09656_));
NAND_g _15999_ (.A(resetn), .B(_09656_), .Y(_09657_));
NOR_g _16000_ (.A(_09655_), .B(_09657_), .Y(_00123_));
NAND_g _16001_ (.A(count_cycle[9]), .B(_09655_), .Y(_09658_));
NOR_g _16002_ (.A(count_cycle[9]), .B(_09655_), .Y(_09659_));
NOR_g _16003_ (.A(_08811_), .B(_09659_), .Y(_09660_));
AND_g _16004_ (.A(_09658_), .B(_09660_), .Y(_00124_));
NOR_g _16005_ (.A(_09038_), .B(_09658_), .Y(_09661_));
NAND_g _16006_ (.A(_09038_), .B(_09658_), .Y(_09662_));
NAND_g _16007_ (.A(resetn), .B(_09662_), .Y(_09663_));
NOR_g _16008_ (.A(_09661_), .B(_09663_), .Y(_00125_));
NAND_g _16009_ (.A(count_cycle[11]), .B(_09661_), .Y(_09664_));
NOR_g _16010_ (.A(count_cycle[11]), .B(_09661_), .Y(_09665_));
NOR_g _16011_ (.A(_08811_), .B(_09665_), .Y(_09666_));
AND_g _16012_ (.A(_09664_), .B(_09666_), .Y(_00126_));
NOR_g _16013_ (.A(_09039_), .B(_09664_), .Y(_09667_));
NAND_g _16014_ (.A(_09039_), .B(_09664_), .Y(_09668_));
NAND_g _16015_ (.A(resetn), .B(_09668_), .Y(_09669_));
NOR_g _16016_ (.A(_09667_), .B(_09669_), .Y(_00127_));
NAND_g _16017_ (.A(count_cycle[13]), .B(_09667_), .Y(_09670_));
NOR_g _16018_ (.A(count_cycle[13]), .B(_09667_), .Y(_09671_));
NOR_g _16019_ (.A(_08811_), .B(_09671_), .Y(_09672_));
AND_g _16020_ (.A(_09670_), .B(_09672_), .Y(_00128_));
NOR_g _16021_ (.A(_09040_), .B(_09670_), .Y(_09673_));
NAND_g _16022_ (.A(_09040_), .B(_09670_), .Y(_09674_));
NAND_g _16023_ (.A(resetn), .B(_09674_), .Y(_09675_));
NOR_g _16024_ (.A(_09673_), .B(_09675_), .Y(_00129_));
NAND_g _16025_ (.A(count_cycle[15]), .B(_09673_), .Y(_09676_));
NOR_g _16026_ (.A(count_cycle[15]), .B(_09673_), .Y(_09677_));
NOR_g _16027_ (.A(_08811_), .B(_09677_), .Y(_09678_));
AND_g _16028_ (.A(_09676_), .B(_09678_), .Y(_00130_));
NOR_g _16029_ (.A(_09041_), .B(_09676_), .Y(_09679_));
NAND_g _16030_ (.A(_09041_), .B(_09676_), .Y(_09680_));
NAND_g _16031_ (.A(resetn), .B(_09680_), .Y(_09681_));
NOR_g _16032_ (.A(_09679_), .B(_09681_), .Y(_00131_));
NAND_g _16033_ (.A(count_cycle[17]), .B(_09679_), .Y(_09682_));
NOR_g _16034_ (.A(count_cycle[17]), .B(_09679_), .Y(_09683_));
NOR_g _16035_ (.A(_08811_), .B(_09683_), .Y(_09684_));
AND_g _16036_ (.A(_09682_), .B(_09684_), .Y(_00132_));
NOR_g _16037_ (.A(_09042_), .B(_09682_), .Y(_09685_));
NAND_g _16038_ (.A(_09042_), .B(_09682_), .Y(_09686_));
NAND_g _16039_ (.A(resetn), .B(_09686_), .Y(_09687_));
NOR_g _16040_ (.A(_09685_), .B(_09687_), .Y(_00133_));
NAND_g _16041_ (.A(count_cycle[19]), .B(_09685_), .Y(_09688_));
NOR_g _16042_ (.A(count_cycle[19]), .B(_09685_), .Y(_09689_));
NOR_g _16043_ (.A(_08811_), .B(_09689_), .Y(_09690_));
AND_g _16044_ (.A(_09688_), .B(_09690_), .Y(_00134_));
NOR_g _16045_ (.A(_09043_), .B(_09688_), .Y(_09691_));
NAND_g _16046_ (.A(_09043_), .B(_09688_), .Y(_09692_));
NAND_g _16047_ (.A(resetn), .B(_09692_), .Y(_09693_));
NOR_g _16048_ (.A(_09691_), .B(_09693_), .Y(_00135_));
NAND_g _16049_ (.A(count_cycle[21]), .B(_09691_), .Y(_09694_));
NOR_g _16050_ (.A(count_cycle[21]), .B(_09691_), .Y(_09695_));
NOR_g _16051_ (.A(_08811_), .B(_09695_), .Y(_09696_));
AND_g _16052_ (.A(_09694_), .B(_09696_), .Y(_00136_));
NOR_g _16053_ (.A(_09044_), .B(_09694_), .Y(_09697_));
NAND_g _16054_ (.A(_09044_), .B(_09694_), .Y(_09698_));
NAND_g _16055_ (.A(resetn), .B(_09698_), .Y(_09699_));
NOR_g _16056_ (.A(_09697_), .B(_09699_), .Y(_00137_));
NAND_g _16057_ (.A(count_cycle[23]), .B(_09697_), .Y(_09700_));
NOR_g _16058_ (.A(count_cycle[23]), .B(_09697_), .Y(_09701_));
NOR_g _16059_ (.A(_08811_), .B(_09701_), .Y(_09702_));
AND_g _16060_ (.A(_09700_), .B(_09702_), .Y(_00138_));
NOR_g _16061_ (.A(_09045_), .B(_09700_), .Y(_09703_));
NAND_g _16062_ (.A(_09045_), .B(_09700_), .Y(_09704_));
NAND_g _16063_ (.A(resetn), .B(_09704_), .Y(_09705_));
NOR_g _16064_ (.A(_09703_), .B(_09705_), .Y(_00139_));
NAND_g _16065_ (.A(count_cycle[25]), .B(_09703_), .Y(_09706_));
NOR_g _16066_ (.A(count_cycle[25]), .B(_09703_), .Y(_09707_));
NOR_g _16067_ (.A(_08811_), .B(_09707_), .Y(_09708_));
AND_g _16068_ (.A(_09706_), .B(_09708_), .Y(_00140_));
NOR_g _16069_ (.A(_09046_), .B(_09706_), .Y(_09709_));
NAND_g _16070_ (.A(_09046_), .B(_09706_), .Y(_09710_));
NAND_g _16071_ (.A(resetn), .B(_09710_), .Y(_09711_));
NOR_g _16072_ (.A(_09709_), .B(_09711_), .Y(_00141_));
NAND_g _16073_ (.A(count_cycle[27]), .B(_09709_), .Y(_09712_));
NOR_g _16074_ (.A(count_cycle[27]), .B(_09709_), .Y(_09713_));
NOR_g _16075_ (.A(_08811_), .B(_09713_), .Y(_09714_));
AND_g _16076_ (.A(_09712_), .B(_09714_), .Y(_00142_));
NOR_g _16077_ (.A(_09047_), .B(_09712_), .Y(_09715_));
NAND_g _16078_ (.A(_09047_), .B(_09712_), .Y(_09716_));
NAND_g _16079_ (.A(resetn), .B(_09716_), .Y(_09717_));
NOR_g _16080_ (.A(_09715_), .B(_09717_), .Y(_00143_));
NAND_g _16081_ (.A(count_cycle[29]), .B(_09715_), .Y(_09718_));
NOR_g _16082_ (.A(count_cycle[29]), .B(_09715_), .Y(_09719_));
NOR_g _16083_ (.A(_08811_), .B(_09719_), .Y(_09720_));
AND_g _16084_ (.A(_09718_), .B(_09720_), .Y(_00144_));
NOR_g _16085_ (.A(_09048_), .B(_09718_), .Y(_09721_));
NAND_g _16086_ (.A(_09048_), .B(_09718_), .Y(_09722_));
NAND_g _16087_ (.A(resetn), .B(_09722_), .Y(_09723_));
NOR_g _16088_ (.A(_09721_), .B(_09723_), .Y(_00145_));
NAND_g _16089_ (.A(count_cycle[31]), .B(_09721_), .Y(_09724_));
NOR_g _16090_ (.A(count_cycle[31]), .B(_09721_), .Y(_09725_));
NOR_g _16091_ (.A(_08811_), .B(_09725_), .Y(_09726_));
AND_g _16092_ (.A(_09724_), .B(_09726_), .Y(_00146_));
NOR_g _16093_ (.A(_09049_), .B(_09724_), .Y(_09727_));
NAND_g _16094_ (.A(_09049_), .B(_09724_), .Y(_09728_));
NAND_g _16095_ (.A(resetn), .B(_09728_), .Y(_09729_));
NOR_g _16096_ (.A(_09727_), .B(_09729_), .Y(_00147_));
NAND_g _16097_ (.A(count_cycle[33]), .B(_09727_), .Y(_09730_));
NOR_g _16098_ (.A(count_cycle[33]), .B(_09727_), .Y(_09731_));
NOR_g _16099_ (.A(_08811_), .B(_09731_), .Y(_09732_));
AND_g _16100_ (.A(_09730_), .B(_09732_), .Y(_00148_));
NOR_g _16101_ (.A(_09050_), .B(_09730_), .Y(_09733_));
NAND_g _16102_ (.A(_09050_), .B(_09730_), .Y(_09734_));
NAND_g _16103_ (.A(resetn), .B(_09734_), .Y(_09735_));
NOR_g _16104_ (.A(_09733_), .B(_09735_), .Y(_00149_));
NAND_g _16105_ (.A(count_cycle[35]), .B(_09733_), .Y(_09736_));
NOR_g _16106_ (.A(count_cycle[35]), .B(_09733_), .Y(_09737_));
NOR_g _16107_ (.A(_08811_), .B(_09737_), .Y(_09738_));
AND_g _16108_ (.A(_09736_), .B(_09738_), .Y(_00150_));
NOR_g _16109_ (.A(_09051_), .B(_09736_), .Y(_09739_));
NAND_g _16110_ (.A(_09051_), .B(_09736_), .Y(_09740_));
NAND_g _16111_ (.A(resetn), .B(_09740_), .Y(_09741_));
NOR_g _16112_ (.A(_09739_), .B(_09741_), .Y(_00151_));
NAND_g _16113_ (.A(count_cycle[37]), .B(_09739_), .Y(_09742_));
NOR_g _16114_ (.A(count_cycle[37]), .B(_09739_), .Y(_09743_));
NOR_g _16115_ (.A(_08811_), .B(_09743_), .Y(_09744_));
AND_g _16116_ (.A(_09742_), .B(_09744_), .Y(_00152_));
NOR_g _16117_ (.A(_09052_), .B(_09742_), .Y(_09745_));
NAND_g _16118_ (.A(_09052_), .B(_09742_), .Y(_09746_));
NAND_g _16119_ (.A(resetn), .B(_09746_), .Y(_09747_));
NOR_g _16120_ (.A(_09745_), .B(_09747_), .Y(_00153_));
NAND_g _16121_ (.A(count_cycle[39]), .B(_09745_), .Y(_09748_));
NOR_g _16122_ (.A(count_cycle[39]), .B(_09745_), .Y(_09749_));
NOR_g _16123_ (.A(_08811_), .B(_09749_), .Y(_09750_));
AND_g _16124_ (.A(_09748_), .B(_09750_), .Y(_00154_));
NOR_g _16125_ (.A(_09053_), .B(_09748_), .Y(_09751_));
NAND_g _16126_ (.A(_09053_), .B(_09748_), .Y(_09752_));
NAND_g _16127_ (.A(resetn), .B(_09752_), .Y(_09753_));
NOR_g _16128_ (.A(_09751_), .B(_09753_), .Y(_00155_));
NAND_g _16129_ (.A(count_cycle[41]), .B(_09751_), .Y(_09754_));
NOR_g _16130_ (.A(count_cycle[41]), .B(_09751_), .Y(_09755_));
NOR_g _16131_ (.A(_08811_), .B(_09755_), .Y(_09756_));
AND_g _16132_ (.A(_09754_), .B(_09756_), .Y(_00156_));
NOR_g _16133_ (.A(_09054_), .B(_09754_), .Y(_09757_));
NAND_g _16134_ (.A(_09054_), .B(_09754_), .Y(_09758_));
NAND_g _16135_ (.A(resetn), .B(_09758_), .Y(_09759_));
NOR_g _16136_ (.A(_09757_), .B(_09759_), .Y(_00157_));
NAND_g _16137_ (.A(count_cycle[43]), .B(_09757_), .Y(_09760_));
NOR_g _16138_ (.A(count_cycle[43]), .B(_09757_), .Y(_09761_));
NOR_g _16139_ (.A(_08811_), .B(_09761_), .Y(_09762_));
AND_g _16140_ (.A(_09760_), .B(_09762_), .Y(_00158_));
NOR_g _16141_ (.A(_09055_), .B(_09760_), .Y(_09763_));
NAND_g _16142_ (.A(_09055_), .B(_09760_), .Y(_09764_));
NAND_g _16143_ (.A(resetn), .B(_09764_), .Y(_09765_));
NOR_g _16144_ (.A(_09763_), .B(_09765_), .Y(_00159_));
NAND_g _16145_ (.A(count_cycle[45]), .B(_09763_), .Y(_09766_));
NOR_g _16146_ (.A(count_cycle[45]), .B(_09763_), .Y(_09767_));
NOR_g _16147_ (.A(_08811_), .B(_09767_), .Y(_09768_));
AND_g _16148_ (.A(_09766_), .B(_09768_), .Y(_00160_));
NOR_g _16149_ (.A(_09056_), .B(_09766_), .Y(_09769_));
NAND_g _16150_ (.A(_09056_), .B(_09766_), .Y(_09770_));
NAND_g _16151_ (.A(resetn), .B(_09770_), .Y(_09771_));
NOR_g _16152_ (.A(_09769_), .B(_09771_), .Y(_00161_));
NAND_g _16153_ (.A(count_cycle[47]), .B(_09769_), .Y(_09772_));
NOR_g _16154_ (.A(count_cycle[47]), .B(_09769_), .Y(_09773_));
NOR_g _16155_ (.A(_08811_), .B(_09773_), .Y(_09774_));
AND_g _16156_ (.A(_09772_), .B(_09774_), .Y(_00162_));
NOR_g _16157_ (.A(_09057_), .B(_09772_), .Y(_09775_));
NAND_g _16158_ (.A(_09057_), .B(_09772_), .Y(_09776_));
NAND_g _16159_ (.A(resetn), .B(_09776_), .Y(_09777_));
NOR_g _16160_ (.A(_09775_), .B(_09777_), .Y(_00163_));
NAND_g _16161_ (.A(count_cycle[49]), .B(_09775_), .Y(_09778_));
NOR_g _16162_ (.A(count_cycle[49]), .B(_09775_), .Y(_09779_));
NOR_g _16163_ (.A(_08811_), .B(_09779_), .Y(_09780_));
AND_g _16164_ (.A(_09778_), .B(_09780_), .Y(_00164_));
NOR_g _16165_ (.A(_09058_), .B(_09778_), .Y(_09781_));
NAND_g _16166_ (.A(_09058_), .B(_09778_), .Y(_09782_));
NAND_g _16167_ (.A(resetn), .B(_09782_), .Y(_09783_));
NOR_g _16168_ (.A(_09781_), .B(_09783_), .Y(_00165_));
NAND_g _16169_ (.A(count_cycle[51]), .B(_09781_), .Y(_09784_));
NOR_g _16170_ (.A(count_cycle[51]), .B(_09781_), .Y(_09785_));
NOR_g _16171_ (.A(_08811_), .B(_09785_), .Y(_09786_));
AND_g _16172_ (.A(_09784_), .B(_09786_), .Y(_00166_));
NOR_g _16173_ (.A(_09059_), .B(_09784_), .Y(_09787_));
NAND_g _16174_ (.A(_09059_), .B(_09784_), .Y(_09788_));
NAND_g _16175_ (.A(resetn), .B(_09788_), .Y(_09789_));
NOR_g _16176_ (.A(_09787_), .B(_09789_), .Y(_00167_));
NAND_g _16177_ (.A(count_cycle[53]), .B(_09787_), .Y(_09790_));
NOR_g _16178_ (.A(count_cycle[53]), .B(_09787_), .Y(_09791_));
NOR_g _16179_ (.A(_08811_), .B(_09791_), .Y(_09792_));
AND_g _16180_ (.A(_09790_), .B(_09792_), .Y(_00168_));
NOR_g _16181_ (.A(_09060_), .B(_09790_), .Y(_09793_));
NAND_g _16182_ (.A(_09060_), .B(_09790_), .Y(_09794_));
NAND_g _16183_ (.A(resetn), .B(_09794_), .Y(_09795_));
NOR_g _16184_ (.A(_09793_), .B(_09795_), .Y(_00169_));
NAND_g _16185_ (.A(count_cycle[55]), .B(_09793_), .Y(_09796_));
NOR_g _16186_ (.A(count_cycle[55]), .B(_09793_), .Y(_09797_));
NOR_g _16187_ (.A(_08811_), .B(_09797_), .Y(_09798_));
AND_g _16188_ (.A(_09796_), .B(_09798_), .Y(_00170_));
NOR_g _16189_ (.A(_09061_), .B(_09796_), .Y(_09799_));
NAND_g _16190_ (.A(_09061_), .B(_09796_), .Y(_09800_));
NAND_g _16191_ (.A(resetn), .B(_09800_), .Y(_09801_));
NOR_g _16192_ (.A(_09799_), .B(_09801_), .Y(_00171_));
NAND_g _16193_ (.A(count_cycle[57]), .B(_09799_), .Y(_09802_));
NOR_g _16194_ (.A(count_cycle[57]), .B(_09799_), .Y(_09803_));
NOR_g _16195_ (.A(_08811_), .B(_09803_), .Y(_09804_));
AND_g _16196_ (.A(_09802_), .B(_09804_), .Y(_00172_));
NOR_g _16197_ (.A(_09062_), .B(_09802_), .Y(_09805_));
NAND_g _16198_ (.A(_09062_), .B(_09802_), .Y(_09806_));
NAND_g _16199_ (.A(resetn), .B(_09806_), .Y(_09807_));
NOR_g _16200_ (.A(_09805_), .B(_09807_), .Y(_00173_));
NAND_g _16201_ (.A(count_cycle[59]), .B(_09805_), .Y(_09808_));
NOR_g _16202_ (.A(count_cycle[59]), .B(_09805_), .Y(_09809_));
NOR_g _16203_ (.A(_08811_), .B(_09809_), .Y(_09810_));
AND_g _16204_ (.A(_09808_), .B(_09810_), .Y(_00174_));
NOR_g _16205_ (.A(_09063_), .B(_09808_), .Y(_09811_));
NAND_g _16206_ (.A(_09063_), .B(_09808_), .Y(_09812_));
NAND_g _16207_ (.A(resetn), .B(_09812_), .Y(_09813_));
NOR_g _16208_ (.A(_09811_), .B(_09813_), .Y(_00175_));
NAND_g _16209_ (.A(count_cycle[61]), .B(_09811_), .Y(_09814_));
NOT_g _16210_ (.A(_09814_), .Y(_09815_));
NOR_g _16211_ (.A(count_cycle[61]), .B(_09811_), .Y(_09816_));
NOR_g _16212_ (.A(_08811_), .B(_09816_), .Y(_09817_));
AND_g _16213_ (.A(_09814_), .B(_09817_), .Y(_00176_));
NAND_g _16214_ (.A(count_cycle[62]), .B(_09815_), .Y(_09818_));
NAND_g _16215_ (.A(_09064_), .B(_09814_), .Y(_09819_));
AND_g _16216_ (.A(resetn), .B(_09819_), .Y(_09820_));
AND_g _16217_ (.A(_09818_), .B(_09820_), .Y(_00177_));
XNOR_g _16218_ (.A(count_cycle[63]), .B(_09818_), .Y(_09821_));
AND_g _16219_ (.A(resetn), .B(_09821_), .Y(_00178_));
NAND_g _16220_ (.A(resetn), .B(cpu_state[7]), .Y(_09822_));
NAND_g _16221_ (.A(_09018_), .B(_09070_), .Y(_09823_));
NOR_g _16222_ (.A(_09822_), .B(_09823_), .Y(_09824_));
AND_g _16223_ (.A(_09069_), .B(_09824_), .Y(_00179_));
NOR_g _16224_ (.A(latched_rd[1]), .B(_09083_), .Y(_09825_));
AND_g _16225_ (.A(_09567_), .B(_09825_), .Y(_09826_));
NAND_g _16226_ (.A(_09567_), .B(_09825_), .Y(_09827_));
NAND_g _16227_ (.A(_09098_), .B(_09826_), .Y(_09828_));
NAND_g _16228_ (.A(cpuregs[1][0]), .B(_09827_), .Y(_09829_));
NAND_g _16229_ (.A(_09828_), .B(_09829_), .Y(_00180_));
NAND_g _16230_ (.A(_09109_), .B(_09826_), .Y(_09830_));
NAND_g _16231_ (.A(cpuregs[1][1]), .B(_09827_), .Y(_09831_));
NAND_g _16232_ (.A(_09830_), .B(_09831_), .Y(_00181_));
NAND_g _16233_ (.A(_09118_), .B(_09826_), .Y(_09832_));
NAND_g _16234_ (.A(cpuregs[1][2]), .B(_09827_), .Y(_09833_));
NAND_g _16235_ (.A(_09832_), .B(_09833_), .Y(_00182_));
NAND_g _16236_ (.A(_09131_), .B(_09826_), .Y(_09834_));
NAND_g _16237_ (.A(cpuregs[1][3]), .B(_09827_), .Y(_09835_));
NAND_g _16238_ (.A(_09834_), .B(_09835_), .Y(_00183_));
NAND_g _16239_ (.A(_09144_), .B(_09826_), .Y(_09836_));
NAND_g _16240_ (.A(cpuregs[1][4]), .B(_09827_), .Y(_09837_));
NAND_g _16241_ (.A(_09836_), .B(_09837_), .Y(_00184_));
NAND_g _16242_ (.A(_09157_), .B(_09826_), .Y(_09838_));
NAND_g _16243_ (.A(cpuregs[1][5]), .B(_09827_), .Y(_09839_));
NAND_g _16244_ (.A(_09838_), .B(_09839_), .Y(_00185_));
NAND_g _16245_ (.A(_09170_), .B(_09826_), .Y(_09840_));
NAND_g _16246_ (.A(cpuregs[1][6]), .B(_09827_), .Y(_09841_));
NAND_g _16247_ (.A(_09840_), .B(_09841_), .Y(_00186_));
NAND_g _16248_ (.A(_09183_), .B(_09826_), .Y(_09842_));
NAND_g _16249_ (.A(cpuregs[1][7]), .B(_09827_), .Y(_09843_));
NAND_g _16250_ (.A(_09842_), .B(_09843_), .Y(_00187_));
NAND_g _16251_ (.A(_09196_), .B(_09826_), .Y(_09844_));
NAND_g _16252_ (.A(cpuregs[1][8]), .B(_09827_), .Y(_09845_));
NAND_g _16253_ (.A(_09844_), .B(_09845_), .Y(_00188_));
NAND_g _16254_ (.A(_09209_), .B(_09826_), .Y(_09846_));
NAND_g _16255_ (.A(cpuregs[1][9]), .B(_09827_), .Y(_09847_));
NAND_g _16256_ (.A(_09846_), .B(_09847_), .Y(_00189_));
NAND_g _16257_ (.A(_09222_), .B(_09826_), .Y(_09848_));
NAND_g _16258_ (.A(cpuregs[1][10]), .B(_09827_), .Y(_09849_));
NAND_g _16259_ (.A(_09848_), .B(_09849_), .Y(_00190_));
NAND_g _16260_ (.A(_09235_), .B(_09826_), .Y(_09850_));
NAND_g _16261_ (.A(cpuregs[1][11]), .B(_09827_), .Y(_09851_));
NAND_g _16262_ (.A(_09850_), .B(_09851_), .Y(_00191_));
NAND_g _16263_ (.A(_09248_), .B(_09826_), .Y(_09852_));
NAND_g _16264_ (.A(cpuregs[1][12]), .B(_09827_), .Y(_09853_));
NAND_g _16265_ (.A(_09852_), .B(_09853_), .Y(_00192_));
NAND_g _16266_ (.A(_09261_), .B(_09826_), .Y(_09854_));
NAND_g _16267_ (.A(cpuregs[1][13]), .B(_09827_), .Y(_09855_));
NAND_g _16268_ (.A(_09854_), .B(_09855_), .Y(_00193_));
NAND_g _16269_ (.A(_09274_), .B(_09826_), .Y(_09856_));
NAND_g _16270_ (.A(cpuregs[1][14]), .B(_09827_), .Y(_09857_));
NAND_g _16271_ (.A(_09856_), .B(_09857_), .Y(_00194_));
NAND_g _16272_ (.A(_09287_), .B(_09826_), .Y(_09858_));
NAND_g _16273_ (.A(cpuregs[1][15]), .B(_09827_), .Y(_09859_));
NAND_g _16274_ (.A(_09858_), .B(_09859_), .Y(_00195_));
NAND_g _16275_ (.A(_09300_), .B(_09826_), .Y(_09860_));
NAND_g _16276_ (.A(cpuregs[1][16]), .B(_09827_), .Y(_09861_));
NAND_g _16277_ (.A(_09860_), .B(_09861_), .Y(_00196_));
NOR_g _16278_ (.A(cpuregs[1][17]), .B(_09826_), .Y(_09862_));
NOR_g _16279_ (.A(_09313_), .B(_09827_), .Y(_09863_));
NOR_g _16280_ (.A(_09862_), .B(_09863_), .Y(_00197_));
NOR_g _16281_ (.A(cpuregs[1][18]), .B(_09826_), .Y(_09864_));
NOR_g _16282_ (.A(_09325_), .B(_09827_), .Y(_09865_));
NOR_g _16283_ (.A(_09864_), .B(_09865_), .Y(_00198_));
NAND_g _16284_ (.A(_09338_), .B(_09826_), .Y(_09866_));
NAND_g _16285_ (.A(cpuregs[1][19]), .B(_09827_), .Y(_09867_));
NAND_g _16286_ (.A(_09866_), .B(_09867_), .Y(_00199_));
NAND_g _16287_ (.A(_09351_), .B(_09826_), .Y(_09868_));
NAND_g _16288_ (.A(cpuregs[1][20]), .B(_09827_), .Y(_09869_));
NAND_g _16289_ (.A(_09868_), .B(_09869_), .Y(_00200_));
NAND_g _16290_ (.A(_09364_), .B(_09826_), .Y(_09870_));
NAND_g _16291_ (.A(cpuregs[1][21]), .B(_09827_), .Y(_09871_));
NAND_g _16292_ (.A(_09870_), .B(_09871_), .Y(_00201_));
NAND_g _16293_ (.A(_09377_), .B(_09826_), .Y(_09872_));
NAND_g _16294_ (.A(cpuregs[1][22]), .B(_09827_), .Y(_09873_));
NAND_g _16295_ (.A(_09872_), .B(_09873_), .Y(_00202_));
NAND_g _16296_ (.A(_09390_), .B(_09826_), .Y(_09874_));
NAND_g _16297_ (.A(cpuregs[1][23]), .B(_09827_), .Y(_09875_));
NAND_g _16298_ (.A(_09874_), .B(_09875_), .Y(_00203_));
NAND_g _16299_ (.A(_09403_), .B(_09826_), .Y(_09876_));
NAND_g _16300_ (.A(cpuregs[1][24]), .B(_09827_), .Y(_09877_));
NAND_g _16301_ (.A(_09876_), .B(_09877_), .Y(_00204_));
NAND_g _16302_ (.A(_09416_), .B(_09826_), .Y(_09878_));
NAND_g _16303_ (.A(cpuregs[1][25]), .B(_09827_), .Y(_09879_));
NAND_g _16304_ (.A(_09878_), .B(_09879_), .Y(_00205_));
NAND_g _16305_ (.A(_09429_), .B(_09826_), .Y(_09880_));
NAND_g _16306_ (.A(cpuregs[1][26]), .B(_09827_), .Y(_09881_));
NAND_g _16307_ (.A(_09880_), .B(_09881_), .Y(_00206_));
NAND_g _16308_ (.A(_09442_), .B(_09826_), .Y(_09882_));
NAND_g _16309_ (.A(cpuregs[1][27]), .B(_09827_), .Y(_09883_));
NAND_g _16310_ (.A(_09882_), .B(_09883_), .Y(_00207_));
NAND_g _16311_ (.A(_09455_), .B(_09826_), .Y(_09884_));
NAND_g _16312_ (.A(cpuregs[1][28]), .B(_09827_), .Y(_09885_));
NAND_g _16313_ (.A(_09884_), .B(_09885_), .Y(_00208_));
NAND_g _16314_ (.A(_09468_), .B(_09826_), .Y(_09886_));
NAND_g _16315_ (.A(cpuregs[1][29]), .B(_09827_), .Y(_09887_));
NAND_g _16316_ (.A(_09886_), .B(_09887_), .Y(_00209_));
NAND_g _16317_ (.A(_09481_), .B(_09826_), .Y(_09888_));
NAND_g _16318_ (.A(cpuregs[1][30]), .B(_09827_), .Y(_09889_));
NAND_g _16319_ (.A(_09888_), .B(_09889_), .Y(_00210_));
NAND_g _16320_ (.A(_09493_), .B(_09826_), .Y(_09890_));
NAND_g _16321_ (.A(cpuregs[1][31]), .B(_09827_), .Y(_09891_));
NAND_g _16322_ (.A(_09890_), .B(_09891_), .Y(_00211_));
NAND_g _16323_ (.A(_08857_), .B(decoder_trigger), .Y(_09892_));
AND_g _16324_ (.A(decoder_trigger), .B(_09073_), .Y(_09893_));
AND_g _16325_ (.A(_08857_), .B(_09893_), .Y(_09894_));
NAND_g _16326_ (.A(resetn), .B(_09894_), .Y(_09895_));
NAND_g _16327_ (.A(_08807_), .B(_09895_), .Y(_09896_));
AND_g _16328_ (.A(mem_state[0]), .B(mem_state[1]), .Y(_09897_));
NAND_g _16329_ (.A(mem_do_rinst), .B(_09897_), .Y(_09898_));
NOR_g _16330_ (.A(mem_do_rdata), .B(mem_do_rinst), .Y(_09899_));
NAND_g _16331_ (.A(_08789_), .B(_09899_), .Y(_09900_));
NOR_g _16332_ (.A(mem_state[0]), .B(mem_state[1]), .Y(_09901_));
NOT_g _16333_ (.A(_09901_), .Y(_09902_));
AND_g _16334_ (.A(mem_valid), .B(mem_ready), .Y(_09903_));
NAND_g _16335_ (.A(mem_valid), .B(mem_ready), .Y(_09904_));
NOR_g _16336_ (.A(_09901_), .B(_09904_), .Y(_09905_));
NAND_g _16337_ (.A(_09900_), .B(_09905_), .Y(_09906_));
AND_g _16338_ (.A(_09898_), .B(_09906_), .Y(_09907_));
NAND_g _16339_ (.A(_09898_), .B(_09906_), .Y(_09908_));
AND_g _16340_ (.A(resetn), .B(_09907_), .Y(_09909_));
NAND_g _16341_ (.A(resetn), .B(_09907_), .Y(_09910_));
AND_g _16342_ (.A(_09896_), .B(_09909_), .Y(_09911_));
NAND_g _16343_ (.A(instr_jalr), .B(_09894_), .Y(_09912_));
AND_g _16344_ (.A(_09911_), .B(_09912_), .Y(_00212_));
AND_g _16345_ (.A(latched_branch), .B(latched_store), .Y(_09913_));
NAND_g _16346_ (.A(latched_branch), .B(latched_store), .Y(_09914_));
NAND_g _16347_ (.A(_09105_), .B(_09913_), .Y(_09915_));
NAND_g _16348_ (.A(reg_next_pc[1]), .B(_09914_), .Y(_09916_));
NAND_g _16349_ (.A(_09915_), .B(_09916_), .Y(_09917_));
AND_g _16350_ (.A(_09075_), .B(_09917_), .Y(_09918_));
NOT_g _16351_ (.A(_09918_), .Y(_09919_));
AND_g _16352_ (.A(resetn), .B(_09074_), .Y(_09920_));
NAND_g _16353_ (.A(reg_pc[1]), .B(_09920_), .Y(_09921_));
NAND_g _16354_ (.A(_09919_), .B(_09921_), .Y(_00213_));
NAND_g _16355_ (.A(reg_next_pc[2]), .B(_09914_), .Y(_09922_));
NAND_g _16356_ (.A(_09114_), .B(_09913_), .Y(_09923_));
NAND_g _16357_ (.A(_09922_), .B(_09923_), .Y(_09924_));
AND_g _16358_ (.A(_09075_), .B(_09924_), .Y(_09925_));
NAND_g _16359_ (.A(_09075_), .B(_09924_), .Y(_09926_));
NAND_g _16360_ (.A(reg_pc[2]), .B(_09920_), .Y(_09927_));
NAND_g _16361_ (.A(_09926_), .B(_09927_), .Y(_00214_));
NAND_g _16362_ (.A(reg_next_pc[3]), .B(_09914_), .Y(_09928_));
NAND_g _16363_ (.A(_09123_), .B(_09913_), .Y(_09929_));
NAND_g _16364_ (.A(_09928_), .B(_09929_), .Y(_09930_));
AND_g _16365_ (.A(_09075_), .B(_09930_), .Y(_09931_));
NAND_g _16366_ (.A(_09075_), .B(_09930_), .Y(_09932_));
NAND_g _16367_ (.A(reg_pc[3]), .B(_09920_), .Y(_09933_));
NAND_g _16368_ (.A(_09932_), .B(_09933_), .Y(_00215_));
NAND_g _16369_ (.A(reg_next_pc[4]), .B(_09914_), .Y(_09934_));
NAND_g _16370_ (.A(_09136_), .B(_09913_), .Y(_09935_));
NAND_g _16371_ (.A(_09934_), .B(_09935_), .Y(_09936_));
AND_g _16372_ (.A(_09075_), .B(_09936_), .Y(_09937_));
NAND_g _16373_ (.A(_09075_), .B(_09936_), .Y(_09938_));
NAND_g _16374_ (.A(reg_pc[4]), .B(_09920_), .Y(_09939_));
NAND_g _16375_ (.A(_09938_), .B(_09939_), .Y(_00216_));
NAND_g _16376_ (.A(reg_next_pc[5]), .B(_09914_), .Y(_09940_));
NAND_g _16377_ (.A(_09149_), .B(_09913_), .Y(_09941_));
NAND_g _16378_ (.A(_09940_), .B(_09941_), .Y(_09942_));
AND_g _16379_ (.A(_09075_), .B(_09942_), .Y(_09943_));
NAND_g _16380_ (.A(_09075_), .B(_09942_), .Y(_09944_));
NAND_g _16381_ (.A(reg_pc[5]), .B(_09920_), .Y(_09945_));
NAND_g _16382_ (.A(_09944_), .B(_09945_), .Y(_00217_));
NAND_g _16383_ (.A(reg_next_pc[6]), .B(_09914_), .Y(_09946_));
NAND_g _16384_ (.A(_09162_), .B(_09913_), .Y(_09947_));
NAND_g _16385_ (.A(_09946_), .B(_09947_), .Y(_09948_));
AND_g _16386_ (.A(_09075_), .B(_09948_), .Y(_09949_));
NOT_g _16387_ (.A(_09949_), .Y(_09950_));
NAND_g _16388_ (.A(reg_pc[6]), .B(_09920_), .Y(_09951_));
NAND_g _16389_ (.A(_09950_), .B(_09951_), .Y(_00218_));
NAND_g _16390_ (.A(reg_next_pc[7]), .B(_09914_), .Y(_09952_));
NAND_g _16391_ (.A(_09175_), .B(_09913_), .Y(_09953_));
NAND_g _16392_ (.A(_09952_), .B(_09953_), .Y(_09954_));
AND_g _16393_ (.A(_09075_), .B(_09954_), .Y(_09955_));
NAND_g _16394_ (.A(_09075_), .B(_09954_), .Y(_09956_));
NAND_g _16395_ (.A(reg_pc[7]), .B(_09920_), .Y(_09957_));
NAND_g _16396_ (.A(_09956_), .B(_09957_), .Y(_00219_));
NAND_g _16397_ (.A(reg_next_pc[8]), .B(_09914_), .Y(_09958_));
NAND_g _16398_ (.A(_09188_), .B(_09913_), .Y(_09959_));
NAND_g _16399_ (.A(_09958_), .B(_09959_), .Y(_09960_));
AND_g _16400_ (.A(_09075_), .B(_09960_), .Y(_09961_));
NOT_g _16401_ (.A(_09961_), .Y(_09962_));
NAND_g _16402_ (.A(reg_pc[8]), .B(_09920_), .Y(_09963_));
NAND_g _16403_ (.A(_09962_), .B(_09963_), .Y(_00220_));
NAND_g _16404_ (.A(reg_next_pc[9]), .B(_09914_), .Y(_09964_));
NAND_g _16405_ (.A(_09201_), .B(_09913_), .Y(_09965_));
NAND_g _16406_ (.A(_09964_), .B(_09965_), .Y(_09966_));
AND_g _16407_ (.A(_09075_), .B(_09966_), .Y(_09967_));
NAND_g _16408_ (.A(_09075_), .B(_09966_), .Y(_09968_));
NAND_g _16409_ (.A(reg_pc[9]), .B(_09920_), .Y(_09969_));
NAND_g _16410_ (.A(_09968_), .B(_09969_), .Y(_00221_));
NAND_g _16411_ (.A(reg_next_pc[10]), .B(_09914_), .Y(_09970_));
NAND_g _16412_ (.A(_09214_), .B(_09913_), .Y(_09971_));
NAND_g _16413_ (.A(_09970_), .B(_09971_), .Y(_09972_));
AND_g _16414_ (.A(_09075_), .B(_09972_), .Y(_09973_));
NOT_g _16415_ (.A(_09973_), .Y(_09974_));
NAND_g _16416_ (.A(reg_pc[10]), .B(_09920_), .Y(_09975_));
NAND_g _16417_ (.A(_09974_), .B(_09975_), .Y(_00222_));
NAND_g _16418_ (.A(reg_next_pc[11]), .B(_09914_), .Y(_09976_));
NAND_g _16419_ (.A(_09227_), .B(_09913_), .Y(_09977_));
NAND_g _16420_ (.A(_09976_), .B(_09977_), .Y(_09978_));
AND_g _16421_ (.A(_09075_), .B(_09978_), .Y(_09979_));
NAND_g _16422_ (.A(_09075_), .B(_09978_), .Y(_09980_));
NAND_g _16423_ (.A(reg_pc[11]), .B(_09920_), .Y(_09981_));
NAND_g _16424_ (.A(_09980_), .B(_09981_), .Y(_00223_));
NAND_g _16425_ (.A(reg_next_pc[12]), .B(_09914_), .Y(_09982_));
NAND_g _16426_ (.A(_09240_), .B(_09913_), .Y(_09983_));
NAND_g _16427_ (.A(_09982_), .B(_09983_), .Y(_09984_));
AND_g _16428_ (.A(_09075_), .B(_09984_), .Y(_09985_));
NOT_g _16429_ (.A(_09985_), .Y(_09986_));
NAND_g _16430_ (.A(reg_pc[12]), .B(_09920_), .Y(_09987_));
NAND_g _16431_ (.A(_09986_), .B(_09987_), .Y(_00224_));
NAND_g _16432_ (.A(reg_next_pc[13]), .B(_09914_), .Y(_09988_));
NAND_g _16433_ (.A(_09253_), .B(_09913_), .Y(_09989_));
NAND_g _16434_ (.A(_09988_), .B(_09989_), .Y(_09990_));
AND_g _16435_ (.A(_09075_), .B(_09990_), .Y(_09991_));
NAND_g _16436_ (.A(_09075_), .B(_09990_), .Y(_09992_));
NAND_g _16437_ (.A(reg_pc[13]), .B(_09920_), .Y(_09993_));
NAND_g _16438_ (.A(_09992_), .B(_09993_), .Y(_00225_));
NAND_g _16439_ (.A(reg_next_pc[14]), .B(_09914_), .Y(_09994_));
NAND_g _16440_ (.A(_09266_), .B(_09913_), .Y(_09995_));
NAND_g _16441_ (.A(_09994_), .B(_09995_), .Y(_09996_));
AND_g _16442_ (.A(_09075_), .B(_09996_), .Y(_09997_));
NOT_g _16443_ (.A(_09997_), .Y(_09998_));
NAND_g _16444_ (.A(reg_pc[14]), .B(_09920_), .Y(_09999_));
NAND_g _16445_ (.A(_09998_), .B(_09999_), .Y(_00226_));
NAND_g _16446_ (.A(reg_next_pc[15]), .B(_09914_), .Y(_10000_));
NAND_g _16447_ (.A(_09279_), .B(_09913_), .Y(_10001_));
NAND_g _16448_ (.A(_10000_), .B(_10001_), .Y(_10002_));
AND_g _16449_ (.A(_09075_), .B(_10002_), .Y(_10003_));
NAND_g _16450_ (.A(_09075_), .B(_10002_), .Y(_10004_));
NAND_g _16451_ (.A(reg_pc[15]), .B(_09920_), .Y(_10005_));
NAND_g _16452_ (.A(_10004_), .B(_10005_), .Y(_00227_));
NAND_g _16453_ (.A(reg_next_pc[16]), .B(_09914_), .Y(_10006_));
NAND_g _16454_ (.A(_09292_), .B(_09913_), .Y(_10007_));
NAND_g _16455_ (.A(_10006_), .B(_10007_), .Y(_10008_));
AND_g _16456_ (.A(_09075_), .B(_10008_), .Y(_10009_));
NOT_g _16457_ (.A(_10009_), .Y(_10010_));
NAND_g _16458_ (.A(reg_pc[16]), .B(_09920_), .Y(_10011_));
NAND_g _16459_ (.A(_10010_), .B(_10011_), .Y(_00228_));
NAND_g _16460_ (.A(reg_next_pc[17]), .B(_09914_), .Y(_10012_));
NAND_g _16461_ (.A(_09305_), .B(_09913_), .Y(_10013_));
NAND_g _16462_ (.A(_10012_), .B(_10013_), .Y(_10014_));
AND_g _16463_ (.A(_09075_), .B(_10014_), .Y(_10015_));
NAND_g _16464_ (.A(_09075_), .B(_10014_), .Y(_10016_));
NAND_g _16465_ (.A(reg_pc[17]), .B(_09920_), .Y(_10017_));
NAND_g _16466_ (.A(_10016_), .B(_10017_), .Y(_00229_));
NAND_g _16467_ (.A(reg_next_pc[18]), .B(_09914_), .Y(_10018_));
NAND_g _16468_ (.A(_09317_), .B(_09913_), .Y(_10019_));
NAND_g _16469_ (.A(_10018_), .B(_10019_), .Y(_10020_));
AND_g _16470_ (.A(_09075_), .B(_10020_), .Y(_10021_));
NOT_g _16471_ (.A(_10021_), .Y(_10022_));
NAND_g _16472_ (.A(reg_pc[18]), .B(_09920_), .Y(_10023_));
NAND_g _16473_ (.A(_10022_), .B(_10023_), .Y(_00230_));
NAND_g _16474_ (.A(reg_next_pc[19]), .B(_09914_), .Y(_10024_));
NAND_g _16475_ (.A(_09330_), .B(_09913_), .Y(_10025_));
NAND_g _16476_ (.A(_10024_), .B(_10025_), .Y(_10026_));
NAND_g _16477_ (.A(_09075_), .B(_10026_), .Y(_10027_));
NOT_g _16478_ (.A(_10027_), .Y(_10028_));
NAND_g _16479_ (.A(reg_pc[19]), .B(_09920_), .Y(_10029_));
NAND_g _16480_ (.A(_10027_), .B(_10029_), .Y(_00231_));
NAND_g _16481_ (.A(reg_next_pc[20]), .B(_09914_), .Y(_10030_));
NAND_g _16482_ (.A(_09343_), .B(_09913_), .Y(_10031_));
NAND_g _16483_ (.A(_10030_), .B(_10031_), .Y(_10032_));
AND_g _16484_ (.A(_09075_), .B(_10032_), .Y(_10033_));
NOT_g _16485_ (.A(_10033_), .Y(_10034_));
NAND_g _16486_ (.A(reg_pc[20]), .B(_09920_), .Y(_10035_));
NAND_g _16487_ (.A(_10034_), .B(_10035_), .Y(_00232_));
NAND_g _16488_ (.A(reg_next_pc[21]), .B(_09914_), .Y(_10036_));
NAND_g _16489_ (.A(_09356_), .B(_09913_), .Y(_10037_));
NAND_g _16490_ (.A(_10036_), .B(_10037_), .Y(_10038_));
NAND_g _16491_ (.A(_09075_), .B(_10038_), .Y(_10039_));
NOT_g _16492_ (.A(_10039_), .Y(_10040_));
NAND_g _16493_ (.A(reg_pc[21]), .B(_09920_), .Y(_10041_));
NAND_g _16494_ (.A(_10039_), .B(_10041_), .Y(_00233_));
NAND_g _16495_ (.A(reg_next_pc[22]), .B(_09914_), .Y(_10042_));
NAND_g _16496_ (.A(_09369_), .B(_09913_), .Y(_10043_));
NAND_g _16497_ (.A(_10042_), .B(_10043_), .Y(_10044_));
AND_g _16498_ (.A(_09075_), .B(_10044_), .Y(_10045_));
NOT_g _16499_ (.A(_10045_), .Y(_10046_));
NAND_g _16500_ (.A(reg_pc[22]), .B(_09920_), .Y(_10047_));
NAND_g _16501_ (.A(_10046_), .B(_10047_), .Y(_00234_));
NAND_g _16502_ (.A(reg_next_pc[23]), .B(_09914_), .Y(_10048_));
NAND_g _16503_ (.A(_09382_), .B(_09913_), .Y(_10049_));
NAND_g _16504_ (.A(_10048_), .B(_10049_), .Y(_10050_));
NAND_g _16505_ (.A(_09075_), .B(_10050_), .Y(_10051_));
NOT_g _16506_ (.A(_10051_), .Y(_10052_));
NAND_g _16507_ (.A(reg_pc[23]), .B(_09920_), .Y(_10053_));
NAND_g _16508_ (.A(_10051_), .B(_10053_), .Y(_00235_));
NAND_g _16509_ (.A(reg_next_pc[24]), .B(_09914_), .Y(_10054_));
NAND_g _16510_ (.A(_09395_), .B(_09913_), .Y(_10055_));
NAND_g _16511_ (.A(_10054_), .B(_10055_), .Y(_10056_));
AND_g _16512_ (.A(_09075_), .B(_10056_), .Y(_10057_));
NAND_g _16513_ (.A(_09075_), .B(_10056_), .Y(_10058_));
NAND_g _16514_ (.A(reg_pc[24]), .B(_09920_), .Y(_10059_));
NAND_g _16515_ (.A(_10058_), .B(_10059_), .Y(_00236_));
NAND_g _16516_ (.A(reg_next_pc[25]), .B(_09914_), .Y(_10060_));
NAND_g _16517_ (.A(_09408_), .B(_09913_), .Y(_10061_));
NAND_g _16518_ (.A(_10060_), .B(_10061_), .Y(_10062_));
NAND_g _16519_ (.A(_09075_), .B(_10062_), .Y(_10063_));
NAND_g _16520_ (.A(reg_pc[25]), .B(_09920_), .Y(_10064_));
NAND_g _16521_ (.A(_10063_), .B(_10064_), .Y(_00237_));
NAND_g _16522_ (.A(reg_next_pc[26]), .B(_09914_), .Y(_10065_));
NAND_g _16523_ (.A(_09421_), .B(_09913_), .Y(_10066_));
NAND_g _16524_ (.A(_10065_), .B(_10066_), .Y(_10067_));
AND_g _16525_ (.A(_09075_), .B(_10067_), .Y(_10068_));
NAND_g _16526_ (.A(_09075_), .B(_10067_), .Y(_10069_));
NAND_g _16527_ (.A(reg_pc[26]), .B(_09920_), .Y(_10070_));
NAND_g _16528_ (.A(_10069_), .B(_10070_), .Y(_00238_));
NAND_g _16529_ (.A(reg_next_pc[27]), .B(_09914_), .Y(_10071_));
NAND_g _16530_ (.A(_09434_), .B(_09913_), .Y(_10072_));
NAND_g _16531_ (.A(_10071_), .B(_10072_), .Y(_10073_));
NAND_g _16532_ (.A(_09075_), .B(_10073_), .Y(_10074_));
NAND_g _16533_ (.A(reg_pc[27]), .B(_09920_), .Y(_10075_));
NAND_g _16534_ (.A(_10074_), .B(_10075_), .Y(_00239_));
NAND_g _16535_ (.A(reg_next_pc[28]), .B(_09914_), .Y(_10076_));
NAND_g _16536_ (.A(_09447_), .B(_09913_), .Y(_10077_));
NAND_g _16537_ (.A(_10076_), .B(_10077_), .Y(_10078_));
AND_g _16538_ (.A(_09075_), .B(_10078_), .Y(_10079_));
NOT_g _16539_ (.A(_10079_), .Y(_10080_));
NAND_g _16540_ (.A(reg_pc[28]), .B(_09920_), .Y(_10081_));
NAND_g _16541_ (.A(_10080_), .B(_10081_), .Y(_00240_));
NAND_g _16542_ (.A(reg_next_pc[29]), .B(_09914_), .Y(_10082_));
NAND_g _16543_ (.A(_09460_), .B(_09913_), .Y(_10083_));
NAND_g _16544_ (.A(_10082_), .B(_10083_), .Y(_10084_));
AND_g _16545_ (.A(_09075_), .B(_10084_), .Y(_10085_));
NAND_g _16546_ (.A(_09075_), .B(_10084_), .Y(_10086_));
NAND_g _16547_ (.A(reg_pc[29]), .B(_09920_), .Y(_10087_));
NAND_g _16548_ (.A(_10086_), .B(_10087_), .Y(_00241_));
NAND_g _16549_ (.A(reg_next_pc[30]), .B(_09914_), .Y(_10088_));
NAND_g _16550_ (.A(_09473_), .B(_09913_), .Y(_10089_));
NAND_g _16551_ (.A(_10088_), .B(_10089_), .Y(_10090_));
NAND_g _16552_ (.A(_09075_), .B(_10090_), .Y(_10091_));
NAND_g _16553_ (.A(reg_pc[30]), .B(_09920_), .Y(_10092_));
NAND_g _16554_ (.A(_10091_), .B(_10092_), .Y(_00242_));
NAND_g _16555_ (.A(reg_next_pc[31]), .B(_09914_), .Y(_10093_));
NAND_g _16556_ (.A(_09486_), .B(_09913_), .Y(_10094_));
NAND_g _16557_ (.A(_10093_), .B(_10094_), .Y(_10095_));
NAND_g _16558_ (.A(_09075_), .B(_10095_), .Y(_10096_));
NAND_g _16559_ (.A(reg_pc[31]), .B(_09920_), .Y(_10097_));
NAND_g _16560_ (.A(_10096_), .B(_10097_), .Y(_00243_));
NAND_g _16561_ (.A(reg_next_pc[1]), .B(_09920_), .Y(_10098_));
AND_g _16562_ (.A(instr_jal), .B(decoded_imm_j[1]), .Y(_10099_));
NAND_g _16563_ (.A(decoder_trigger), .B(_10099_), .Y(_10100_));
XNOR_g _16564_ (.A(_09917_), .B(_10100_), .Y(_10101_));
NAND_g _16565_ (.A(_09075_), .B(_10101_), .Y(_10102_));
NAND_g _16566_ (.A(_10098_), .B(_10102_), .Y(_00244_));
AND_g _16567_ (.A(decoded_imm_j[1]), .B(_09918_), .Y(_10103_));
NAND_g _16568_ (.A(decoded_imm_j[2]), .B(_09925_), .Y(_10104_));
XNOR_g _16569_ (.A(decoded_imm_j[2]), .B(_09926_), .Y(_10105_));
NAND_g _16570_ (.A(_10103_), .B(_10105_), .Y(_10106_));
XOR_g _16571_ (.A(_10103_), .B(_10105_), .Y(_10107_));
NAND_g _16572_ (.A(_08857_), .B(_09926_), .Y(_10108_));
AND_g _16573_ (.A(decoder_trigger), .B(_10108_), .Y(_10109_));
NAND_g _16574_ (.A(instr_jal), .B(_10107_), .Y(_10110_));
NAND_g _16575_ (.A(_10109_), .B(_10110_), .Y(_10111_));
NAND_g _16576_ (.A(resetn), .B(_09893_), .Y(_10112_));
NAND_g _16577_ (.A(_09926_), .B(_10112_), .Y(_10113_));
NAND_g _16578_ (.A(_10111_), .B(_10113_), .Y(_10114_));
NAND_g _16579_ (.A(reg_next_pc[2]), .B(_09920_), .Y(_10115_));
NAND_g _16580_ (.A(_10114_), .B(_10115_), .Y(_00245_));
NAND_g _16581_ (.A(reg_next_pc[3]), .B(_09920_), .Y(_10116_));
NAND_g _16582_ (.A(_10104_), .B(_10106_), .Y(_10117_));
NAND_g _16583_ (.A(decoded_imm_j[3]), .B(_09931_), .Y(_10118_));
XNOR_g _16584_ (.A(decoded_imm_j[3]), .B(_09932_), .Y(_10119_));
NAND_g _16585_ (.A(_10117_), .B(_10119_), .Y(_10120_));
XOR_g _16586_ (.A(_10117_), .B(_10119_), .Y(_10121_));
NAND_g _16587_ (.A(instr_jal), .B(_10121_), .Y(_10122_));
AND_g _16588_ (.A(_09924_), .B(_09931_), .Y(_10123_));
AND_g _16589_ (.A(_09926_), .B(_09932_), .Y(_10124_));
AND_g _16590_ (.A(_09925_), .B(_09930_), .Y(_10125_));
NOR_g _16591_ (.A(_10123_), .B(_10124_), .Y(_10126_));
NAND_g _16592_ (.A(_08857_), .B(_10126_), .Y(_10127_));
AND_g _16593_ (.A(decoder_trigger), .B(_10127_), .Y(_10128_));
NAND_g _16594_ (.A(_10122_), .B(_10128_), .Y(_10129_));
NAND_g _16595_ (.A(_09932_), .B(_10112_), .Y(_10130_));
NAND_g _16596_ (.A(_10129_), .B(_10130_), .Y(_10131_));
NAND_g _16597_ (.A(_10116_), .B(_10131_), .Y(_00246_));
NAND_g _16598_ (.A(reg_next_pc[4]), .B(_09920_), .Y(_10132_));
NAND_g _16599_ (.A(_10118_), .B(_10120_), .Y(_10133_));
NAND_g _16600_ (.A(decoded_imm_j[4]), .B(_09937_), .Y(_10134_));
XNOR_g _16601_ (.A(_08879_), .B(_09937_), .Y(_10135_));
NAND_g _16602_ (.A(_10133_), .B(_10135_), .Y(_10136_));
XOR_g _16603_ (.A(_10133_), .B(_10135_), .Y(_10137_));
NAND_g _16604_ (.A(instr_jal), .B(_10137_), .Y(_10138_));
AND_g _16605_ (.A(_09936_), .B(_10123_), .Y(_10139_));
AND_g _16606_ (.A(_09937_), .B(_10125_), .Y(_10140_));
XNOR_g _16607_ (.A(_09938_), .B(_10123_), .Y(_10141_));
NAND_g _16608_ (.A(_08857_), .B(_10141_), .Y(_10142_));
AND_g _16609_ (.A(decoder_trigger), .B(_10142_), .Y(_10143_));
NAND_g _16610_ (.A(_10138_), .B(_10143_), .Y(_10144_));
NAND_g _16611_ (.A(_09938_), .B(_10112_), .Y(_10145_));
NAND_g _16612_ (.A(_10144_), .B(_10145_), .Y(_10146_));
NAND_g _16613_ (.A(_10132_), .B(_10146_), .Y(_00247_));
NAND_g _16614_ (.A(reg_next_pc[5]), .B(_09920_), .Y(_10147_));
NAND_g _16615_ (.A(_10134_), .B(_10136_), .Y(_10148_));
NAND_g _16616_ (.A(decoded_imm_j[5]), .B(_09943_), .Y(_10149_));
XNOR_g _16617_ (.A(decoded_imm_j[5]), .B(_09944_), .Y(_10150_));
NAND_g _16618_ (.A(_10148_), .B(_10150_), .Y(_10151_));
XOR_g _16619_ (.A(_10148_), .B(_10150_), .Y(_10152_));
NOR_g _16620_ (.A(_09943_), .B(_10140_), .Y(_10153_));
AND_g _16621_ (.A(_09942_), .B(_10139_), .Y(_10154_));
AND_g _16622_ (.A(_09942_), .B(_10140_), .Y(_10155_));
NOR_g _16623_ (.A(_10153_), .B(_10155_), .Y(_10156_));
NAND_g _16624_ (.A(_08857_), .B(_10156_), .Y(_10157_));
AND_g _16625_ (.A(decoder_trigger), .B(_10157_), .Y(_10158_));
NAND_g _16626_ (.A(instr_jal), .B(_10152_), .Y(_10159_));
NAND_g _16627_ (.A(_10158_), .B(_10159_), .Y(_10160_));
NAND_g _16628_ (.A(_09944_), .B(_10112_), .Y(_10161_));
NAND_g _16629_ (.A(_10160_), .B(_10161_), .Y(_10162_));
NAND_g _16630_ (.A(_10147_), .B(_10162_), .Y(_00248_));
NAND_g _16631_ (.A(reg_next_pc[6]), .B(_09920_), .Y(_10163_));
NAND_g _16632_ (.A(_10149_), .B(_10151_), .Y(_10164_));
NAND_g _16633_ (.A(decoded_imm_j[6]), .B(_09949_), .Y(_10165_));
XOR_g _16634_ (.A(decoded_imm_j[6]), .B(_09949_), .Y(_10166_));
NAND_g _16635_ (.A(_10164_), .B(_10166_), .Y(_10167_));
XOR_g _16636_ (.A(_10164_), .B(_10166_), .Y(_10168_));
NAND_g _16637_ (.A(instr_jal), .B(_10168_), .Y(_10169_));
AND_g _16638_ (.A(_09949_), .B(_10154_), .Y(_10170_));
AND_g _16639_ (.A(_09949_), .B(_10155_), .Y(_10171_));
XNOR_g _16640_ (.A(_09950_), .B(_10155_), .Y(_10172_));
NAND_g _16641_ (.A(_08857_), .B(_10172_), .Y(_10173_));
AND_g _16642_ (.A(decoder_trigger), .B(_10173_), .Y(_10174_));
NAND_g _16643_ (.A(_10169_), .B(_10174_), .Y(_10175_));
NAND_g _16644_ (.A(_09950_), .B(_10112_), .Y(_10176_));
NAND_g _16645_ (.A(_10175_), .B(_10176_), .Y(_10177_));
NAND_g _16646_ (.A(_10163_), .B(_10177_), .Y(_00249_));
NAND_g _16647_ (.A(reg_next_pc[7]), .B(_09920_), .Y(_10178_));
AND_g _16648_ (.A(_10165_), .B(_10167_), .Y(_10179_));
NAND_g _16649_ (.A(decoded_imm_j[7]), .B(_09955_), .Y(_10180_));
NOR_g _16650_ (.A(decoded_imm_j[7]), .B(_09955_), .Y(_10181_));
XNOR_g _16651_ (.A(decoded_imm_j[7]), .B(_09956_), .Y(_10182_));
XNOR_g _16652_ (.A(_10179_), .B(_10182_), .Y(_10183_));
NAND_g _16653_ (.A(instr_jal), .B(_10183_), .Y(_10184_));
AND_g _16654_ (.A(_09954_), .B(_10170_), .Y(_10185_));
NOR_g _16655_ (.A(_09955_), .B(_10171_), .Y(_10186_));
AND_g _16656_ (.A(_09954_), .B(_10171_), .Y(_10187_));
NOR_g _16657_ (.A(_10186_), .B(_10187_), .Y(_10188_));
NAND_g _16658_ (.A(_08857_), .B(_10188_), .Y(_10189_));
AND_g _16659_ (.A(decoder_trigger), .B(_10189_), .Y(_10190_));
NAND_g _16660_ (.A(_10184_), .B(_10190_), .Y(_10191_));
NAND_g _16661_ (.A(_09956_), .B(_10112_), .Y(_10192_));
NAND_g _16662_ (.A(_10191_), .B(_10192_), .Y(_10193_));
NAND_g _16663_ (.A(_10178_), .B(_10193_), .Y(_00250_));
NAND_g _16664_ (.A(reg_next_pc[8]), .B(_09920_), .Y(_10194_));
NAND_g _16665_ (.A(decoded_imm_j[8]), .B(_09961_), .Y(_10195_));
XOR_g _16666_ (.A(decoded_imm_j[8]), .B(_09961_), .Y(_10196_));
AND_g _16667_ (.A(_10179_), .B(_10180_), .Y(_10197_));
NOR_g _16668_ (.A(_10181_), .B(_10197_), .Y(_10198_));
NAND_g _16669_ (.A(_10196_), .B(_10198_), .Y(_10199_));
XOR_g _16670_ (.A(_10196_), .B(_10198_), .Y(_10200_));
NAND_g _16671_ (.A(instr_jal), .B(_10200_), .Y(_10201_));
AND_g _16672_ (.A(_09961_), .B(_10185_), .Y(_10202_));
AND_g _16673_ (.A(_09961_), .B(_10187_), .Y(_10203_));
XNOR_g _16674_ (.A(_09962_), .B(_10187_), .Y(_10204_));
NAND_g _16675_ (.A(_08857_), .B(_10204_), .Y(_10205_));
AND_g _16676_ (.A(decoder_trigger), .B(_10205_), .Y(_10206_));
NAND_g _16677_ (.A(_10201_), .B(_10206_), .Y(_10207_));
NAND_g _16678_ (.A(_09962_), .B(_10112_), .Y(_10208_));
AND_g _16679_ (.A(_10207_), .B(_10208_), .Y(_10209_));
NOT_g _16680_ (.A(_10209_), .Y(_10210_));
NAND_g _16681_ (.A(_10194_), .B(_10210_), .Y(_00251_));
NAND_g _16682_ (.A(reg_next_pc[9]), .B(_09920_), .Y(_10211_));
AND_g _16683_ (.A(_10195_), .B(_10199_), .Y(_10212_));
NAND_g _16684_ (.A(decoded_imm_j[9]), .B(_09967_), .Y(_10213_));
NOR_g _16685_ (.A(decoded_imm_j[9]), .B(_09967_), .Y(_10214_));
XNOR_g _16686_ (.A(decoded_imm_j[9]), .B(_09968_), .Y(_10215_));
XNOR_g _16687_ (.A(_10212_), .B(_10215_), .Y(_10216_));
NAND_g _16688_ (.A(instr_jal), .B(_10216_), .Y(_10217_));
NOR_g _16689_ (.A(_09967_), .B(_10202_), .Y(_10218_));
AND_g _16690_ (.A(_09966_), .B(_10202_), .Y(_10219_));
AND_g _16691_ (.A(_09966_), .B(_10203_), .Y(_10220_));
NOR_g _16692_ (.A(_10218_), .B(_10220_), .Y(_10221_));
NAND_g _16693_ (.A(_08857_), .B(_10221_), .Y(_10222_));
AND_g _16694_ (.A(decoder_trigger), .B(_10222_), .Y(_10223_));
NAND_g _16695_ (.A(_10217_), .B(_10223_), .Y(_10224_));
NAND_g _16696_ (.A(_09968_), .B(_10112_), .Y(_10225_));
NAND_g _16697_ (.A(_10224_), .B(_10225_), .Y(_10226_));
NAND_g _16698_ (.A(_10211_), .B(_10226_), .Y(_00252_));
NAND_g _16699_ (.A(reg_next_pc[10]), .B(_09920_), .Y(_10227_));
NAND_g _16700_ (.A(decoded_imm_j[10]), .B(_09973_), .Y(_10228_));
XOR_g _16701_ (.A(decoded_imm_j[10]), .B(_09973_), .Y(_10229_));
AND_g _16702_ (.A(_10212_), .B(_10213_), .Y(_10230_));
NOR_g _16703_ (.A(_10214_), .B(_10230_), .Y(_10231_));
NAND_g _16704_ (.A(_10229_), .B(_10231_), .Y(_10232_));
XOR_g _16705_ (.A(_10229_), .B(_10231_), .Y(_10233_));
NAND_g _16706_ (.A(instr_jal), .B(_10233_), .Y(_10234_));
AND_g _16707_ (.A(_09973_), .B(_10219_), .Y(_10235_));
AND_g _16708_ (.A(_09973_), .B(_10220_), .Y(_10236_));
XNOR_g _16709_ (.A(_09974_), .B(_10220_), .Y(_10237_));
NAND_g _16710_ (.A(_08857_), .B(_10237_), .Y(_10238_));
AND_g _16711_ (.A(decoder_trigger), .B(_10238_), .Y(_10239_));
NAND_g _16712_ (.A(_10234_), .B(_10239_), .Y(_10240_));
NAND_g _16713_ (.A(_09974_), .B(_10112_), .Y(_10241_));
AND_g _16714_ (.A(_10240_), .B(_10241_), .Y(_10242_));
NOT_g _16715_ (.A(_10242_), .Y(_10243_));
NAND_g _16716_ (.A(_10227_), .B(_10243_), .Y(_00253_));
NAND_g _16717_ (.A(reg_next_pc[11]), .B(_09920_), .Y(_10244_));
AND_g _16718_ (.A(_10228_), .B(_10232_), .Y(_10245_));
NAND_g _16719_ (.A(decoded_imm_j[11]), .B(_09979_), .Y(_10246_));
NOR_g _16720_ (.A(decoded_imm_j[11]), .B(_09979_), .Y(_10247_));
XNOR_g _16721_ (.A(decoded_imm_j[11]), .B(_09980_), .Y(_10248_));
XNOR_g _16722_ (.A(_10245_), .B(_10248_), .Y(_10249_));
NAND_g _16723_ (.A(instr_jal), .B(_10249_), .Y(_10250_));
NOR_g _16724_ (.A(_09979_), .B(_10235_), .Y(_10251_));
AND_g _16725_ (.A(_09978_), .B(_10235_), .Y(_10252_));
AND_g _16726_ (.A(_09978_), .B(_10236_), .Y(_10253_));
NOR_g _16727_ (.A(_10251_), .B(_10253_), .Y(_10254_));
NAND_g _16728_ (.A(_08857_), .B(_10254_), .Y(_10255_));
AND_g _16729_ (.A(decoder_trigger), .B(_10255_), .Y(_10256_));
NAND_g _16730_ (.A(_10250_), .B(_10256_), .Y(_10257_));
NAND_g _16731_ (.A(_09980_), .B(_10112_), .Y(_10258_));
NAND_g _16732_ (.A(_10257_), .B(_10258_), .Y(_10259_));
NAND_g _16733_ (.A(_10244_), .B(_10259_), .Y(_00254_));
NAND_g _16734_ (.A(reg_next_pc[12]), .B(_09920_), .Y(_10260_));
NAND_g _16735_ (.A(decoded_imm_j[12]), .B(_09985_), .Y(_10261_));
XOR_g _16736_ (.A(decoded_imm_j[12]), .B(_09985_), .Y(_10262_));
AND_g _16737_ (.A(_10245_), .B(_10246_), .Y(_10263_));
NOR_g _16738_ (.A(_10247_), .B(_10263_), .Y(_10264_));
NAND_g _16739_ (.A(_10262_), .B(_10264_), .Y(_10265_));
XOR_g _16740_ (.A(_10262_), .B(_10264_), .Y(_10266_));
NAND_g _16741_ (.A(instr_jal), .B(_10266_), .Y(_10267_));
AND_g _16742_ (.A(_09985_), .B(_10252_), .Y(_10268_));
AND_g _16743_ (.A(_09985_), .B(_10253_), .Y(_10269_));
XNOR_g _16744_ (.A(_09986_), .B(_10253_), .Y(_10270_));
NAND_g _16745_ (.A(_08857_), .B(_10270_), .Y(_10271_));
AND_g _16746_ (.A(decoder_trigger), .B(_10271_), .Y(_10272_));
NAND_g _16747_ (.A(_10267_), .B(_10272_), .Y(_10273_));
NAND_g _16748_ (.A(_09986_), .B(_10112_), .Y(_10274_));
NAND_g _16749_ (.A(_10273_), .B(_10274_), .Y(_10275_));
NAND_g _16750_ (.A(_10260_), .B(_10275_), .Y(_00255_));
NAND_g _16751_ (.A(reg_next_pc[13]), .B(_09920_), .Y(_10276_));
AND_g _16752_ (.A(_10261_), .B(_10265_), .Y(_10277_));
NAND_g _16753_ (.A(decoded_imm_j[13]), .B(_09991_), .Y(_10278_));
NOR_g _16754_ (.A(decoded_imm_j[13]), .B(_09991_), .Y(_10279_));
XNOR_g _16755_ (.A(decoded_imm_j[13]), .B(_09992_), .Y(_10280_));
XNOR_g _16756_ (.A(_10277_), .B(_10280_), .Y(_10281_));
NAND_g _16757_ (.A(instr_jal), .B(_10281_), .Y(_10282_));
NOR_g _16758_ (.A(_09991_), .B(_10268_), .Y(_10283_));
AND_g _16759_ (.A(_09990_), .B(_10268_), .Y(_10284_));
AND_g _16760_ (.A(_09990_), .B(_10269_), .Y(_10285_));
NOR_g _16761_ (.A(_10283_), .B(_10285_), .Y(_10286_));
NAND_g _16762_ (.A(_08857_), .B(_10286_), .Y(_10287_));
AND_g _16763_ (.A(decoder_trigger), .B(_10287_), .Y(_10288_));
NAND_g _16764_ (.A(_10282_), .B(_10288_), .Y(_10289_));
NAND_g _16765_ (.A(_09992_), .B(_10112_), .Y(_10290_));
NAND_g _16766_ (.A(_10289_), .B(_10290_), .Y(_10291_));
NAND_g _16767_ (.A(_10276_), .B(_10291_), .Y(_00256_));
NAND_g _16768_ (.A(reg_next_pc[14]), .B(_09920_), .Y(_10292_));
NAND_g _16769_ (.A(decoded_imm_j[14]), .B(_09997_), .Y(_10293_));
XOR_g _16770_ (.A(decoded_imm_j[14]), .B(_09997_), .Y(_10294_));
AND_g _16771_ (.A(_10277_), .B(_10278_), .Y(_10295_));
NOR_g _16772_ (.A(_10279_), .B(_10295_), .Y(_10296_));
NAND_g _16773_ (.A(_10294_), .B(_10296_), .Y(_10297_));
XOR_g _16774_ (.A(_10294_), .B(_10296_), .Y(_10298_));
NAND_g _16775_ (.A(instr_jal), .B(_10298_), .Y(_10299_));
AND_g _16776_ (.A(_09997_), .B(_10284_), .Y(_10300_));
AND_g _16777_ (.A(_09997_), .B(_10285_), .Y(_10301_));
XNOR_g _16778_ (.A(_09998_), .B(_10285_), .Y(_10302_));
NAND_g _16779_ (.A(_08857_), .B(_10302_), .Y(_10303_));
AND_g _16780_ (.A(decoder_trigger), .B(_10303_), .Y(_10304_));
NAND_g _16781_ (.A(_10299_), .B(_10304_), .Y(_10305_));
NAND_g _16782_ (.A(_09998_), .B(_10112_), .Y(_10306_));
AND_g _16783_ (.A(_10305_), .B(_10306_), .Y(_10307_));
NOT_g _16784_ (.A(_10307_), .Y(_10308_));
NAND_g _16785_ (.A(_10292_), .B(_10308_), .Y(_00257_));
NAND_g _16786_ (.A(reg_next_pc[15]), .B(_09920_), .Y(_10309_));
AND_g _16787_ (.A(_10293_), .B(_10297_), .Y(_10310_));
NAND_g _16788_ (.A(decoded_imm_j[15]), .B(_10003_), .Y(_10311_));
NOR_g _16789_ (.A(decoded_imm_j[15]), .B(_10003_), .Y(_10312_));
XNOR_g _16790_ (.A(decoded_imm_j[15]), .B(_10004_), .Y(_10313_));
XNOR_g _16791_ (.A(_10310_), .B(_10313_), .Y(_10314_));
NAND_g _16792_ (.A(instr_jal), .B(_10314_), .Y(_10315_));
NOR_g _16793_ (.A(_10003_), .B(_10300_), .Y(_10316_));
AND_g _16794_ (.A(_10002_), .B(_10300_), .Y(_10317_));
AND_g _16795_ (.A(_10002_), .B(_10301_), .Y(_10318_));
NOR_g _16796_ (.A(_10316_), .B(_10318_), .Y(_10319_));
NAND_g _16797_ (.A(_08857_), .B(_10319_), .Y(_10320_));
AND_g _16798_ (.A(decoder_trigger), .B(_10320_), .Y(_10321_));
NAND_g _16799_ (.A(_10315_), .B(_10321_), .Y(_10322_));
NAND_g _16800_ (.A(_10004_), .B(_10112_), .Y(_10323_));
NAND_g _16801_ (.A(_10322_), .B(_10323_), .Y(_10324_));
NAND_g _16802_ (.A(_10309_), .B(_10324_), .Y(_00258_));
NAND_g _16803_ (.A(reg_next_pc[16]), .B(_09920_), .Y(_10325_));
NAND_g _16804_ (.A(decoded_imm_j[16]), .B(_10009_), .Y(_10326_));
XOR_g _16805_ (.A(decoded_imm_j[16]), .B(_10009_), .Y(_10327_));
AND_g _16806_ (.A(_10310_), .B(_10311_), .Y(_10328_));
NOR_g _16807_ (.A(_10312_), .B(_10328_), .Y(_10329_));
NAND_g _16808_ (.A(_10327_), .B(_10329_), .Y(_10330_));
XOR_g _16809_ (.A(_10327_), .B(_10329_), .Y(_10331_));
NAND_g _16810_ (.A(instr_jal), .B(_10331_), .Y(_10332_));
AND_g _16811_ (.A(_10009_), .B(_10317_), .Y(_10333_));
AND_g _16812_ (.A(_10009_), .B(_10318_), .Y(_10334_));
XNOR_g _16813_ (.A(_10010_), .B(_10318_), .Y(_10335_));
NAND_g _16814_ (.A(_08857_), .B(_10335_), .Y(_10336_));
AND_g _16815_ (.A(decoder_trigger), .B(_10336_), .Y(_10337_));
NAND_g _16816_ (.A(_10332_), .B(_10337_), .Y(_10338_));
NAND_g _16817_ (.A(_10010_), .B(_10112_), .Y(_10339_));
AND_g _16818_ (.A(_10338_), .B(_10339_), .Y(_10340_));
NOT_g _16819_ (.A(_10340_), .Y(_10341_));
NAND_g _16820_ (.A(_10325_), .B(_10341_), .Y(_00259_));
NAND_g _16821_ (.A(reg_next_pc[17]), .B(_09920_), .Y(_10342_));
AND_g _16822_ (.A(_10326_), .B(_10330_), .Y(_10343_));
NAND_g _16823_ (.A(decoded_imm_j[17]), .B(_10015_), .Y(_10344_));
NOR_g _16824_ (.A(decoded_imm_j[17]), .B(_10015_), .Y(_10345_));
XNOR_g _16825_ (.A(decoded_imm_j[17]), .B(_10016_), .Y(_10346_));
XNOR_g _16826_ (.A(_10343_), .B(_10346_), .Y(_10347_));
NAND_g _16827_ (.A(instr_jal), .B(_10347_), .Y(_10348_));
AND_g _16828_ (.A(_10014_), .B(_10333_), .Y(_10349_));
NOR_g _16829_ (.A(_10015_), .B(_10333_), .Y(_10350_));
AND_g _16830_ (.A(_10014_), .B(_10334_), .Y(_10351_));
NOR_g _16831_ (.A(_10350_), .B(_10351_), .Y(_10352_));
NAND_g _16832_ (.A(_08857_), .B(_10352_), .Y(_10353_));
AND_g _16833_ (.A(decoder_trigger), .B(_10353_), .Y(_10354_));
NAND_g _16834_ (.A(_10348_), .B(_10354_), .Y(_10355_));
NAND_g _16835_ (.A(_10016_), .B(_10112_), .Y(_10356_));
NAND_g _16836_ (.A(_10355_), .B(_10356_), .Y(_10357_));
NAND_g _16837_ (.A(_10342_), .B(_10357_), .Y(_00260_));
NAND_g _16838_ (.A(reg_next_pc[18]), .B(_09920_), .Y(_10358_));
NAND_g _16839_ (.A(decoded_imm_j[18]), .B(_10021_), .Y(_10359_));
XOR_g _16840_ (.A(decoded_imm_j[18]), .B(_10021_), .Y(_10360_));
AND_g _16841_ (.A(_10343_), .B(_10344_), .Y(_10361_));
NOR_g _16842_ (.A(_10345_), .B(_10361_), .Y(_10362_));
NAND_g _16843_ (.A(_10360_), .B(_10362_), .Y(_10363_));
XOR_g _16844_ (.A(_10360_), .B(_10362_), .Y(_10364_));
NAND_g _16845_ (.A(instr_jal), .B(_10364_), .Y(_10365_));
AND_g _16846_ (.A(_10021_), .B(_10349_), .Y(_10366_));
AND_g _16847_ (.A(_10021_), .B(_10351_), .Y(_10367_));
XNOR_g _16848_ (.A(_10022_), .B(_10351_), .Y(_10368_));
NAND_g _16849_ (.A(_08857_), .B(_10368_), .Y(_10369_));
AND_g _16850_ (.A(decoder_trigger), .B(_10369_), .Y(_10370_));
NAND_g _16851_ (.A(_10365_), .B(_10370_), .Y(_10371_));
NAND_g _16852_ (.A(_10022_), .B(_10112_), .Y(_10372_));
AND_g _16853_ (.A(_10371_), .B(_10372_), .Y(_10373_));
NOT_g _16854_ (.A(_10373_), .Y(_10374_));
NAND_g _16855_ (.A(_10358_), .B(_10374_), .Y(_00261_));
NAND_g _16856_ (.A(reg_next_pc[19]), .B(_09920_), .Y(_10375_));
AND_g _16857_ (.A(_10359_), .B(_10363_), .Y(_10376_));
NAND_g _16858_ (.A(decoded_imm_j[19]), .B(_10028_), .Y(_10377_));
NAND_g _16859_ (.A(_08945_), .B(_10027_), .Y(_10378_));
XNOR_g _16860_ (.A(decoded_imm_j[19]), .B(_10027_), .Y(_10379_));
XNOR_g _16861_ (.A(_10376_), .B(_10379_), .Y(_10380_));
NAND_g _16862_ (.A(instr_jal), .B(_10380_), .Y(_10381_));
NOR_g _16863_ (.A(_10028_), .B(_10366_), .Y(_10382_));
AND_g _16864_ (.A(_10026_), .B(_10366_), .Y(_10383_));
AND_g _16865_ (.A(_10026_), .B(_10367_), .Y(_10384_));
NOR_g _16866_ (.A(_10382_), .B(_10384_), .Y(_10385_));
NAND_g _16867_ (.A(_08857_), .B(_10385_), .Y(_10386_));
AND_g _16868_ (.A(decoder_trigger), .B(_10386_), .Y(_10387_));
NAND_g _16869_ (.A(_10381_), .B(_10387_), .Y(_10388_));
NAND_g _16870_ (.A(_10027_), .B(_10112_), .Y(_10389_));
NAND_g _16871_ (.A(_10388_), .B(_10389_), .Y(_10390_));
NAND_g _16872_ (.A(_10375_), .B(_10390_), .Y(_00262_));
NAND_g _16873_ (.A(reg_next_pc[20]), .B(_09920_), .Y(_10391_));
NAND_g _16874_ (.A(decoded_imm_j[31]), .B(_10033_), .Y(_10392_));
XNOR_g _16875_ (.A(_09017_), .B(_10033_), .Y(_10393_));
NAND_g _16876_ (.A(_10376_), .B(_10377_), .Y(_10394_));
NAND_g _16877_ (.A(_10378_), .B(_10394_), .Y(_10395_));
NOT_g _16878_ (.A(_10395_), .Y(_10396_));
NAND_g _16879_ (.A(_10393_), .B(_10396_), .Y(_10397_));
XNOR_g _16880_ (.A(_10393_), .B(_10395_), .Y(_10398_));
NAND_g _16881_ (.A(instr_jal), .B(_10398_), .Y(_10399_));
AND_g _16882_ (.A(_10033_), .B(_10383_), .Y(_10400_));
AND_g _16883_ (.A(_10033_), .B(_10384_), .Y(_10401_));
XNOR_g _16884_ (.A(_10034_), .B(_10384_), .Y(_10402_));
NAND_g _16885_ (.A(_08857_), .B(_10402_), .Y(_10403_));
AND_g _16886_ (.A(decoder_trigger), .B(_10403_), .Y(_10404_));
NAND_g _16887_ (.A(_10399_), .B(_10404_), .Y(_10405_));
NAND_g _16888_ (.A(_10034_), .B(_10112_), .Y(_10406_));
NAND_g _16889_ (.A(_10405_), .B(_10406_), .Y(_10407_));
NAND_g _16890_ (.A(_10391_), .B(_10407_), .Y(_00263_));
NAND_g _16891_ (.A(_10392_), .B(_10397_), .Y(_10408_));
NAND_g _16892_ (.A(decoded_imm_j[31]), .B(_10040_), .Y(_10409_));
XNOR_g _16893_ (.A(_09017_), .B(_10039_), .Y(_10410_));
XNOR_g _16894_ (.A(_10408_), .B(_10410_), .Y(_10411_));
NAND_g _16895_ (.A(instr_jal), .B(_10411_), .Y(_10412_));
NOR_g _16896_ (.A(_10040_), .B(_10400_), .Y(_10413_));
AND_g _16897_ (.A(_10038_), .B(_10400_), .Y(_10414_));
AND_g _16898_ (.A(_10038_), .B(_10401_), .Y(_10415_));
NOR_g _16899_ (.A(_10413_), .B(_10415_), .Y(_10416_));
NAND_g _16900_ (.A(_08857_), .B(_10416_), .Y(_10417_));
AND_g _16901_ (.A(decoder_trigger), .B(_10417_), .Y(_10418_));
NAND_g _16902_ (.A(_10412_), .B(_10418_), .Y(_10419_));
NAND_g _16903_ (.A(_10039_), .B(_10112_), .Y(_10420_));
NAND_g _16904_ (.A(_10419_), .B(_10420_), .Y(_10421_));
NAND_g _16905_ (.A(reg_next_pc[21]), .B(_09920_), .Y(_10422_));
NAND_g _16906_ (.A(_10421_), .B(_10422_), .Y(_00264_));
NAND_g _16907_ (.A(reg_next_pc[22]), .B(_09920_), .Y(_10423_));
NOR_g _16908_ (.A(_10397_), .B(_10410_), .Y(_10424_));
NOT_g _16909_ (.A(_10424_), .Y(_10425_));
AND_g _16910_ (.A(_10392_), .B(_10409_), .Y(_10426_));
NAND_g _16911_ (.A(_10425_), .B(_10426_), .Y(_10427_));
NAND_g _16912_ (.A(decoded_imm_j[31]), .B(_10045_), .Y(_10428_));
XNOR_g _16913_ (.A(_09017_), .B(_10045_), .Y(_10429_));
XNOR_g _16914_ (.A(decoded_imm_j[31]), .B(_10045_), .Y(_10430_));
NAND_g _16915_ (.A(_10427_), .B(_10429_), .Y(_10431_));
XNOR_g _16916_ (.A(_10427_), .B(_10430_), .Y(_10432_));
NAND_g _16917_ (.A(instr_jal), .B(_10432_), .Y(_10433_));
AND_g _16918_ (.A(_10045_), .B(_10414_), .Y(_10434_));
NAND_g _16919_ (.A(_10045_), .B(_10414_), .Y(_10435_));
XNOR_g _16920_ (.A(_10046_), .B(_10415_), .Y(_10436_));
NAND_g _16921_ (.A(_08857_), .B(_10436_), .Y(_10437_));
AND_g _16922_ (.A(decoder_trigger), .B(_10437_), .Y(_10438_));
NAND_g _16923_ (.A(_10433_), .B(_10438_), .Y(_10439_));
NAND_g _16924_ (.A(_10046_), .B(_10112_), .Y(_10440_));
AND_g _16925_ (.A(_10439_), .B(_10440_), .Y(_10441_));
NOT_g _16926_ (.A(_10441_), .Y(_10442_));
NAND_g _16927_ (.A(_10423_), .B(_10442_), .Y(_00265_));
NAND_g _16928_ (.A(reg_next_pc[23]), .B(_09920_), .Y(_10443_));
NAND_g _16929_ (.A(_10428_), .B(_10431_), .Y(_10444_));
NAND_g _16930_ (.A(decoded_imm_j[31]), .B(_10052_), .Y(_10445_));
XNOR_g _16931_ (.A(_09017_), .B(_10051_), .Y(_10446_));
XNOR_g _16932_ (.A(_10444_), .B(_10446_), .Y(_10447_));
NAND_g _16933_ (.A(instr_jal), .B(_10447_), .Y(_10448_));
NAND_g _16934_ (.A(_10051_), .B(_10435_), .Y(_10449_));
AND_g _16935_ (.A(_10050_), .B(_10434_), .Y(_10450_));
NOR_g _16936_ (.A(instr_jal), .B(_10450_), .Y(_10451_));
NAND_g _16937_ (.A(_10449_), .B(_10451_), .Y(_10452_));
AND_g _16938_ (.A(decoder_trigger), .B(_10452_), .Y(_10453_));
NAND_g _16939_ (.A(_10448_), .B(_10453_), .Y(_10454_));
NAND_g _16940_ (.A(_10051_), .B(_10112_), .Y(_10455_));
NAND_g _16941_ (.A(_10454_), .B(_10455_), .Y(_10456_));
NAND_g _16942_ (.A(_10443_), .B(_10456_), .Y(_00266_));
NAND_g _16943_ (.A(reg_next_pc[24]), .B(_09920_), .Y(_10457_));
NOR_g _16944_ (.A(_10430_), .B(_10446_), .Y(_10458_));
NAND_g _16945_ (.A(_10424_), .B(_10458_), .Y(_10459_));
AND_g _16946_ (.A(_10428_), .B(_10445_), .Y(_10460_));
AND_g _16947_ (.A(_10426_), .B(_10460_), .Y(_10461_));
AND_g _16948_ (.A(_10459_), .B(_10461_), .Y(_10462_));
AND_g _16949_ (.A(decoded_imm_j[31]), .B(_10057_), .Y(_10463_));
XNOR_g _16950_ (.A(decoded_imm_j[31]), .B(_10057_), .Y(_10464_));
NOR_g _16951_ (.A(_10462_), .B(_10464_), .Y(_10465_));
XOR_g _16952_ (.A(_10462_), .B(_10464_), .Y(_10466_));
NAND_g _16953_ (.A(instr_jal), .B(_10466_), .Y(_10467_));
NAND_g _16954_ (.A(_10057_), .B(_10450_), .Y(_10468_));
NOT_g _16955_ (.A(_10468_), .Y(_10469_));
NOR_g _16956_ (.A(_10057_), .B(_10450_), .Y(_10470_));
NOR_g _16957_ (.A(instr_jal), .B(_10470_), .Y(_10471_));
NAND_g _16958_ (.A(_10468_), .B(_10471_), .Y(_10472_));
AND_g _16959_ (.A(decoder_trigger), .B(_10472_), .Y(_10473_));
NAND_g _16960_ (.A(_10467_), .B(_10473_), .Y(_10474_));
NAND_g _16961_ (.A(_10058_), .B(_10112_), .Y(_10475_));
NAND_g _16962_ (.A(_10474_), .B(_10475_), .Y(_10476_));
NAND_g _16963_ (.A(_10457_), .B(_10476_), .Y(_00267_));
NOR_g _16964_ (.A(_10463_), .B(_10465_), .Y(_10477_));
NOR_g _16965_ (.A(_09017_), .B(_10063_), .Y(_10478_));
XNOR_g _16966_ (.A(decoded_imm_j[31]), .B(_10063_), .Y(_10479_));
XNOR_g _16967_ (.A(_10477_), .B(_10479_), .Y(_10480_));
NAND_g _16968_ (.A(instr_jal), .B(_10480_), .Y(_10481_));
NAND_g _16969_ (.A(_10063_), .B(_10468_), .Y(_10482_));
AND_g _16970_ (.A(_10062_), .B(_10469_), .Y(_10483_));
NOT_g _16971_ (.A(_10483_), .Y(_10484_));
NOR_g _16972_ (.A(instr_jal), .B(_10483_), .Y(_10485_));
NAND_g _16973_ (.A(_10482_), .B(_10485_), .Y(_10486_));
AND_g _16974_ (.A(decoder_trigger), .B(_10486_), .Y(_10487_));
NAND_g _16975_ (.A(_10481_), .B(_10487_), .Y(_10488_));
NAND_g _16976_ (.A(_10063_), .B(_10112_), .Y(_10489_));
NAND_g _16977_ (.A(_10488_), .B(_10489_), .Y(_10490_));
NAND_g _16978_ (.A(reg_next_pc[25]), .B(_09920_), .Y(_10491_));
NAND_g _16979_ (.A(_10490_), .B(_10491_), .Y(_00268_));
NAND_g _16980_ (.A(reg_next_pc[26]), .B(_09920_), .Y(_10492_));
NAND_g _16981_ (.A(_10465_), .B(_10479_), .Y(_10493_));
NOR_g _16982_ (.A(_10463_), .B(_10478_), .Y(_10494_));
NAND_g _16983_ (.A(_10493_), .B(_10494_), .Y(_10495_));
NAND_g _16984_ (.A(decoded_imm_j[31]), .B(_10068_), .Y(_10496_));
XNOR_g _16985_ (.A(_09017_), .B(_10068_), .Y(_10497_));
NOR_g _16986_ (.A(_10495_), .B(_10497_), .Y(_10498_));
NAND_g _16987_ (.A(_10495_), .B(_10497_), .Y(_10499_));
NAND_g _16988_ (.A(instr_jal), .B(_10499_), .Y(_10500_));
NOR_g _16989_ (.A(_10498_), .B(_10500_), .Y(_10501_));
NAND_g _16990_ (.A(_10069_), .B(_10484_), .Y(_10502_));
AND_g _16991_ (.A(_10068_), .B(_10483_), .Y(_10503_));
NOT_g _16992_ (.A(_10503_), .Y(_10504_));
NOR_g _16993_ (.A(instr_jal), .B(_10503_), .Y(_10505_));
NAND_g _16994_ (.A(_10502_), .B(_10505_), .Y(_10506_));
NAND_g _16995_ (.A(decoder_trigger), .B(_10506_), .Y(_10507_));
NOR_g _16996_ (.A(_10501_), .B(_10507_), .Y(_10508_));
NOR_g _16997_ (.A(_09893_), .B(_10068_), .Y(_10509_));
NOR_g _16998_ (.A(_10508_), .B(_10509_), .Y(_10510_));
NAND_g _16999_ (.A(resetn), .B(_10510_), .Y(_10511_));
NAND_g _17000_ (.A(_10492_), .B(_10511_), .Y(_00269_));
NAND_g _17001_ (.A(_10496_), .B(_10499_), .Y(_10512_));
XNOR_g _17002_ (.A(_09017_), .B(_10074_), .Y(_10513_));
XNOR_g _17003_ (.A(_10512_), .B(_10513_), .Y(_10514_));
NAND_g _17004_ (.A(instr_jal), .B(_10514_), .Y(_10515_));
NAND_g _17005_ (.A(_10073_), .B(_10503_), .Y(_10516_));
NAND_g _17006_ (.A(_10074_), .B(_10504_), .Y(_10517_));
AND_g _17007_ (.A(_08857_), .B(_10517_), .Y(_10518_));
NAND_g _17008_ (.A(_10516_), .B(_10518_), .Y(_10519_));
AND_g _17009_ (.A(decoder_trigger), .B(_10519_), .Y(_10520_));
NAND_g _17010_ (.A(_10515_), .B(_10520_), .Y(_10521_));
NAND_g _17011_ (.A(_10074_), .B(_10112_), .Y(_10522_));
NAND_g _17012_ (.A(_10521_), .B(_10522_), .Y(_10523_));
NAND_g _17013_ (.A(reg_next_pc[27]), .B(_09920_), .Y(_10524_));
NAND_g _17014_ (.A(_10523_), .B(_10524_), .Y(_00270_));
NAND_g _17015_ (.A(reg_next_pc[28]), .B(_09920_), .Y(_10525_));
AND_g _17016_ (.A(_10058_), .B(_10074_), .Y(_10526_));
AND_g _17017_ (.A(_10063_), .B(_10069_), .Y(_10527_));
NAND_g _17018_ (.A(_10526_), .B(_10527_), .Y(_10528_));
NAND_g _17019_ (.A(decoded_imm_j[31]), .B(_10528_), .Y(_10529_));
NOR_g _17020_ (.A(_10493_), .B(_10513_), .Y(_10530_));
NAND_g _17021_ (.A(_10497_), .B(_10530_), .Y(_10531_));
AND_g _17022_ (.A(_10529_), .B(_10531_), .Y(_10532_));
NAND_g _17023_ (.A(_10529_), .B(_10531_), .Y(_10533_));
NAND_g _17024_ (.A(decoded_imm_j[31]), .B(_10079_), .Y(_10534_));
XNOR_g _17025_ (.A(_09017_), .B(_10079_), .Y(_10535_));
XNOR_g _17026_ (.A(decoded_imm_j[31]), .B(_10079_), .Y(_10536_));
NAND_g _17027_ (.A(_10532_), .B(_10536_), .Y(_10537_));
NAND_g _17028_ (.A(_10533_), .B(_10535_), .Y(_10538_));
AND_g _17029_ (.A(instr_jal), .B(_10537_), .Y(_10539_));
NAND_g _17030_ (.A(_10538_), .B(_10539_), .Y(_10540_));
NOR_g _17031_ (.A(_10080_), .B(_10516_), .Y(_10541_));
NOT_g _17032_ (.A(_10541_), .Y(_10542_));
AND_g _17033_ (.A(_10080_), .B(_10516_), .Y(_10543_));
NOR_g _17034_ (.A(instr_jal), .B(_10543_), .Y(_10544_));
NAND_g _17035_ (.A(_10542_), .B(_10544_), .Y(_10545_));
AND_g _17036_ (.A(decoder_trigger), .B(_10545_), .Y(_10546_));
NAND_g _17037_ (.A(_10540_), .B(_10546_), .Y(_10547_));
NAND_g _17038_ (.A(_10080_), .B(_10112_), .Y(_10548_));
NAND_g _17039_ (.A(_10547_), .B(_10548_), .Y(_10549_));
NAND_g _17040_ (.A(_10525_), .B(_10549_), .Y(_00271_));
AND_g _17041_ (.A(decoded_imm_j[31]), .B(_10085_), .Y(_10550_));
XNOR_g _17042_ (.A(decoded_imm_j[31]), .B(_10085_), .Y(_10551_));
NAND_g _17043_ (.A(_10534_), .B(_10538_), .Y(_10552_));
NAND_g _17044_ (.A(_10534_), .B(_10551_), .Y(_10553_));
XNOR_g _17045_ (.A(_10551_), .B(_10552_), .Y(_10554_));
NAND_g _17046_ (.A(instr_jal), .B(_10554_), .Y(_10555_));
NAND_g _17047_ (.A(_10084_), .B(_10541_), .Y(_10556_));
NOR_g _17048_ (.A(_10085_), .B(_10541_), .Y(_10557_));
NOR_g _17049_ (.A(instr_jal), .B(_10557_), .Y(_10558_));
NAND_g _17050_ (.A(_10556_), .B(_10558_), .Y(_10559_));
AND_g _17051_ (.A(decoder_trigger), .B(_10559_), .Y(_10560_));
NAND_g _17052_ (.A(_10555_), .B(_10560_), .Y(_10561_));
NAND_g _17053_ (.A(_10086_), .B(_10112_), .Y(_10562_));
NAND_g _17054_ (.A(_10561_), .B(_10562_), .Y(_10563_));
NAND_g _17055_ (.A(reg_next_pc[29]), .B(_09920_), .Y(_10564_));
NAND_g _17056_ (.A(_10563_), .B(_10564_), .Y(_00272_));
NAND_g _17057_ (.A(reg_next_pc[30]), .B(_09920_), .Y(_10565_));
NOR_g _17058_ (.A(_10091_), .B(_10556_), .Y(_10566_));
NOT_g _17059_ (.A(_10566_), .Y(_10567_));
NAND_g _17060_ (.A(_08857_), .B(_10567_), .Y(_10568_));
AND_g _17061_ (.A(decoder_trigger), .B(_10568_), .Y(_10569_));
NAND_g _17062_ (.A(decoder_trigger), .B(_10568_), .Y(_10570_));
AND_g _17063_ (.A(decoder_trigger), .B(_10091_), .Y(_10571_));
NAND_g _17064_ (.A(_10556_), .B(_10571_), .Y(_10572_));
NAND_g _17065_ (.A(_10570_), .B(_10572_), .Y(_10573_));
AND_g _17066_ (.A(decoded_imm_j[31]), .B(_10091_), .Y(_10574_));
NOR_g _17067_ (.A(decoded_imm_j[31]), .B(_10091_), .Y(_10575_));
XNOR_g _17068_ (.A(decoded_imm_j[31]), .B(_10091_), .Y(_10576_));
AND_g _17069_ (.A(_10552_), .B(_10553_), .Y(_10577_));
NOR_g _17070_ (.A(_10550_), .B(_10577_), .Y(_10578_));
XNOR_g _17071_ (.A(_10576_), .B(_10578_), .Y(_10579_));
NAND_g _17072_ (.A(instr_jal), .B(_10579_), .Y(_10580_));
NAND_g _17073_ (.A(_10573_), .B(_10580_), .Y(_10581_));
NAND_g _17074_ (.A(_10091_), .B(_10112_), .Y(_10582_));
NAND_g _17075_ (.A(_10581_), .B(_10582_), .Y(_10583_));
NAND_g _17076_ (.A(_10565_), .B(_10583_), .Y(_00273_));
NAND_g _17077_ (.A(_10574_), .B(_10578_), .Y(_10584_));
NAND_g _17078_ (.A(_10575_), .B(_10577_), .Y(_10585_));
AND_g _17079_ (.A(instr_jal), .B(_10585_), .Y(_10586_));
NAND_g _17080_ (.A(_10584_), .B(_10586_), .Y(_10587_));
NAND_g _17081_ (.A(_10569_), .B(_10587_), .Y(_10588_));
XNOR_g _17082_ (.A(_10095_), .B(_10588_), .Y(_10589_));
NAND_g _17083_ (.A(_09075_), .B(_10589_), .Y(_10590_));
NAND_g _17084_ (.A(reg_next_pc[31]), .B(_09920_), .Y(_10591_));
NAND_g _17085_ (.A(_10590_), .B(_10591_), .Y(_00274_));
NOR_g _17086_ (.A(cpu_state[6]), .B(cpu_state[7]), .Y(_10592_));
AND_g _17087_ (.A(cpu_state[5]), .B(_09020_), .Y(_10593_));
AND_g _17088_ (.A(_10592_), .B(_10593_), .Y(_10594_));
AND_g _17089_ (.A(_09069_), .B(_10594_), .Y(_10595_));
NAND_g _17090_ (.A(_09069_), .B(_10594_), .Y(_10596_));
NOR_g _17091_ (.A(cpu_state[5]), .B(_09020_), .Y(_10597_));
AND_g _17092_ (.A(_10592_), .B(_10597_), .Y(_10598_));
AND_g _17093_ (.A(_09069_), .B(_10598_), .Y(_10599_));
NAND_g _17094_ (.A(_09069_), .B(_10598_), .Y(_10600_));
AND_g _17095_ (.A(_10596_), .B(_10600_), .Y(_10601_));
NAND_g _17096_ (.A(_10596_), .B(_10600_), .Y(_10602_));
AND_g _17097_ (.A(resetn), .B(_10602_), .Y(_10603_));
NAND_g _17098_ (.A(resetn), .B(_10602_), .Y(_10604_));
NOR_g _17099_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi), .B(is_lui_auipc_jal), .Y(_10605_));
NOR_g _17100_ (.A(_10596_), .B(_10605_), .Y(_10606_));
NAND_g _17101_ (.A(decoded_imm[0]), .B(_10606_), .Y(_10607_));
NOR_g _17102_ (.A(decoded_imm_j[11]), .B(decoded_imm_j[1]), .Y(_10608_));
NOR_g _17103_ (.A(decoded_imm_j[2]), .B(decoded_imm_j[3]), .Y(_10609_));
AND_g _17104_ (.A(_08879_), .B(_10609_), .Y(_10610_));
NAND_g _17105_ (.A(_10608_), .B(_10610_), .Y(_10611_));
NAND_g _17106_ (.A(cpuregs[24][0]), .B(_09027_), .Y(_10612_));
NAND_g _17107_ (.A(cpuregs[28][0]), .B(_00007_[2]), .Y(_10613_));
AND_g _17108_ (.A(_09025_), .B(_10613_), .Y(_10614_));
NAND_g _17109_ (.A(_10612_), .B(_10614_), .Y(_10615_));
NAND_g _17110_ (.A(cpuregs[25][0]), .B(_09027_), .Y(_10616_));
NAND_g _17111_ (.A(cpuregs[29][0]), .B(_00007_[2]), .Y(_10617_));
AND_g _17112_ (.A(_00007_[0]), .B(_10617_), .Y(_10618_));
NAND_g _17113_ (.A(_10616_), .B(_10618_), .Y(_10619_));
NAND_g _17114_ (.A(_10615_), .B(_10619_), .Y(_10620_));
NAND_g _17115_ (.A(_09026_), .B(_10620_), .Y(_10621_));
NAND_g _17116_ (.A(cpuregs[26][0]), .B(_09027_), .Y(_10622_));
NAND_g _17117_ (.A(cpuregs[30][0]), .B(_00007_[2]), .Y(_10623_));
AND_g _17118_ (.A(_09025_), .B(_10623_), .Y(_10624_));
NAND_g _17119_ (.A(_10622_), .B(_10624_), .Y(_10625_));
NAND_g _17120_ (.A(cpuregs[31][0]), .B(_00007_[2]), .Y(_10626_));
NAND_g _17121_ (.A(cpuregs[27][0]), .B(_09027_), .Y(_10627_));
AND_g _17122_ (.A(_00007_[0]), .B(_10627_), .Y(_10628_));
NAND_g _17123_ (.A(_10626_), .B(_10628_), .Y(_10629_));
NAND_g _17124_ (.A(_10625_), .B(_10629_), .Y(_10630_));
NAND_g _17125_ (.A(_00007_[1]), .B(_10630_), .Y(_10631_));
AND_g _17126_ (.A(_00007_[3]), .B(_10621_), .Y(_10632_));
NAND_g _17127_ (.A(_10631_), .B(_10632_), .Y(_10633_));
NAND_g _17128_ (.A(cpuregs[20][0]), .B(_00007_[2]), .Y(_10634_));
NAND_g _17129_ (.A(cpuregs[16][0]), .B(_09027_), .Y(_10635_));
AND_g _17130_ (.A(_10634_), .B(_10635_), .Y(_10636_));
NAND_g _17131_ (.A(_09025_), .B(_10636_), .Y(_10637_));
NAND_g _17132_ (.A(cpuregs[21][0]), .B(_00007_[2]), .Y(_10638_));
NAND_g _17133_ (.A(cpuregs[17][0]), .B(_09027_), .Y(_10639_));
AND_g _17134_ (.A(_00007_[0]), .B(_10639_), .Y(_10640_));
NAND_g _17135_ (.A(_10638_), .B(_10640_), .Y(_10641_));
AND_g _17136_ (.A(_09026_), .B(_10641_), .Y(_10642_));
NAND_g _17137_ (.A(_10637_), .B(_10642_), .Y(_10643_));
NAND_g _17138_ (.A(cpuregs[23][0]), .B(_00007_[2]), .Y(_10644_));
NAND_g _17139_ (.A(cpuregs[19][0]), .B(_09027_), .Y(_10645_));
AND_g _17140_ (.A(_00007_[0]), .B(_10645_), .Y(_10646_));
NAND_g _17141_ (.A(_10644_), .B(_10646_), .Y(_10647_));
NAND_g _17142_ (.A(cpuregs[22][0]), .B(_00007_[2]), .Y(_10648_));
NAND_g _17143_ (.A(cpuregs[18][0]), .B(_09027_), .Y(_10649_));
AND_g _17144_ (.A(_10648_), .B(_10649_), .Y(_10650_));
NAND_g _17145_ (.A(_09025_), .B(_10650_), .Y(_10651_));
AND_g _17146_ (.A(_00007_[1]), .B(_10651_), .Y(_10652_));
NAND_g _17147_ (.A(_10647_), .B(_10652_), .Y(_10653_));
NAND_g _17148_ (.A(_10643_), .B(_10653_), .Y(_10654_));
NAND_g _17149_ (.A(_09028_), .B(_10654_), .Y(_10655_));
AND_g _17150_ (.A(_10633_), .B(_10655_), .Y(_10656_));
NAND_g _17151_ (.A(cpuregs[13][0]), .B(_09026_), .Y(_10657_));
NAND_g _17152_ (.A(cpuregs[15][0]), .B(_00007_[1]), .Y(_10658_));
AND_g _17153_ (.A(_00007_[2]), .B(_10658_), .Y(_10659_));
NAND_g _17154_ (.A(_10657_), .B(_10659_), .Y(_10660_));
NAND_g _17155_ (.A(cpuregs[9][0]), .B(_09026_), .Y(_10661_));
NAND_g _17156_ (.A(cpuregs[11][0]), .B(_00007_[1]), .Y(_10662_));
AND_g _17157_ (.A(_09027_), .B(_10662_), .Y(_10663_));
NAND_g _17158_ (.A(_10661_), .B(_10663_), .Y(_10664_));
AND_g _17159_ (.A(_00007_[0]), .B(_10664_), .Y(_10665_));
NAND_g _17160_ (.A(_10660_), .B(_10665_), .Y(_10666_));
NAND_g _17161_ (.A(cpuregs[12][0]), .B(_09026_), .Y(_10667_));
NAND_g _17162_ (.A(cpuregs[14][0]), .B(_00007_[1]), .Y(_10668_));
AND_g _17163_ (.A(_00007_[2]), .B(_10668_), .Y(_10669_));
NAND_g _17164_ (.A(_10667_), .B(_10669_), .Y(_10670_));
NAND_g _17165_ (.A(cpuregs[8][0]), .B(_09026_), .Y(_10671_));
NAND_g _17166_ (.A(cpuregs[10][0]), .B(_00007_[1]), .Y(_10672_));
AND_g _17167_ (.A(_09027_), .B(_10672_), .Y(_10673_));
NAND_g _17168_ (.A(_10671_), .B(_10673_), .Y(_10674_));
AND_g _17169_ (.A(_09025_), .B(_10674_), .Y(_10675_));
NAND_g _17170_ (.A(_10670_), .B(_10675_), .Y(_10676_));
NAND_g _17171_ (.A(_10666_), .B(_10676_), .Y(_10677_));
NAND_g _17172_ (.A(_00007_[3]), .B(_10677_), .Y(_10678_));
NAND_g _17173_ (.A(_09003_), .B(_00007_[2]), .Y(_10679_));
NOR_g _17174_ (.A(cpuregs[2][0]), .B(_00007_[2]), .Y(_10680_));
NOR_g _17175_ (.A(_00007_[0]), .B(_10680_), .Y(_10681_));
NAND_g _17176_ (.A(_10679_), .B(_10681_), .Y(_10682_));
NAND_g _17177_ (.A(_08963_), .B(_00007_[2]), .Y(_10683_));
NOR_g _17178_ (.A(cpuregs[3][0]), .B(_00007_[2]), .Y(_10684_));
NOR_g _17179_ (.A(_09025_), .B(_10684_), .Y(_10685_));
NAND_g _17180_ (.A(_10683_), .B(_10685_), .Y(_10686_));
AND_g _17181_ (.A(_10682_), .B(_10686_), .Y(_10687_));
NAND_g _17182_ (.A(_08904_), .B(_00007_[2]), .Y(_10688_));
NOR_g _17183_ (.A(cpuregs[0][0]), .B(_00007_[2]), .Y(_10689_));
NOR_g _17184_ (.A(_00007_[0]), .B(_10689_), .Y(_10690_));
NAND_g _17185_ (.A(_10688_), .B(_10690_), .Y(_10691_));
NAND_g _17186_ (.A(_08946_), .B(_00007_[2]), .Y(_10692_));
NOR_g _17187_ (.A(cpuregs[1][0]), .B(_00007_[2]), .Y(_10693_));
NOR_g _17188_ (.A(_09025_), .B(_10693_), .Y(_10694_));
NAND_g _17189_ (.A(_10692_), .B(_10694_), .Y(_10695_));
AND_g _17190_ (.A(_10691_), .B(_10695_), .Y(_10696_));
NAND_g _17191_ (.A(_00007_[1]), .B(_10687_), .Y(_10697_));
NAND_g _17192_ (.A(_09026_), .B(_10696_), .Y(_10698_));
AND_g _17193_ (.A(_10697_), .B(_10698_), .Y(_10699_));
NAND_g _17194_ (.A(_09028_), .B(_10699_), .Y(_10700_));
AND_g _17195_ (.A(_10678_), .B(_10700_), .Y(_10701_));
NAND_g _17196_ (.A(_00007_[4]), .B(_10656_), .Y(_10702_));
NAND_g _17197_ (.A(_09029_), .B(_10701_), .Y(_10703_));
AND_g _17198_ (.A(_10611_), .B(_10703_), .Y(_10704_));
AND_g _17199_ (.A(_10702_), .B(_10704_), .Y(_10705_));
NAND_g _17200_ (.A(_10599_), .B(_10705_), .Y(_10706_));
NOR_g _17201_ (.A(instr_rdcycle), .B(instr_rdcycleh), .Y(_10707_));
NOR_g _17202_ (.A(instr_rdinstr), .B(instr_rdinstrh), .Y(_10708_));
AND_g _17203_ (.A(_10707_), .B(_10708_), .Y(_10709_));
NOT_g _17204_ (.A(_10709_), .Y(_10710_));
NOR_g _17205_ (.A(instr_lb), .B(instr_sb), .Y(_10711_));
AND_g _17206_ (.A(_08859_), .B(_10711_), .Y(_10712_));
NOR_g _17207_ (.A(instr_bge), .B(instr_blt), .Y(_10713_));
NOR_g _17208_ (.A(instr_bne), .B(instr_beq), .Y(_10714_));
AND_g _17209_ (.A(_10713_), .B(_10714_), .Y(_10715_));
AND_g _17210_ (.A(_10712_), .B(_10715_), .Y(_10716_));
NOR_g _17211_ (.A(instr_slt), .B(instr_slti), .Y(_10717_));
NOR_g _17212_ (.A(instr_sltu), .B(instr_sltiu), .Y(_10718_));
AND_g _17213_ (.A(_10717_), .B(_10718_), .Y(_10719_));
AND_g _17214_ (.A(_10709_), .B(_10719_), .Y(_10720_));
AND_g _17215_ (.A(_10716_), .B(_10720_), .Y(_10721_));
NOR_g _17216_ (.A(instr_lw), .B(instr_lbu), .Y(_10722_));
NOR_g _17217_ (.A(instr_sra), .B(instr_srl), .Y(_10723_));
AND_g _17218_ (.A(_10722_), .B(_10723_), .Y(_10724_));
NOR_g _17219_ (.A(instr_sub), .B(instr_add), .Y(_10725_));
NOR_g _17220_ (.A(instr_sw), .B(instr_sh), .Y(_10726_));
AND_g _17221_ (.A(_10725_), .B(_10726_), .Y(_10727_));
AND_g _17222_ (.A(_10724_), .B(_10727_), .Y(_10728_));
NOR_g _17223_ (.A(instr_ori), .B(instr_addi), .Y(_10729_));
NOR_g _17224_ (.A(instr_bgeu), .B(instr_bltu), .Y(_10730_));
AND_g _17225_ (.A(_10729_), .B(_10730_), .Y(_10731_));
NOR_g _17226_ (.A(instr_and), .B(instr_or), .Y(_10732_));
NOR_g _17227_ (.A(instr_sll), .B(instr_andi), .Y(_10733_));
AND_g _17228_ (.A(_10732_), .B(_10733_), .Y(_10734_));
AND_g _17229_ (.A(_10731_), .B(_10734_), .Y(_10735_));
AND_g _17230_ (.A(_10728_), .B(_10735_), .Y(_10736_));
NOR_g _17231_ (.A(instr_lui), .B(instr_auipc), .Y(_10737_));
NAND_g _17232_ (.A(_08855_), .B(_08856_), .Y(_10738_));
NAND_g _17233_ (.A(_08857_), .B(_10737_), .Y(_00002_));
NOR_g _17234_ (.A(instr_jalr), .B(_00002_), .Y(_10739_));
NOR_g _17235_ (.A(instr_lh), .B(instr_lhu), .Y(_10740_));
NOR_g _17236_ (.A(instr_srli), .B(instr_srai), .Y(_10741_));
NOR_g _17237_ (.A(instr_xor), .B(instr_xori), .Y(_10742_));
NAND_g _17238_ (.A(_08792_), .B(_08795_), .Y(_10743_));
AND_g _17239_ (.A(_10741_), .B(_10742_), .Y(_10744_));
AND_g _17240_ (.A(_10740_), .B(_10744_), .Y(_10745_));
AND_g _17241_ (.A(_10739_), .B(_10745_), .Y(_10746_));
AND_g _17242_ (.A(_10736_), .B(_10746_), .Y(_10747_));
NAND_g _17243_ (.A(_10721_), .B(_10747_), .Y(_10748_));
NOT_g _17244_ (.A(_10748_), .Y(_10749_));
AND_g _17245_ (.A(_10709_), .B(_10748_), .Y(_10750_));
NAND_g _17246_ (.A(_08861_), .B(_10750_), .Y(_10751_));
NOR_g _17247_ (.A(is_lb_lh_lw_lbu_lhu), .B(_10751_), .Y(_10752_));
AND_g _17248_ (.A(_10595_), .B(_10752_), .Y(_10753_));
AND_g _17249_ (.A(_10605_), .B(_10753_), .Y(_10754_));
NOT_g _17250_ (.A(_10754_), .Y(_10755_));
NAND_g _17251_ (.A(_10705_), .B(_10754_), .Y(_10756_));
AND_g _17252_ (.A(_10706_), .B(_10756_), .Y(_10757_));
NAND_g _17253_ (.A(_10607_), .B(_10757_), .Y(_10758_));
NAND_g _17254_ (.A(_10603_), .B(_10758_), .Y(_10759_));
NAND_g _17255_ (.A(pcpi_rs2[0]), .B(_10604_), .Y(_10760_));
NAND_g _17256_ (.A(_10759_), .B(_10760_), .Y(_00275_));
NAND_g _17257_ (.A(decoded_imm[1]), .B(_10606_), .Y(_10761_));
NOR_g _17258_ (.A(cpuregs[16][1]), .B(_00007_[2]), .Y(_10762_));
NOR_g _17259_ (.A(cpuregs[20][1]), .B(_09027_), .Y(_10763_));
NOR_g _17260_ (.A(_10762_), .B(_10763_), .Y(_10764_));
NOR_g _17261_ (.A(cpuregs[18][1]), .B(_00007_[2]), .Y(_10765_));
NOR_g _17262_ (.A(cpuregs[22][1]), .B(_09027_), .Y(_10766_));
NOR_g _17263_ (.A(_10765_), .B(_10766_), .Y(_10767_));
NOR_g _17264_ (.A(cpuregs[17][1]), .B(_00007_[2]), .Y(_10768_));
NAND_g _17265_ (.A(_08982_), .B(_00007_[2]), .Y(_10769_));
NAND_g _17266_ (.A(_08885_), .B(_00007_[2]), .Y(_10770_));
NOR_g _17267_ (.A(cpuregs[19][1]), .B(_00007_[2]), .Y(_10771_));
NOR_g _17268_ (.A(_09025_), .B(_10771_), .Y(_10772_));
NAND_g _17269_ (.A(_10770_), .B(_10772_), .Y(_10773_));
NAND_g _17270_ (.A(_09025_), .B(_10767_), .Y(_10774_));
AND_g _17271_ (.A(_10773_), .B(_10774_), .Y(_10775_));
NAND_g _17272_ (.A(_00007_[1]), .B(_10775_), .Y(_10776_));
NOR_g _17273_ (.A(_09025_), .B(_10768_), .Y(_10777_));
NAND_g _17274_ (.A(_10769_), .B(_10777_), .Y(_10778_));
NAND_g _17275_ (.A(_09025_), .B(_10764_), .Y(_10779_));
AND_g _17276_ (.A(_10778_), .B(_10779_), .Y(_10780_));
NAND_g _17277_ (.A(_09026_), .B(_10780_), .Y(_10781_));
AND_g _17278_ (.A(_10776_), .B(_10781_), .Y(_10782_));
NAND_g _17279_ (.A(_09028_), .B(_10782_), .Y(_10783_));
NAND_g _17280_ (.A(cpuregs[27][1]), .B(_00007_[1]), .Y(_10784_));
NAND_g _17281_ (.A(cpuregs[25][1]), .B(_09026_), .Y(_10785_));
NAND_g _17282_ (.A(_10784_), .B(_10785_), .Y(_10786_));
NAND_g _17283_ (.A(_09027_), .B(_10786_), .Y(_10787_));
NAND_g _17284_ (.A(cpuregs[31][1]), .B(_00007_[1]), .Y(_10788_));
NAND_g _17285_ (.A(cpuregs[29][1]), .B(_09026_), .Y(_10789_));
NAND_g _17286_ (.A(_10788_), .B(_10789_), .Y(_10790_));
NAND_g _17287_ (.A(_00007_[2]), .B(_10790_), .Y(_10791_));
AND_g _17288_ (.A(_00007_[0]), .B(_10791_), .Y(_10792_));
NAND_g _17289_ (.A(_10787_), .B(_10792_), .Y(_10793_));
NAND_g _17290_ (.A(cpuregs[26][1]), .B(_00007_[1]), .Y(_10794_));
NAND_g _17291_ (.A(cpuregs[24][1]), .B(_09026_), .Y(_10795_));
NAND_g _17292_ (.A(_10794_), .B(_10795_), .Y(_10796_));
NAND_g _17293_ (.A(_09027_), .B(_10796_), .Y(_10797_));
NAND_g _17294_ (.A(cpuregs[30][1]), .B(_00007_[1]), .Y(_10798_));
NAND_g _17295_ (.A(cpuregs[28][1]), .B(_09026_), .Y(_10799_));
NAND_g _17296_ (.A(_10798_), .B(_10799_), .Y(_10800_));
NAND_g _17297_ (.A(_00007_[2]), .B(_10800_), .Y(_10801_));
AND_g _17298_ (.A(_09025_), .B(_10801_), .Y(_10802_));
NAND_g _17299_ (.A(_10797_), .B(_10802_), .Y(_10803_));
AND_g _17300_ (.A(_00007_[3]), .B(_10803_), .Y(_10804_));
NAND_g _17301_ (.A(_10793_), .B(_10804_), .Y(_10805_));
AND_g _17302_ (.A(_10783_), .B(_10805_), .Y(_10806_));
NAND_g _17303_ (.A(cpuregs[1][1]), .B(_09027_), .Y(_10807_));
NAND_g _17304_ (.A(cpuregs[5][1]), .B(_00007_[2]), .Y(_10808_));
AND_g _17305_ (.A(_00007_[0]), .B(_10808_), .Y(_10809_));
NAND_g _17306_ (.A(_10807_), .B(_10809_), .Y(_10810_));
NAND_g _17307_ (.A(cpuregs[0][1]), .B(_09027_), .Y(_10811_));
NAND_g _17308_ (.A(cpuregs[4][1]), .B(_00007_[2]), .Y(_10812_));
AND_g _17309_ (.A(_09025_), .B(_10812_), .Y(_10813_));
NAND_g _17310_ (.A(_10811_), .B(_10813_), .Y(_10814_));
AND_g _17311_ (.A(_09026_), .B(_10814_), .Y(_10815_));
NAND_g _17312_ (.A(_10810_), .B(_10815_), .Y(_10816_));
NAND_g _17313_ (.A(cpuregs[3][1]), .B(_09027_), .Y(_10817_));
NAND_g _17314_ (.A(cpuregs[7][1]), .B(_00007_[2]), .Y(_10818_));
AND_g _17315_ (.A(_00007_[0]), .B(_10818_), .Y(_10819_));
NAND_g _17316_ (.A(_10817_), .B(_10819_), .Y(_10820_));
NAND_g _17317_ (.A(cpuregs[2][1]), .B(_09027_), .Y(_10821_));
NAND_g _17318_ (.A(cpuregs[6][1]), .B(_00007_[2]), .Y(_10822_));
AND_g _17319_ (.A(_09025_), .B(_10822_), .Y(_10823_));
NAND_g _17320_ (.A(_10821_), .B(_10823_), .Y(_10824_));
AND_g _17321_ (.A(_00007_[1]), .B(_10824_), .Y(_10825_));
NAND_g _17322_ (.A(_10820_), .B(_10825_), .Y(_10826_));
NAND_g _17323_ (.A(_10816_), .B(_10826_), .Y(_10827_));
NAND_g _17324_ (.A(_09028_), .B(_10827_), .Y(_10828_));
NAND_g _17325_ (.A(cpuregs[14][1]), .B(_09025_), .Y(_10829_));
NAND_g _17326_ (.A(cpuregs[15][1]), .B(_00007_[0]), .Y(_10830_));
NAND_g _17327_ (.A(_10829_), .B(_10830_), .Y(_10831_));
NAND_g _17328_ (.A(_00007_[2]), .B(_10831_), .Y(_10832_));
NAND_g _17329_ (.A(cpuregs[10][1]), .B(_09025_), .Y(_10833_));
NAND_g _17330_ (.A(cpuregs[11][1]), .B(_00007_[0]), .Y(_10834_));
NAND_g _17331_ (.A(_10833_), .B(_10834_), .Y(_10835_));
NAND_g _17332_ (.A(_09027_), .B(_10835_), .Y(_10836_));
AND_g _17333_ (.A(_10832_), .B(_10836_), .Y(_10837_));
NAND_g _17334_ (.A(cpuregs[12][1]), .B(_09025_), .Y(_10838_));
NAND_g _17335_ (.A(cpuregs[13][1]), .B(_00007_[0]), .Y(_10839_));
NAND_g _17336_ (.A(_10838_), .B(_10839_), .Y(_10840_));
NAND_g _17337_ (.A(_00007_[2]), .B(_10840_), .Y(_10841_));
NAND_g _17338_ (.A(cpuregs[8][1]), .B(_09025_), .Y(_10842_));
NAND_g _17339_ (.A(cpuregs[9][1]), .B(_00007_[0]), .Y(_10843_));
NAND_g _17340_ (.A(_10842_), .B(_10843_), .Y(_10844_));
NAND_g _17341_ (.A(_09027_), .B(_10844_), .Y(_10845_));
AND_g _17342_ (.A(_10841_), .B(_10845_), .Y(_10846_));
NAND_g _17343_ (.A(_09026_), .B(_10846_), .Y(_10847_));
NAND_g _17344_ (.A(_00007_[1]), .B(_10837_), .Y(_10848_));
AND_g _17345_ (.A(_00007_[3]), .B(_10847_), .Y(_10849_));
NAND_g _17346_ (.A(_10848_), .B(_10849_), .Y(_10850_));
NAND_g _17347_ (.A(_00007_[4]), .B(_10806_), .Y(_10851_));
AND_g _17348_ (.A(_09029_), .B(_10828_), .Y(_10852_));
NAND_g _17349_ (.A(_10850_), .B(_10852_), .Y(_10853_));
AND_g _17350_ (.A(_10611_), .B(_10853_), .Y(_10854_));
AND_g _17351_ (.A(_10851_), .B(_10854_), .Y(_10855_));
NAND_g _17352_ (.A(_10599_), .B(_10855_), .Y(_10856_));
NAND_g _17353_ (.A(_10754_), .B(_10855_), .Y(_10857_));
AND_g _17354_ (.A(_10856_), .B(_10857_), .Y(_10858_));
AND_g _17355_ (.A(_10761_), .B(_10858_), .Y(_10859_));
NAND_g _17356_ (.A(_08812_), .B(_10604_), .Y(_10860_));
NAND_g _17357_ (.A(_10603_), .B(_10859_), .Y(_10861_));
AND_g _17358_ (.A(_10860_), .B(_10861_), .Y(_00276_));
NAND_g _17359_ (.A(decoded_imm[2]), .B(_10606_), .Y(_10862_));
NAND_g _17360_ (.A(cpuregs[19][2]), .B(_09027_), .Y(_10863_));
NAND_g _17361_ (.A(cpuregs[23][2]), .B(_00007_[2]), .Y(_10864_));
AND_g _17362_ (.A(_00007_[0]), .B(_10864_), .Y(_10865_));
NAND_g _17363_ (.A(_10863_), .B(_10865_), .Y(_10866_));
NAND_g _17364_ (.A(cpuregs[18][2]), .B(_09027_), .Y(_10867_));
NAND_g _17365_ (.A(cpuregs[22][2]), .B(_00007_[2]), .Y(_10868_));
AND_g _17366_ (.A(_09025_), .B(_10868_), .Y(_10869_));
NAND_g _17367_ (.A(_10867_), .B(_10869_), .Y(_10870_));
AND_g _17368_ (.A(_09028_), .B(_10870_), .Y(_10871_));
NAND_g _17369_ (.A(_10866_), .B(_10871_), .Y(_10872_));
NAND_g _17370_ (.A(cpuregs[27][2]), .B(_09027_), .Y(_10873_));
NAND_g _17371_ (.A(cpuregs[31][2]), .B(_00007_[2]), .Y(_10874_));
AND_g _17372_ (.A(_00007_[0]), .B(_10874_), .Y(_10875_));
NAND_g _17373_ (.A(_10873_), .B(_10875_), .Y(_10876_));
NAND_g _17374_ (.A(cpuregs[26][2]), .B(_09027_), .Y(_10877_));
NAND_g _17375_ (.A(cpuregs[30][2]), .B(_00007_[2]), .Y(_10878_));
AND_g _17376_ (.A(_09025_), .B(_10878_), .Y(_10879_));
NAND_g _17377_ (.A(_10877_), .B(_10879_), .Y(_10880_));
AND_g _17378_ (.A(_00007_[3]), .B(_10880_), .Y(_10881_));
NAND_g _17379_ (.A(_10876_), .B(_10881_), .Y(_10882_));
NAND_g _17380_ (.A(_10872_), .B(_10882_), .Y(_10883_));
NAND_g _17381_ (.A(_00007_[1]), .B(_10883_), .Y(_10884_));
NOR_g _17382_ (.A(cpuregs[16][2]), .B(_00007_[2]), .Y(_10885_));
NOR_g _17383_ (.A(cpuregs[20][2]), .B(_09027_), .Y(_10886_));
NOR_g _17384_ (.A(_10885_), .B(_10886_), .Y(_10887_));
NOR_g _17385_ (.A(cpuregs[17][2]), .B(_00007_[2]), .Y(_10888_));
NAND_g _17386_ (.A(_08983_), .B(_00007_[2]), .Y(_10889_));
NOR_g _17387_ (.A(cpuregs[24][2]), .B(_00007_[2]), .Y(_10890_));
NOR_g _17388_ (.A(cpuregs[28][2]), .B(_09027_), .Y(_10891_));
NOR_g _17389_ (.A(_10890_), .B(_10891_), .Y(_10892_));
NOR_g _17390_ (.A(cpuregs[25][2]), .B(_00007_[2]), .Y(_10893_));
NAND_g _17391_ (.A(_08876_), .B(_00007_[2]), .Y(_10894_));
NAND_g _17392_ (.A(_09025_), .B(_10887_), .Y(_10895_));
NOR_g _17393_ (.A(_09025_), .B(_10888_), .Y(_10896_));
NAND_g _17394_ (.A(_10889_), .B(_10896_), .Y(_10897_));
AND_g _17395_ (.A(_10895_), .B(_10897_), .Y(_10898_));
NAND_g _17396_ (.A(_09028_), .B(_10898_), .Y(_10899_));
NOR_g _17397_ (.A(_09025_), .B(_10893_), .Y(_10900_));
NAND_g _17398_ (.A(_10894_), .B(_10900_), .Y(_10901_));
NAND_g _17399_ (.A(_09025_), .B(_10892_), .Y(_10902_));
AND_g _17400_ (.A(_10901_), .B(_10902_), .Y(_10903_));
NAND_g _17401_ (.A(_00007_[3]), .B(_10903_), .Y(_10904_));
AND_g _17402_ (.A(_10899_), .B(_10904_), .Y(_10905_));
NAND_g _17403_ (.A(_09026_), .B(_10905_), .Y(_10906_));
NAND_g _17404_ (.A(cpuregs[6][2]), .B(_00007_[2]), .Y(_10907_));
NAND_g _17405_ (.A(cpuregs[2][2]), .B(_09027_), .Y(_10908_));
AND_g _17406_ (.A(_10907_), .B(_10908_), .Y(_10909_));
NAND_g _17407_ (.A(_09025_), .B(_10909_), .Y(_10910_));
NAND_g _17408_ (.A(cpuregs[7][2]), .B(_00007_[2]), .Y(_10911_));
NAND_g _17409_ (.A(cpuregs[3][2]), .B(_09027_), .Y(_10912_));
AND_g _17410_ (.A(_00007_[0]), .B(_10912_), .Y(_10913_));
NAND_g _17411_ (.A(_10911_), .B(_10913_), .Y(_10914_));
AND_g _17412_ (.A(_09028_), .B(_10914_), .Y(_10915_));
NAND_g _17413_ (.A(_10910_), .B(_10915_), .Y(_10916_));
NOR_g _17414_ (.A(cpuregs[10][2]), .B(_00007_[2]), .Y(_10917_));
NOR_g _17415_ (.A(cpuregs[14][2]), .B(_09027_), .Y(_10918_));
NOR_g _17416_ (.A(_10917_), .B(_10918_), .Y(_10919_));
NOR_g _17417_ (.A(cpuregs[11][2]), .B(_00007_[2]), .Y(_10920_));
NOT_g _17418_ (.A(_10920_), .Y(_10921_));
NAND_g _17419_ (.A(_08808_), .B(_00007_[2]), .Y(_10922_));
AND_g _17420_ (.A(_00007_[0]), .B(_10922_), .Y(_10923_));
NAND_g _17421_ (.A(_10921_), .B(_10923_), .Y(_10924_));
NAND_g _17422_ (.A(_09025_), .B(_10919_), .Y(_10925_));
NAND_g _17423_ (.A(_10924_), .B(_10925_), .Y(_10926_));
NAND_g _17424_ (.A(_00007_[3]), .B(_10926_), .Y(_10927_));
NAND_g _17425_ (.A(_10916_), .B(_10927_), .Y(_10928_));
NAND_g _17426_ (.A(_00007_[1]), .B(_10928_), .Y(_10929_));
NAND_g _17427_ (.A(cpuregs[4][2]), .B(_00007_[2]), .Y(_10930_));
NAND_g _17428_ (.A(cpuregs[0][2]), .B(_09027_), .Y(_10931_));
AND_g _17429_ (.A(_09025_), .B(_10931_), .Y(_10932_));
NAND_g _17430_ (.A(_10930_), .B(_10932_), .Y(_10933_));
NAND_g _17431_ (.A(cpuregs[1][2]), .B(_09027_), .Y(_10934_));
NAND_g _17432_ (.A(cpuregs[5][2]), .B(_00007_[2]), .Y(_10935_));
AND_g _17433_ (.A(_00007_[0]), .B(_10935_), .Y(_10936_));
NAND_g _17434_ (.A(_10934_), .B(_10936_), .Y(_10937_));
NOR_g _17435_ (.A(cpuregs[9][2]), .B(_00007_[2]), .Y(_10938_));
NAND_g _17436_ (.A(_08926_), .B(_00007_[2]), .Y(_10939_));
NOR_g _17437_ (.A(cpuregs[8][2]), .B(_00007_[2]), .Y(_10940_));
NOR_g _17438_ (.A(cpuregs[12][2]), .B(_09027_), .Y(_10941_));
NOR_g _17439_ (.A(_10940_), .B(_10941_), .Y(_10942_));
NAND_g _17440_ (.A(_10933_), .B(_10937_), .Y(_10943_));
NAND_g _17441_ (.A(_09028_), .B(_10943_), .Y(_10944_));
NAND_g _17442_ (.A(_09025_), .B(_10942_), .Y(_10945_));
NOR_g _17443_ (.A(_09025_), .B(_10938_), .Y(_10946_));
NAND_g _17444_ (.A(_10939_), .B(_10946_), .Y(_10947_));
AND_g _17445_ (.A(_00007_[3]), .B(_10947_), .Y(_10948_));
NAND_g _17446_ (.A(_10945_), .B(_10948_), .Y(_10949_));
AND_g _17447_ (.A(_10944_), .B(_10949_), .Y(_10950_));
NAND_g _17448_ (.A(_09026_), .B(_10950_), .Y(_10951_));
AND_g _17449_ (.A(_10929_), .B(_10951_), .Y(_10952_));
AND_g _17450_ (.A(_00007_[4]), .B(_10884_), .Y(_10953_));
NAND_g _17451_ (.A(_10906_), .B(_10953_), .Y(_10954_));
NAND_g _17452_ (.A(_09029_), .B(_10952_), .Y(_10955_));
AND_g _17453_ (.A(_10954_), .B(_10955_), .Y(_10956_));
AND_g _17454_ (.A(_10611_), .B(_10956_), .Y(_10957_));
NAND_g _17455_ (.A(_10599_), .B(_10957_), .Y(_10958_));
NAND_g _17456_ (.A(_10754_), .B(_10957_), .Y(_10959_));
AND_g _17457_ (.A(_10958_), .B(_10959_), .Y(_10960_));
NAND_g _17458_ (.A(_10862_), .B(_10960_), .Y(_10961_));
NAND_g _17459_ (.A(_10603_), .B(_10961_), .Y(_10962_));
NAND_g _17460_ (.A(pcpi_rs2[2]), .B(_10604_), .Y(_10963_));
NAND_g _17461_ (.A(_10962_), .B(_10963_), .Y(_00277_));
NAND_g _17462_ (.A(cpuregs[29][3]), .B(_00007_[2]), .Y(_10964_));
NAND_g _17463_ (.A(cpuregs[25][3]), .B(_09027_), .Y(_10965_));
AND_g _17464_ (.A(_00007_[0]), .B(_10965_), .Y(_10966_));
NAND_g _17465_ (.A(_10964_), .B(_10966_), .Y(_10967_));
NAND_g _17466_ (.A(cpuregs[24][3]), .B(_09027_), .Y(_10968_));
NAND_g _17467_ (.A(cpuregs[28][3]), .B(_00007_[2]), .Y(_10969_));
AND_g _17468_ (.A(_09025_), .B(_10969_), .Y(_10970_));
NAND_g _17469_ (.A(_10968_), .B(_10970_), .Y(_10971_));
AND_g _17470_ (.A(_09026_), .B(_10971_), .Y(_10972_));
NAND_g _17471_ (.A(_10967_), .B(_10972_), .Y(_10973_));
NAND_g _17472_ (.A(cpuregs[27][3]), .B(_09027_), .Y(_10974_));
NAND_g _17473_ (.A(cpuregs[31][3]), .B(_00007_[2]), .Y(_10975_));
AND_g _17474_ (.A(_00007_[0]), .B(_10975_), .Y(_10976_));
NAND_g _17475_ (.A(_10974_), .B(_10976_), .Y(_10977_));
NAND_g _17476_ (.A(cpuregs[26][3]), .B(_09027_), .Y(_10978_));
NAND_g _17477_ (.A(cpuregs[30][3]), .B(_00007_[2]), .Y(_10979_));
AND_g _17478_ (.A(_09025_), .B(_10979_), .Y(_10980_));
NAND_g _17479_ (.A(_10978_), .B(_10980_), .Y(_10981_));
AND_g _17480_ (.A(_00007_[1]), .B(_10981_), .Y(_10982_));
NAND_g _17481_ (.A(_10977_), .B(_10982_), .Y(_10983_));
NAND_g _17482_ (.A(_10973_), .B(_10983_), .Y(_10984_));
NAND_g _17483_ (.A(_00007_[4]), .B(_10984_), .Y(_10985_));
NAND_g _17484_ (.A(cpuregs[14][3]), .B(_09025_), .Y(_10986_));
NAND_g _17485_ (.A(cpuregs[15][3]), .B(_00007_[0]), .Y(_10987_));
NAND_g _17486_ (.A(_10986_), .B(_10987_), .Y(_10988_));
NAND_g _17487_ (.A(_00007_[2]), .B(_10988_), .Y(_10989_));
NAND_g _17488_ (.A(cpuregs[10][3]), .B(_09025_), .Y(_10990_));
NAND_g _17489_ (.A(cpuregs[11][3]), .B(_00007_[0]), .Y(_10991_));
NAND_g _17490_ (.A(_10990_), .B(_10991_), .Y(_10992_));
NAND_g _17491_ (.A(_09027_), .B(_10992_), .Y(_10993_));
NAND_g _17492_ (.A(_10989_), .B(_10993_), .Y(_10994_));
NAND_g _17493_ (.A(_00007_[1]), .B(_10994_), .Y(_10995_));
NAND_g _17494_ (.A(cpuregs[12][3]), .B(_09025_), .Y(_10996_));
NAND_g _17495_ (.A(cpuregs[13][3]), .B(_00007_[0]), .Y(_10997_));
NAND_g _17496_ (.A(_10996_), .B(_10997_), .Y(_10998_));
NAND_g _17497_ (.A(_00007_[2]), .B(_10998_), .Y(_10999_));
NAND_g _17498_ (.A(cpuregs[8][3]), .B(_09025_), .Y(_11000_));
NAND_g _17499_ (.A(cpuregs[9][3]), .B(_00007_[0]), .Y(_11001_));
NAND_g _17500_ (.A(_11000_), .B(_11001_), .Y(_11002_));
NAND_g _17501_ (.A(_09027_), .B(_11002_), .Y(_11003_));
NAND_g _17502_ (.A(_10999_), .B(_11003_), .Y(_11004_));
NAND_g _17503_ (.A(_09026_), .B(_11004_), .Y(_11005_));
NAND_g _17504_ (.A(_10995_), .B(_11005_), .Y(_11006_));
AND_g _17505_ (.A(_09029_), .B(_11006_), .Y(_11007_));
NOT_g _17506_ (.A(_11007_), .Y(_11008_));
NAND_g _17507_ (.A(_10985_), .B(_11008_), .Y(_11009_));
NAND_g _17508_ (.A(_00007_[3]), .B(_11009_), .Y(_11010_));
NAND_g _17509_ (.A(cpuregs[1][3]), .B(_09027_), .Y(_11011_));
NAND_g _17510_ (.A(cpuregs[5][3]), .B(_00007_[2]), .Y(_11012_));
AND_g _17511_ (.A(_00007_[0]), .B(_11012_), .Y(_11013_));
NAND_g _17512_ (.A(_11011_), .B(_11013_), .Y(_11014_));
NAND_g _17513_ (.A(cpuregs[0][3]), .B(_09027_), .Y(_11015_));
NAND_g _17514_ (.A(cpuregs[4][3]), .B(_00007_[2]), .Y(_11016_));
AND_g _17515_ (.A(_09025_), .B(_11016_), .Y(_11017_));
NAND_g _17516_ (.A(_11015_), .B(_11017_), .Y(_11018_));
AND_g _17517_ (.A(_09026_), .B(_11018_), .Y(_11019_));
NAND_g _17518_ (.A(_11014_), .B(_11019_), .Y(_11020_));
NAND_g _17519_ (.A(cpuregs[3][3]), .B(_09027_), .Y(_11021_));
NAND_g _17520_ (.A(cpuregs[7][3]), .B(_00007_[2]), .Y(_11022_));
AND_g _17521_ (.A(_00007_[0]), .B(_11022_), .Y(_11023_));
NAND_g _17522_ (.A(_11021_), .B(_11023_), .Y(_11024_));
NAND_g _17523_ (.A(cpuregs[2][3]), .B(_09027_), .Y(_11025_));
NAND_g _17524_ (.A(cpuregs[6][3]), .B(_00007_[2]), .Y(_11026_));
AND_g _17525_ (.A(_09025_), .B(_11026_), .Y(_11027_));
NAND_g _17526_ (.A(_11025_), .B(_11027_), .Y(_11028_));
AND_g _17527_ (.A(_00007_[1]), .B(_11028_), .Y(_11029_));
NAND_g _17528_ (.A(_11024_), .B(_11029_), .Y(_11030_));
NAND_g _17529_ (.A(_11020_), .B(_11030_), .Y(_11031_));
NAND_g _17530_ (.A(_09029_), .B(_11031_), .Y(_11032_));
NAND_g _17531_ (.A(cpuregs[19][3]), .B(_00007_[1]), .Y(_11033_));
NAND_g _17532_ (.A(cpuregs[17][3]), .B(_09026_), .Y(_11034_));
NAND_g _17533_ (.A(_11033_), .B(_11034_), .Y(_11035_));
NAND_g _17534_ (.A(_09027_), .B(_11035_), .Y(_11036_));
NAND_g _17535_ (.A(cpuregs[23][3]), .B(_00007_[1]), .Y(_11037_));
NAND_g _17536_ (.A(cpuregs[21][3]), .B(_09026_), .Y(_11038_));
NAND_g _17537_ (.A(_11037_), .B(_11038_), .Y(_11039_));
NAND_g _17538_ (.A(_00007_[2]), .B(_11039_), .Y(_11040_));
AND_g _17539_ (.A(_00007_[0]), .B(_11040_), .Y(_11041_));
NAND_g _17540_ (.A(_11036_), .B(_11041_), .Y(_11042_));
NAND_g _17541_ (.A(cpuregs[18][3]), .B(_00007_[1]), .Y(_11043_));
NAND_g _17542_ (.A(cpuregs[16][3]), .B(_09026_), .Y(_11044_));
NAND_g _17543_ (.A(_11043_), .B(_11044_), .Y(_11045_));
NAND_g _17544_ (.A(_09027_), .B(_11045_), .Y(_11046_));
NAND_g _17545_ (.A(cpuregs[22][3]), .B(_00007_[1]), .Y(_11047_));
NAND_g _17546_ (.A(cpuregs[20][3]), .B(_09026_), .Y(_11048_));
NAND_g _17547_ (.A(_11047_), .B(_11048_), .Y(_11049_));
NAND_g _17548_ (.A(_00007_[2]), .B(_11049_), .Y(_11050_));
AND_g _17549_ (.A(_09025_), .B(_11050_), .Y(_11051_));
NAND_g _17550_ (.A(_11046_), .B(_11051_), .Y(_11052_));
AND_g _17551_ (.A(_00007_[4]), .B(_11052_), .Y(_11053_));
NAND_g _17552_ (.A(_11042_), .B(_11053_), .Y(_11054_));
NAND_g _17553_ (.A(_11032_), .B(_11054_), .Y(_11055_));
NAND_g _17554_ (.A(_09028_), .B(_11055_), .Y(_11056_));
NAND_g _17555_ (.A(_11010_), .B(_11056_), .Y(_11057_));
AND_g _17556_ (.A(_10611_), .B(_11057_), .Y(_11058_));
NAND_g _17557_ (.A(_10754_), .B(_11058_), .Y(_11059_));
NAND_g _17558_ (.A(_10599_), .B(_11058_), .Y(_11060_));
NAND_g _17559_ (.A(decoded_imm[3]), .B(_10606_), .Y(_11061_));
NOR_g _17560_ (.A(pcpi_rs2[3]), .B(_10603_), .Y(_11062_));
AND_g _17561_ (.A(_10603_), .B(_11061_), .Y(_11063_));
AND_g _17562_ (.A(_11059_), .B(_11063_), .Y(_11064_));
AND_g _17563_ (.A(_11060_), .B(_11064_), .Y(_11065_));
NOR_g _17564_ (.A(_11062_), .B(_11065_), .Y(_00278_));
NAND_g _17565_ (.A(decoded_imm[4]), .B(_10606_), .Y(_11066_));
NAND_g _17566_ (.A(cpuregs[19][4]), .B(_09027_), .Y(_11067_));
NAND_g _17567_ (.A(cpuregs[23][4]), .B(_00007_[2]), .Y(_11068_));
AND_g _17568_ (.A(_00007_[0]), .B(_11068_), .Y(_11069_));
NAND_g _17569_ (.A(_11067_), .B(_11069_), .Y(_11070_));
NAND_g _17570_ (.A(cpuregs[18][4]), .B(_09027_), .Y(_11071_));
NAND_g _17571_ (.A(cpuregs[22][4]), .B(_00007_[2]), .Y(_11072_));
AND_g _17572_ (.A(_09025_), .B(_11072_), .Y(_11073_));
NAND_g _17573_ (.A(_11071_), .B(_11073_), .Y(_11074_));
AND_g _17574_ (.A(_09028_), .B(_11074_), .Y(_11075_));
NAND_g _17575_ (.A(_11070_), .B(_11075_), .Y(_11076_));
NAND_g _17576_ (.A(cpuregs[27][4]), .B(_09027_), .Y(_11077_));
NAND_g _17577_ (.A(cpuregs[31][4]), .B(_00007_[2]), .Y(_11078_));
AND_g _17578_ (.A(_00007_[0]), .B(_11078_), .Y(_11079_));
NAND_g _17579_ (.A(_11077_), .B(_11079_), .Y(_11080_));
NAND_g _17580_ (.A(cpuregs[26][4]), .B(_09027_), .Y(_11081_));
NAND_g _17581_ (.A(cpuregs[30][4]), .B(_00007_[2]), .Y(_11082_));
AND_g _17582_ (.A(_09025_), .B(_11082_), .Y(_11083_));
NAND_g _17583_ (.A(_11081_), .B(_11083_), .Y(_11084_));
AND_g _17584_ (.A(_00007_[3]), .B(_11084_), .Y(_11085_));
NAND_g _17585_ (.A(_11080_), .B(_11085_), .Y(_11086_));
NAND_g _17586_ (.A(_11076_), .B(_11086_), .Y(_11087_));
NAND_g _17587_ (.A(_00007_[1]), .B(_11087_), .Y(_11088_));
NOR_g _17588_ (.A(cpuregs[16][4]), .B(_00007_[2]), .Y(_11089_));
NOR_g _17589_ (.A(cpuregs[20][4]), .B(_09027_), .Y(_11090_));
NOR_g _17590_ (.A(_11089_), .B(_11090_), .Y(_11091_));
NOR_g _17591_ (.A(cpuregs[17][4]), .B(_00007_[2]), .Y(_11092_));
NAND_g _17592_ (.A(_08984_), .B(_00007_[2]), .Y(_11093_));
NOR_g _17593_ (.A(cpuregs[24][4]), .B(_00007_[2]), .Y(_11094_));
NOR_g _17594_ (.A(cpuregs[28][4]), .B(_09027_), .Y(_11095_));
NOR_g _17595_ (.A(_11094_), .B(_11095_), .Y(_11096_));
NOR_g _17596_ (.A(cpuregs[25][4]), .B(_00007_[2]), .Y(_11097_));
NAND_g _17597_ (.A(_08877_), .B(_00007_[2]), .Y(_11098_));
NAND_g _17598_ (.A(_09025_), .B(_11091_), .Y(_11099_));
NOR_g _17599_ (.A(_09025_), .B(_11092_), .Y(_11100_));
NAND_g _17600_ (.A(_11093_), .B(_11100_), .Y(_11101_));
AND_g _17601_ (.A(_11099_), .B(_11101_), .Y(_11102_));
NAND_g _17602_ (.A(_09028_), .B(_11102_), .Y(_11103_));
NOR_g _17603_ (.A(_09025_), .B(_11097_), .Y(_11104_));
NAND_g _17604_ (.A(_11098_), .B(_11104_), .Y(_11105_));
NAND_g _17605_ (.A(_09025_), .B(_11096_), .Y(_11106_));
AND_g _17606_ (.A(_11105_), .B(_11106_), .Y(_11107_));
NAND_g _17607_ (.A(_00007_[3]), .B(_11107_), .Y(_11108_));
AND_g _17608_ (.A(_11103_), .B(_11108_), .Y(_11109_));
NAND_g _17609_ (.A(_09026_), .B(_11109_), .Y(_11110_));
NAND_g _17610_ (.A(cpuregs[14][4]), .B(_09025_), .Y(_11111_));
NAND_g _17611_ (.A(cpuregs[15][4]), .B(_00007_[0]), .Y(_11112_));
NAND_g _17612_ (.A(_11111_), .B(_11112_), .Y(_11113_));
NAND_g _17613_ (.A(_00007_[2]), .B(_11113_), .Y(_11114_));
NAND_g _17614_ (.A(cpuregs[10][4]), .B(_09025_), .Y(_11115_));
NAND_g _17615_ (.A(cpuregs[11][4]), .B(_00007_[0]), .Y(_11116_));
NAND_g _17616_ (.A(_11115_), .B(_11116_), .Y(_11117_));
NAND_g _17617_ (.A(_09027_), .B(_11117_), .Y(_11118_));
NAND_g _17618_ (.A(_11114_), .B(_11118_), .Y(_11119_));
NAND_g _17619_ (.A(_00007_[3]), .B(_11119_), .Y(_11120_));
NAND_g _17620_ (.A(cpuregs[6][4]), .B(_09025_), .Y(_11121_));
NAND_g _17621_ (.A(cpuregs[7][4]), .B(_00007_[0]), .Y(_11122_));
NAND_g _17622_ (.A(_11121_), .B(_11122_), .Y(_11123_));
NAND_g _17623_ (.A(_00007_[2]), .B(_11123_), .Y(_11124_));
NAND_g _17624_ (.A(cpuregs[2][4]), .B(_09025_), .Y(_11125_));
NAND_g _17625_ (.A(cpuregs[3][4]), .B(_00007_[0]), .Y(_11126_));
NAND_g _17626_ (.A(_11125_), .B(_11126_), .Y(_11127_));
NAND_g _17627_ (.A(_09027_), .B(_11127_), .Y(_11128_));
NAND_g _17628_ (.A(_11124_), .B(_11128_), .Y(_11129_));
NAND_g _17629_ (.A(_09028_), .B(_11129_), .Y(_11130_));
NAND_g _17630_ (.A(_11120_), .B(_11130_), .Y(_11131_));
NAND_g _17631_ (.A(_00007_[1]), .B(_11131_), .Y(_11132_));
NOR_g _17632_ (.A(cpuregs[9][4]), .B(_00007_[2]), .Y(_11133_));
NOT_g _17633_ (.A(_11133_), .Y(_11134_));
NAND_g _17634_ (.A(_08927_), .B(_00007_[2]), .Y(_11135_));
AND_g _17635_ (.A(_00007_[0]), .B(_11135_), .Y(_11136_));
NAND_g _17636_ (.A(_11134_), .B(_11136_), .Y(_11137_));
NOR_g _17637_ (.A(cpuregs[8][4]), .B(_00007_[2]), .Y(_11138_));
NOR_g _17638_ (.A(cpuregs[12][4]), .B(_09027_), .Y(_11139_));
NOR_g _17639_ (.A(_11138_), .B(_11139_), .Y(_11140_));
NAND_g _17640_ (.A(_09025_), .B(_11140_), .Y(_11141_));
NAND_g _17641_ (.A(_11137_), .B(_11141_), .Y(_11142_));
NAND_g _17642_ (.A(_00007_[3]), .B(_11142_), .Y(_11143_));
NAND_g _17643_ (.A(cpuregs[4][4]), .B(_00007_[2]), .Y(_11144_));
NAND_g _17644_ (.A(cpuregs[0][4]), .B(_09027_), .Y(_11145_));
AND_g _17645_ (.A(_11144_), .B(_11145_), .Y(_11146_));
NAND_g _17646_ (.A(_09025_), .B(_11146_), .Y(_11147_));
NAND_g _17647_ (.A(cpuregs[5][4]), .B(_00007_[2]), .Y(_11148_));
NAND_g _17648_ (.A(cpuregs[1][4]), .B(_09027_), .Y(_11149_));
AND_g _17649_ (.A(_00007_[0]), .B(_11149_), .Y(_11150_));
NAND_g _17650_ (.A(_11148_), .B(_11150_), .Y(_11151_));
AND_g _17651_ (.A(_09028_), .B(_11151_), .Y(_11152_));
NAND_g _17652_ (.A(_11147_), .B(_11152_), .Y(_11153_));
NAND_g _17653_ (.A(_11143_), .B(_11153_), .Y(_11154_));
NAND_g _17654_ (.A(_09026_), .B(_11154_), .Y(_11155_));
AND_g _17655_ (.A(_11132_), .B(_11155_), .Y(_11156_));
AND_g _17656_ (.A(_00007_[4]), .B(_11088_), .Y(_11157_));
NAND_g _17657_ (.A(_11110_), .B(_11157_), .Y(_11158_));
NAND_g _17658_ (.A(_09029_), .B(_11156_), .Y(_11159_));
AND_g _17659_ (.A(_11158_), .B(_11159_), .Y(_11160_));
AND_g _17660_ (.A(_10611_), .B(_11160_), .Y(_11161_));
NAND_g _17661_ (.A(_10599_), .B(_11161_), .Y(_11162_));
NAND_g _17662_ (.A(_10754_), .B(_11161_), .Y(_11163_));
AND_g _17663_ (.A(_11162_), .B(_11163_), .Y(_11164_));
NAND_g _17664_ (.A(_11066_), .B(_11164_), .Y(_11165_));
NAND_g _17665_ (.A(_10603_), .B(_11165_), .Y(_11166_));
NAND_g _17666_ (.A(pcpi_rs2[4]), .B(_10604_), .Y(_11167_));
NAND_g _17667_ (.A(_11166_), .B(_11167_), .Y(_00279_));
NAND_g _17668_ (.A(_08815_), .B(_10604_), .Y(_11168_));
NAND_g _17669_ (.A(_10600_), .B(_10755_), .Y(_11169_));
AND_g _17670_ (.A(_10611_), .B(_11169_), .Y(_11170_));
NAND_g _17671_ (.A(cpuregs[13][5]), .B(_00007_[2]), .Y(_11171_));
NAND_g _17672_ (.A(cpuregs[9][5]), .B(_09027_), .Y(_11172_));
AND_g _17673_ (.A(_00007_[0]), .B(_11172_), .Y(_11173_));
NAND_g _17674_ (.A(_11171_), .B(_11173_), .Y(_11174_));
NAND_g _17675_ (.A(cpuregs[8][5]), .B(_09027_), .Y(_11175_));
NAND_g _17676_ (.A(cpuregs[12][5]), .B(_00007_[2]), .Y(_11176_));
AND_g _17677_ (.A(_09025_), .B(_11176_), .Y(_11177_));
NAND_g _17678_ (.A(_11175_), .B(_11177_), .Y(_11178_));
AND_g _17679_ (.A(_00007_[3]), .B(_11178_), .Y(_11179_));
NAND_g _17680_ (.A(_11174_), .B(_11179_), .Y(_11180_));
NAND_g _17681_ (.A(cpuregs[1][5]), .B(_09027_), .Y(_11181_));
NAND_g _17682_ (.A(cpuregs[5][5]), .B(_00007_[2]), .Y(_11182_));
AND_g _17683_ (.A(_00007_[0]), .B(_11182_), .Y(_11183_));
NAND_g _17684_ (.A(_11181_), .B(_11183_), .Y(_11184_));
NAND_g _17685_ (.A(cpuregs[0][5]), .B(_09027_), .Y(_11185_));
NAND_g _17686_ (.A(cpuregs[4][5]), .B(_00007_[2]), .Y(_11186_));
AND_g _17687_ (.A(_09025_), .B(_11186_), .Y(_11187_));
NAND_g _17688_ (.A(_11185_), .B(_11187_), .Y(_11188_));
AND_g _17689_ (.A(_09028_), .B(_11184_), .Y(_11189_));
NAND_g _17690_ (.A(_11188_), .B(_11189_), .Y(_11190_));
NAND_g _17691_ (.A(cpuregs[3][5]), .B(_09027_), .Y(_11191_));
NAND_g _17692_ (.A(cpuregs[7][5]), .B(_00007_[2]), .Y(_11192_));
AND_g _17693_ (.A(_00007_[0]), .B(_11192_), .Y(_11193_));
NAND_g _17694_ (.A(_11191_), .B(_11193_), .Y(_11194_));
NAND_g _17695_ (.A(cpuregs[2][5]), .B(_09027_), .Y(_11195_));
NAND_g _17696_ (.A(cpuregs[6][5]), .B(_00007_[2]), .Y(_11196_));
AND_g _17697_ (.A(_09025_), .B(_11196_), .Y(_11197_));
NAND_g _17698_ (.A(_11195_), .B(_11197_), .Y(_11198_));
AND_g _17699_ (.A(_09028_), .B(_11194_), .Y(_11199_));
NAND_g _17700_ (.A(_11198_), .B(_11199_), .Y(_11200_));
NAND_g _17701_ (.A(cpuregs[15][5]), .B(_00007_[2]), .Y(_11201_));
NAND_g _17702_ (.A(cpuregs[11][5]), .B(_09027_), .Y(_11202_));
AND_g _17703_ (.A(_00007_[0]), .B(_11202_), .Y(_11203_));
NAND_g _17704_ (.A(_11201_), .B(_11203_), .Y(_11204_));
NAND_g _17705_ (.A(cpuregs[10][5]), .B(_09027_), .Y(_11205_));
NAND_g _17706_ (.A(cpuregs[14][5]), .B(_00007_[2]), .Y(_11206_));
AND_g _17707_ (.A(_09025_), .B(_11206_), .Y(_11207_));
NAND_g _17708_ (.A(_11205_), .B(_11207_), .Y(_11208_));
AND_g _17709_ (.A(_00007_[3]), .B(_11208_), .Y(_11209_));
NAND_g _17710_ (.A(_11204_), .B(_11209_), .Y(_11210_));
NAND_g _17711_ (.A(_11200_), .B(_11210_), .Y(_11211_));
NAND_g _17712_ (.A(_00007_[1]), .B(_11211_), .Y(_11212_));
NAND_g _17713_ (.A(_11180_), .B(_11190_), .Y(_11213_));
NAND_g _17714_ (.A(_09026_), .B(_11213_), .Y(_11214_));
AND_g _17715_ (.A(_11212_), .B(_11214_), .Y(_11215_));
NAND_g _17716_ (.A(_09029_), .B(_11215_), .Y(_11216_));
NAND_g _17717_ (.A(cpuregs[25][5]), .B(_09027_), .Y(_11217_));
NAND_g _17718_ (.A(cpuregs[29][5]), .B(_00007_[2]), .Y(_11218_));
AND_g _17719_ (.A(_00007_[0]), .B(_11218_), .Y(_11219_));
NAND_g _17720_ (.A(_11217_), .B(_11219_), .Y(_11220_));
NAND_g _17721_ (.A(cpuregs[24][5]), .B(_09027_), .Y(_11221_));
NAND_g _17722_ (.A(cpuregs[28][5]), .B(_00007_[2]), .Y(_11222_));
AND_g _17723_ (.A(_09025_), .B(_11222_), .Y(_11223_));
NAND_g _17724_ (.A(_11221_), .B(_11223_), .Y(_11224_));
AND_g _17725_ (.A(_00007_[3]), .B(_11224_), .Y(_11225_));
NAND_g _17726_ (.A(_11220_), .B(_11225_), .Y(_11226_));
NAND_g _17727_ (.A(cpuregs[21][5]), .B(_00007_[2]), .Y(_11227_));
NAND_g _17728_ (.A(cpuregs[17][5]), .B(_09027_), .Y(_11228_));
AND_g _17729_ (.A(_00007_[0]), .B(_11228_), .Y(_11229_));
NAND_g _17730_ (.A(_11227_), .B(_11229_), .Y(_11230_));
NAND_g _17731_ (.A(cpuregs[20][5]), .B(_00007_[2]), .Y(_11231_));
NAND_g _17732_ (.A(cpuregs[16][5]), .B(_09027_), .Y(_11232_));
AND_g _17733_ (.A(_09025_), .B(_11232_), .Y(_11233_));
NAND_g _17734_ (.A(_11231_), .B(_11233_), .Y(_11234_));
AND_g _17735_ (.A(_09028_), .B(_11234_), .Y(_11235_));
NAND_g _17736_ (.A(_11230_), .B(_11235_), .Y(_11236_));
AND_g _17737_ (.A(_09026_), .B(_11236_), .Y(_11237_));
NAND_g _17738_ (.A(_11226_), .B(_11237_), .Y(_11238_));
NAND_g _17739_ (.A(cpuregs[27][5]), .B(_09027_), .Y(_11239_));
NAND_g _17740_ (.A(cpuregs[31][5]), .B(_00007_[2]), .Y(_11240_));
AND_g _17741_ (.A(_00007_[0]), .B(_11240_), .Y(_11241_));
NAND_g _17742_ (.A(_11239_), .B(_11241_), .Y(_11242_));
NAND_g _17743_ (.A(cpuregs[26][5]), .B(_09027_), .Y(_11243_));
NAND_g _17744_ (.A(cpuregs[30][5]), .B(_00007_[2]), .Y(_11244_));
AND_g _17745_ (.A(_09025_), .B(_11244_), .Y(_11245_));
NAND_g _17746_ (.A(_11243_), .B(_11245_), .Y(_11246_));
AND_g _17747_ (.A(_00007_[3]), .B(_11246_), .Y(_11247_));
NAND_g _17748_ (.A(_11242_), .B(_11247_), .Y(_11248_));
NAND_g _17749_ (.A(cpuregs[19][5]), .B(_09027_), .Y(_11249_));
NAND_g _17750_ (.A(cpuregs[23][5]), .B(_00007_[2]), .Y(_11250_));
AND_g _17751_ (.A(_00007_[0]), .B(_11250_), .Y(_11251_));
NAND_g _17752_ (.A(_11249_), .B(_11251_), .Y(_11252_));
NAND_g _17753_ (.A(cpuregs[18][5]), .B(_09027_), .Y(_11253_));
NAND_g _17754_ (.A(cpuregs[22][5]), .B(_00007_[2]), .Y(_11254_));
AND_g _17755_ (.A(_09025_), .B(_11254_), .Y(_11255_));
NAND_g _17756_ (.A(_11253_), .B(_11255_), .Y(_11256_));
AND_g _17757_ (.A(_09028_), .B(_11256_), .Y(_11257_));
NAND_g _17758_ (.A(_11252_), .B(_11257_), .Y(_11258_));
AND_g _17759_ (.A(_00007_[1]), .B(_11258_), .Y(_11259_));
NAND_g _17760_ (.A(_11248_), .B(_11259_), .Y(_11260_));
NAND_g _17761_ (.A(_11238_), .B(_11260_), .Y(_11261_));
NAND_g _17762_ (.A(_00007_[4]), .B(_11261_), .Y(_11262_));
AND_g _17763_ (.A(_11216_), .B(_11262_), .Y(_11263_));
NAND_g _17764_ (.A(_11170_), .B(_11263_), .Y(_11264_));
NAND_g _17765_ (.A(decoded_imm[5]), .B(_10606_), .Y(_11265_));
AND_g _17766_ (.A(_10603_), .B(_11265_), .Y(_11266_));
NAND_g _17767_ (.A(_11264_), .B(_11266_), .Y(_11267_));
AND_g _17768_ (.A(_11168_), .B(_11267_), .Y(_00280_));
NAND_g _17769_ (.A(_08816_), .B(_10604_), .Y(_11268_));
NAND_g _17770_ (.A(_09004_), .B(_00007_[2]), .Y(_11269_));
NOR_g _17771_ (.A(cpuregs[2][6]), .B(_00007_[2]), .Y(_11270_));
NOR_g _17772_ (.A(_00007_[0]), .B(_11270_), .Y(_11271_));
NAND_g _17773_ (.A(_11269_), .B(_11271_), .Y(_11272_));
NAND_g _17774_ (.A(_08964_), .B(_00007_[2]), .Y(_11273_));
NOR_g _17775_ (.A(cpuregs[3][6]), .B(_00007_[2]), .Y(_11274_));
NOR_g _17776_ (.A(_09025_), .B(_11274_), .Y(_11275_));
NAND_g _17777_ (.A(_11273_), .B(_11275_), .Y(_11276_));
NAND_g _17778_ (.A(_11272_), .B(_11276_), .Y(_11277_));
NAND_g _17779_ (.A(_09028_), .B(_11277_), .Y(_11278_));
NAND_g _17780_ (.A(cpuregs[11][6]), .B(_09027_), .Y(_11279_));
NAND_g _17781_ (.A(cpuregs[15][6]), .B(_00007_[2]), .Y(_11280_));
NAND_g _17782_ (.A(_11279_), .B(_11280_), .Y(_11281_));
NAND_g _17783_ (.A(_00007_[0]), .B(_11281_), .Y(_11282_));
NAND_g _17784_ (.A(cpuregs[14][6]), .B(_00007_[2]), .Y(_11283_));
NAND_g _17785_ (.A(cpuregs[10][6]), .B(_09027_), .Y(_11284_));
NAND_g _17786_ (.A(_11283_), .B(_11284_), .Y(_11285_));
NAND_g _17787_ (.A(_09025_), .B(_11285_), .Y(_11286_));
NAND_g _17788_ (.A(_11282_), .B(_11286_), .Y(_11287_));
NAND_g _17789_ (.A(_00007_[3]), .B(_11287_), .Y(_11288_));
AND_g _17790_ (.A(_09029_), .B(_11288_), .Y(_11289_));
NAND_g _17791_ (.A(_11278_), .B(_11289_), .Y(_11290_));
NAND_g _17792_ (.A(cpuregs[31][6]), .B(_00007_[2]), .Y(_11291_));
NAND_g _17793_ (.A(cpuregs[27][6]), .B(_09027_), .Y(_11292_));
AND_g _17794_ (.A(_00007_[0]), .B(_11292_), .Y(_11293_));
NAND_g _17795_ (.A(_11291_), .B(_11293_), .Y(_11294_));
NAND_g _17796_ (.A(cpuregs[26][6]), .B(_09027_), .Y(_11295_));
NAND_g _17797_ (.A(cpuregs[30][6]), .B(_00007_[2]), .Y(_11296_));
AND_g _17798_ (.A(_09025_), .B(_11296_), .Y(_11297_));
NAND_g _17799_ (.A(_11295_), .B(_11297_), .Y(_11298_));
AND_g _17800_ (.A(_00007_[3]), .B(_11298_), .Y(_11299_));
NAND_g _17801_ (.A(_11294_), .B(_11299_), .Y(_11300_));
NOR_g _17802_ (.A(cpuregs[18][6]), .B(_00007_[2]), .Y(_11301_));
NOT_g _17803_ (.A(_11301_), .Y(_11302_));
NAND_g _17804_ (.A(_08918_), .B(_00007_[2]), .Y(_11303_));
NAND_g _17805_ (.A(_11302_), .B(_11303_), .Y(_11304_));
NAND_g _17806_ (.A(_09025_), .B(_11304_), .Y(_11305_));
NAND_g _17807_ (.A(_08886_), .B(_00007_[2]), .Y(_11306_));
NOR_g _17808_ (.A(cpuregs[19][6]), .B(_00007_[2]), .Y(_11307_));
NOT_g _17809_ (.A(_11307_), .Y(_11308_));
NAND_g _17810_ (.A(_11306_), .B(_11308_), .Y(_11309_));
NAND_g _17811_ (.A(_00007_[0]), .B(_11309_), .Y(_11310_));
AND_g _17812_ (.A(_09028_), .B(_11310_), .Y(_11311_));
NAND_g _17813_ (.A(_11305_), .B(_11311_), .Y(_11312_));
AND_g _17814_ (.A(_00007_[4]), .B(_11312_), .Y(_11313_));
NAND_g _17815_ (.A(_11300_), .B(_11313_), .Y(_11314_));
NAND_g _17816_ (.A(_11290_), .B(_11314_), .Y(_11315_));
NAND_g _17817_ (.A(_00007_[1]), .B(_11315_), .Y(_11316_));
NAND_g _17818_ (.A(_08905_), .B(_00007_[2]), .Y(_11317_));
NOR_g _17819_ (.A(cpuregs[0][6]), .B(_00007_[2]), .Y(_11318_));
NOR_g _17820_ (.A(_00007_[0]), .B(_11318_), .Y(_11319_));
NAND_g _17821_ (.A(_11317_), .B(_11319_), .Y(_11320_));
NOR_g _17822_ (.A(cpuregs[1][6]), .B(_00007_[2]), .Y(_11321_));
NOT_g _17823_ (.A(_11321_), .Y(_11322_));
NAND_g _17824_ (.A(_08947_), .B(_00007_[2]), .Y(_11323_));
AND_g _17825_ (.A(_00007_[0]), .B(_11323_), .Y(_11324_));
NAND_g _17826_ (.A(_11322_), .B(_11324_), .Y(_11325_));
NAND_g _17827_ (.A(_11320_), .B(_11325_), .Y(_11326_));
NAND_g _17828_ (.A(_09028_), .B(_11326_), .Y(_11327_));
NAND_g _17829_ (.A(cpuregs[9][6]), .B(_09027_), .Y(_11328_));
NAND_g _17830_ (.A(cpuregs[13][6]), .B(_00007_[2]), .Y(_11329_));
NAND_g _17831_ (.A(_11328_), .B(_11329_), .Y(_11330_));
NAND_g _17832_ (.A(_00007_[0]), .B(_11330_), .Y(_11331_));
NAND_g _17833_ (.A(cpuregs[12][6]), .B(_00007_[2]), .Y(_11332_));
NAND_g _17834_ (.A(cpuregs[8][6]), .B(_09027_), .Y(_11333_));
NAND_g _17835_ (.A(_11332_), .B(_11333_), .Y(_11334_));
NAND_g _17836_ (.A(_09025_), .B(_11334_), .Y(_11335_));
NAND_g _17837_ (.A(_11331_), .B(_11335_), .Y(_11336_));
NAND_g _17838_ (.A(_00007_[3]), .B(_11336_), .Y(_11337_));
AND_g _17839_ (.A(_09029_), .B(_11337_), .Y(_11338_));
NAND_g _17840_ (.A(_11327_), .B(_11338_), .Y(_11339_));
NAND_g _17841_ (.A(cpuregs[29][6]), .B(_00007_[2]), .Y(_11340_));
NAND_g _17842_ (.A(cpuregs[25][6]), .B(_09027_), .Y(_11341_));
AND_g _17843_ (.A(_00007_[0]), .B(_11341_), .Y(_11342_));
NAND_g _17844_ (.A(_11340_), .B(_11342_), .Y(_11343_));
NAND_g _17845_ (.A(cpuregs[24][6]), .B(_09027_), .Y(_11344_));
NAND_g _17846_ (.A(cpuregs[28][6]), .B(_00007_[2]), .Y(_11345_));
AND_g _17847_ (.A(_09025_), .B(_11345_), .Y(_11346_));
NAND_g _17848_ (.A(_11344_), .B(_11346_), .Y(_11347_));
AND_g _17849_ (.A(_00007_[3]), .B(_11347_), .Y(_11348_));
NAND_g _17850_ (.A(_11343_), .B(_11348_), .Y(_11349_));
NOR_g _17851_ (.A(cpuregs[16][6]), .B(_00007_[2]), .Y(_11350_));
NOT_g _17852_ (.A(_11350_), .Y(_11351_));
NAND_g _17853_ (.A(_08844_), .B(_00007_[2]), .Y(_11352_));
NAND_g _17854_ (.A(_11351_), .B(_11352_), .Y(_11353_));
NAND_g _17855_ (.A(_09025_), .B(_11353_), .Y(_11354_));
NAND_g _17856_ (.A(_08941_), .B(_09027_), .Y(_11355_));
NAND_g _17857_ (.A(_08985_), .B(_00007_[2]), .Y(_11356_));
NAND_g _17858_ (.A(_11355_), .B(_11356_), .Y(_11357_));
NAND_g _17859_ (.A(_00007_[0]), .B(_11357_), .Y(_11358_));
AND_g _17860_ (.A(_09028_), .B(_11358_), .Y(_11359_));
NAND_g _17861_ (.A(_11354_), .B(_11359_), .Y(_11360_));
AND_g _17862_ (.A(_00007_[4]), .B(_11360_), .Y(_11361_));
NAND_g _17863_ (.A(_11349_), .B(_11361_), .Y(_11362_));
NAND_g _17864_ (.A(_11339_), .B(_11362_), .Y(_11363_));
NAND_g _17865_ (.A(_09026_), .B(_11363_), .Y(_11364_));
AND_g _17866_ (.A(_11316_), .B(_11364_), .Y(_11365_));
NAND_g _17867_ (.A(_11170_), .B(_11365_), .Y(_11366_));
NAND_g _17868_ (.A(decoded_imm[6]), .B(_10606_), .Y(_11367_));
AND_g _17869_ (.A(_10603_), .B(_11367_), .Y(_11368_));
NAND_g _17870_ (.A(_11366_), .B(_11368_), .Y(_11369_));
AND_g _17871_ (.A(_11268_), .B(_11369_), .Y(_00281_));
NAND_g _17872_ (.A(_08817_), .B(_10604_), .Y(_11370_));
NAND_g _17873_ (.A(cpuregs[14][7]), .B(_09025_), .Y(_11371_));
NAND_g _17874_ (.A(cpuregs[15][7]), .B(_00007_[0]), .Y(_11372_));
NAND_g _17875_ (.A(_11371_), .B(_11372_), .Y(_11373_));
NAND_g _17876_ (.A(_00007_[2]), .B(_11373_), .Y(_11374_));
NAND_g _17877_ (.A(cpuregs[10][7]), .B(_09025_), .Y(_11375_));
NAND_g _17878_ (.A(cpuregs[11][7]), .B(_00007_[0]), .Y(_11376_));
NAND_g _17879_ (.A(_11375_), .B(_11376_), .Y(_11377_));
NAND_g _17880_ (.A(_09027_), .B(_11377_), .Y(_11378_));
NAND_g _17881_ (.A(_11374_), .B(_11378_), .Y(_11379_));
NAND_g _17882_ (.A(_00007_[3]), .B(_11379_), .Y(_11380_));
NAND_g _17883_ (.A(cpuregs[6][7]), .B(_09025_), .Y(_11381_));
NAND_g _17884_ (.A(cpuregs[7][7]), .B(_00007_[0]), .Y(_11382_));
NAND_g _17885_ (.A(_11381_), .B(_11382_), .Y(_11383_));
NAND_g _17886_ (.A(_00007_[2]), .B(_11383_), .Y(_11384_));
NAND_g _17887_ (.A(cpuregs[2][7]), .B(_09025_), .Y(_11385_));
NAND_g _17888_ (.A(cpuregs[3][7]), .B(_00007_[0]), .Y(_11386_));
NAND_g _17889_ (.A(_11385_), .B(_11386_), .Y(_11387_));
NAND_g _17890_ (.A(_09027_), .B(_11387_), .Y(_11388_));
NAND_g _17891_ (.A(_11384_), .B(_11388_), .Y(_11389_));
NAND_g _17892_ (.A(_09028_), .B(_11389_), .Y(_11390_));
AND_g _17893_ (.A(_09029_), .B(_11390_), .Y(_11391_));
NAND_g _17894_ (.A(_11380_), .B(_11391_), .Y(_11392_));
NAND_g _17895_ (.A(cpuregs[27][7]), .B(_09027_), .Y(_11393_));
NAND_g _17896_ (.A(cpuregs[31][7]), .B(_00007_[2]), .Y(_11394_));
AND_g _17897_ (.A(_00007_[0]), .B(_11394_), .Y(_11395_));
NAND_g _17898_ (.A(_11393_), .B(_11395_), .Y(_11396_));
NAND_g _17899_ (.A(cpuregs[26][7]), .B(_09027_), .Y(_11397_));
NAND_g _17900_ (.A(cpuregs[30][7]), .B(_00007_[2]), .Y(_11398_));
AND_g _17901_ (.A(_09025_), .B(_11398_), .Y(_11399_));
NAND_g _17902_ (.A(_11397_), .B(_11399_), .Y(_11400_));
AND_g _17903_ (.A(_00007_[3]), .B(_11400_), .Y(_11401_));
NAND_g _17904_ (.A(_11396_), .B(_11401_), .Y(_11402_));
NAND_g _17905_ (.A(cpuregs[19][7]), .B(_09027_), .Y(_11403_));
NAND_g _17906_ (.A(cpuregs[23][7]), .B(_00007_[2]), .Y(_11404_));
AND_g _17907_ (.A(_00007_[0]), .B(_11404_), .Y(_11405_));
NAND_g _17908_ (.A(_11403_), .B(_11405_), .Y(_11406_));
NAND_g _17909_ (.A(cpuregs[18][7]), .B(_09027_), .Y(_11407_));
NAND_g _17910_ (.A(cpuregs[22][7]), .B(_00007_[2]), .Y(_11408_));
AND_g _17911_ (.A(_09025_), .B(_11408_), .Y(_11409_));
NAND_g _17912_ (.A(_11407_), .B(_11409_), .Y(_11410_));
AND_g _17913_ (.A(_09028_), .B(_11410_), .Y(_11411_));
NAND_g _17914_ (.A(_11406_), .B(_11411_), .Y(_11412_));
AND_g _17915_ (.A(_00007_[4]), .B(_11412_), .Y(_11413_));
NAND_g _17916_ (.A(_11402_), .B(_11413_), .Y(_11414_));
NAND_g _17917_ (.A(_11392_), .B(_11414_), .Y(_11415_));
NAND_g _17918_ (.A(_00007_[1]), .B(_11415_), .Y(_11416_));
NAND_g _17919_ (.A(cpuregs[13][7]), .B(_00007_[2]), .Y(_11417_));
NAND_g _17920_ (.A(cpuregs[9][7]), .B(_09027_), .Y(_11418_));
AND_g _17921_ (.A(_00007_[0]), .B(_11418_), .Y(_11419_));
NAND_g _17922_ (.A(_11417_), .B(_11419_), .Y(_11420_));
NAND_g _17923_ (.A(cpuregs[8][7]), .B(_09027_), .Y(_11421_));
NAND_g _17924_ (.A(cpuregs[12][7]), .B(_00007_[2]), .Y(_11422_));
AND_g _17925_ (.A(_09025_), .B(_11422_), .Y(_11423_));
NAND_g _17926_ (.A(_11421_), .B(_11423_), .Y(_11424_));
AND_g _17927_ (.A(_00007_[3]), .B(_11424_), .Y(_11425_));
NAND_g _17928_ (.A(_11420_), .B(_11425_), .Y(_11426_));
NAND_g _17929_ (.A(cpuregs[1][7]), .B(_09027_), .Y(_11427_));
NAND_g _17930_ (.A(cpuregs[5][7]), .B(_00007_[2]), .Y(_11428_));
AND_g _17931_ (.A(_00007_[0]), .B(_11428_), .Y(_11429_));
NAND_g _17932_ (.A(_11427_), .B(_11429_), .Y(_11430_));
NAND_g _17933_ (.A(cpuregs[0][7]), .B(_09027_), .Y(_11431_));
NAND_g _17934_ (.A(cpuregs[4][7]), .B(_00007_[2]), .Y(_11432_));
AND_g _17935_ (.A(_09025_), .B(_11432_), .Y(_11433_));
NAND_g _17936_ (.A(_11431_), .B(_11433_), .Y(_11434_));
AND_g _17937_ (.A(_09028_), .B(_11434_), .Y(_11435_));
NAND_g _17938_ (.A(_11430_), .B(_11435_), .Y(_11436_));
AND_g _17939_ (.A(_09029_), .B(_11436_), .Y(_11437_));
NAND_g _17940_ (.A(_11426_), .B(_11437_), .Y(_11438_));
NAND_g _17941_ (.A(cpuregs[25][7]), .B(_09027_), .Y(_11439_));
NAND_g _17942_ (.A(cpuregs[29][7]), .B(_00007_[2]), .Y(_11440_));
AND_g _17943_ (.A(_00007_[0]), .B(_11440_), .Y(_11441_));
NAND_g _17944_ (.A(_11439_), .B(_11441_), .Y(_11442_));
NAND_g _17945_ (.A(cpuregs[24][7]), .B(_09027_), .Y(_11443_));
NAND_g _17946_ (.A(cpuregs[28][7]), .B(_00007_[2]), .Y(_11444_));
AND_g _17947_ (.A(_09025_), .B(_11444_), .Y(_11445_));
NAND_g _17948_ (.A(_11443_), .B(_11445_), .Y(_11446_));
AND_g _17949_ (.A(_00007_[3]), .B(_11446_), .Y(_11447_));
NAND_g _17950_ (.A(_11442_), .B(_11447_), .Y(_11448_));
NAND_g _17951_ (.A(cpuregs[21][7]), .B(_00007_[2]), .Y(_11449_));
NAND_g _17952_ (.A(cpuregs[17][7]), .B(_09027_), .Y(_11450_));
AND_g _17953_ (.A(_00007_[0]), .B(_11450_), .Y(_11451_));
NAND_g _17954_ (.A(_11449_), .B(_11451_), .Y(_11452_));
NAND_g _17955_ (.A(cpuregs[20][7]), .B(_00007_[2]), .Y(_11453_));
NAND_g _17956_ (.A(cpuregs[16][7]), .B(_09027_), .Y(_11454_));
AND_g _17957_ (.A(_09025_), .B(_11454_), .Y(_11455_));
NAND_g _17958_ (.A(_11453_), .B(_11455_), .Y(_11456_));
AND_g _17959_ (.A(_09028_), .B(_11456_), .Y(_11457_));
NAND_g _17960_ (.A(_11452_), .B(_11457_), .Y(_11458_));
AND_g _17961_ (.A(_00007_[4]), .B(_11458_), .Y(_11459_));
NAND_g _17962_ (.A(_11448_), .B(_11459_), .Y(_11460_));
NAND_g _17963_ (.A(_11438_), .B(_11460_), .Y(_11461_));
NAND_g _17964_ (.A(_09026_), .B(_11461_), .Y(_11462_));
AND_g _17965_ (.A(_11416_), .B(_11462_), .Y(_11463_));
NAND_g _17966_ (.A(_11170_), .B(_11463_), .Y(_11464_));
NAND_g _17967_ (.A(decoded_imm[7]), .B(_10606_), .Y(_11465_));
AND_g _17968_ (.A(_10603_), .B(_11465_), .Y(_11466_));
NAND_g _17969_ (.A(_11464_), .B(_11466_), .Y(_11467_));
AND_g _17970_ (.A(_11370_), .B(_11467_), .Y(_00282_));
NAND_g _17971_ (.A(_08818_), .B(_10604_), .Y(_11468_));
NAND_g _17972_ (.A(cpuregs[14][8]), .B(_09025_), .Y(_11469_));
NAND_g _17973_ (.A(cpuregs[15][8]), .B(_00007_[0]), .Y(_11470_));
NAND_g _17974_ (.A(_11469_), .B(_11470_), .Y(_11471_));
NAND_g _17975_ (.A(_00007_[2]), .B(_11471_), .Y(_11472_));
NAND_g _17976_ (.A(cpuregs[10][8]), .B(_09025_), .Y(_11473_));
NAND_g _17977_ (.A(cpuregs[11][8]), .B(_00007_[0]), .Y(_11474_));
NAND_g _17978_ (.A(_11473_), .B(_11474_), .Y(_11475_));
NAND_g _17979_ (.A(_09027_), .B(_11475_), .Y(_11476_));
NAND_g _17980_ (.A(_11472_), .B(_11476_), .Y(_11477_));
NAND_g _17981_ (.A(_00007_[3]), .B(_11477_), .Y(_11478_));
NAND_g _17982_ (.A(cpuregs[6][8]), .B(_09025_), .Y(_11479_));
NAND_g _17983_ (.A(cpuregs[7][8]), .B(_00007_[0]), .Y(_11480_));
NAND_g _17984_ (.A(_11479_), .B(_11480_), .Y(_11481_));
NAND_g _17985_ (.A(_00007_[2]), .B(_11481_), .Y(_11482_));
NAND_g _17986_ (.A(cpuregs[2][8]), .B(_09025_), .Y(_11483_));
NAND_g _17987_ (.A(cpuregs[3][8]), .B(_00007_[0]), .Y(_11484_));
NAND_g _17988_ (.A(_11483_), .B(_11484_), .Y(_11485_));
NAND_g _17989_ (.A(_09027_), .B(_11485_), .Y(_11486_));
NAND_g _17990_ (.A(_11482_), .B(_11486_), .Y(_11487_));
NAND_g _17991_ (.A(_09028_), .B(_11487_), .Y(_11488_));
AND_g _17992_ (.A(_09029_), .B(_11488_), .Y(_11489_));
NAND_g _17993_ (.A(_11478_), .B(_11489_), .Y(_11490_));
NAND_g _17994_ (.A(cpuregs[27][8]), .B(_09027_), .Y(_11491_));
NAND_g _17995_ (.A(cpuregs[31][8]), .B(_00007_[2]), .Y(_11492_));
AND_g _17996_ (.A(_00007_[0]), .B(_11492_), .Y(_11493_));
NAND_g _17997_ (.A(_11491_), .B(_11493_), .Y(_11494_));
NAND_g _17998_ (.A(cpuregs[26][8]), .B(_09027_), .Y(_11495_));
NAND_g _17999_ (.A(cpuregs[30][8]), .B(_00007_[2]), .Y(_11496_));
AND_g _18000_ (.A(_09025_), .B(_11496_), .Y(_11497_));
NAND_g _18001_ (.A(_11495_), .B(_11497_), .Y(_11498_));
AND_g _18002_ (.A(_00007_[3]), .B(_11498_), .Y(_11499_));
NAND_g _18003_ (.A(_11494_), .B(_11499_), .Y(_11500_));
NAND_g _18004_ (.A(cpuregs[19][8]), .B(_09027_), .Y(_11501_));
NAND_g _18005_ (.A(cpuregs[23][8]), .B(_00007_[2]), .Y(_11502_));
AND_g _18006_ (.A(_00007_[0]), .B(_11502_), .Y(_11503_));
NAND_g _18007_ (.A(_11501_), .B(_11503_), .Y(_11504_));
NAND_g _18008_ (.A(cpuregs[18][8]), .B(_09027_), .Y(_11505_));
NAND_g _18009_ (.A(cpuregs[22][8]), .B(_00007_[2]), .Y(_11506_));
AND_g _18010_ (.A(_09025_), .B(_11506_), .Y(_11507_));
NAND_g _18011_ (.A(_11505_), .B(_11507_), .Y(_11508_));
AND_g _18012_ (.A(_09028_), .B(_11508_), .Y(_11509_));
NAND_g _18013_ (.A(_11504_), .B(_11509_), .Y(_11510_));
AND_g _18014_ (.A(_00007_[4]), .B(_11510_), .Y(_11511_));
NAND_g _18015_ (.A(_11500_), .B(_11511_), .Y(_11512_));
NAND_g _18016_ (.A(_11490_), .B(_11512_), .Y(_11513_));
NAND_g _18017_ (.A(_00007_[1]), .B(_11513_), .Y(_11514_));
NAND_g _18018_ (.A(cpuregs[13][8]), .B(_00007_[2]), .Y(_11515_));
NAND_g _18019_ (.A(cpuregs[9][8]), .B(_09027_), .Y(_11516_));
AND_g _18020_ (.A(_00007_[0]), .B(_11516_), .Y(_11517_));
NAND_g _18021_ (.A(_11515_), .B(_11517_), .Y(_11518_));
NAND_g _18022_ (.A(cpuregs[8][8]), .B(_09027_), .Y(_11519_));
NAND_g _18023_ (.A(cpuregs[12][8]), .B(_00007_[2]), .Y(_11520_));
AND_g _18024_ (.A(_09025_), .B(_11520_), .Y(_11521_));
NAND_g _18025_ (.A(_11519_), .B(_11521_), .Y(_11522_));
AND_g _18026_ (.A(_00007_[3]), .B(_11522_), .Y(_11523_));
NAND_g _18027_ (.A(_11518_), .B(_11523_), .Y(_11524_));
NAND_g _18028_ (.A(cpuregs[1][8]), .B(_09027_), .Y(_11525_));
NAND_g _18029_ (.A(cpuregs[5][8]), .B(_00007_[2]), .Y(_11526_));
AND_g _18030_ (.A(_00007_[0]), .B(_11526_), .Y(_11527_));
NAND_g _18031_ (.A(_11525_), .B(_11527_), .Y(_11528_));
NAND_g _18032_ (.A(cpuregs[0][8]), .B(_09027_), .Y(_11529_));
NAND_g _18033_ (.A(cpuregs[4][8]), .B(_00007_[2]), .Y(_11530_));
AND_g _18034_ (.A(_09025_), .B(_11530_), .Y(_11531_));
NAND_g _18035_ (.A(_11529_), .B(_11531_), .Y(_11532_));
AND_g _18036_ (.A(_09028_), .B(_11528_), .Y(_11533_));
NAND_g _18037_ (.A(_11532_), .B(_11533_), .Y(_11534_));
AND_g _18038_ (.A(_09029_), .B(_11534_), .Y(_11535_));
NAND_g _18039_ (.A(_11524_), .B(_11535_), .Y(_11536_));
NAND_g _18040_ (.A(cpuregs[25][8]), .B(_09027_), .Y(_11537_));
NAND_g _18041_ (.A(cpuregs[29][8]), .B(_00007_[2]), .Y(_11538_));
AND_g _18042_ (.A(_00007_[0]), .B(_11538_), .Y(_11539_));
NAND_g _18043_ (.A(_11537_), .B(_11539_), .Y(_11540_));
NAND_g _18044_ (.A(cpuregs[24][8]), .B(_09027_), .Y(_11541_));
NAND_g _18045_ (.A(cpuregs[28][8]), .B(_00007_[2]), .Y(_11542_));
AND_g _18046_ (.A(_09025_), .B(_11542_), .Y(_11543_));
NAND_g _18047_ (.A(_11541_), .B(_11543_), .Y(_11544_));
AND_g _18048_ (.A(_00007_[3]), .B(_11544_), .Y(_11545_));
NAND_g _18049_ (.A(_11540_), .B(_11545_), .Y(_11546_));
NAND_g _18050_ (.A(cpuregs[21][8]), .B(_00007_[2]), .Y(_11547_));
NAND_g _18051_ (.A(cpuregs[17][8]), .B(_09027_), .Y(_11548_));
AND_g _18052_ (.A(_00007_[0]), .B(_11548_), .Y(_11549_));
NAND_g _18053_ (.A(_11547_), .B(_11549_), .Y(_11550_));
NAND_g _18054_ (.A(cpuregs[20][8]), .B(_00007_[2]), .Y(_11551_));
NAND_g _18055_ (.A(cpuregs[16][8]), .B(_09027_), .Y(_11552_));
AND_g _18056_ (.A(_09025_), .B(_11552_), .Y(_11553_));
NAND_g _18057_ (.A(_11551_), .B(_11553_), .Y(_11554_));
AND_g _18058_ (.A(_09028_), .B(_11554_), .Y(_11555_));
NAND_g _18059_ (.A(_11550_), .B(_11555_), .Y(_11556_));
AND_g _18060_ (.A(_00007_[4]), .B(_11556_), .Y(_11557_));
NAND_g _18061_ (.A(_11546_), .B(_11557_), .Y(_11558_));
NAND_g _18062_ (.A(_11536_), .B(_11558_), .Y(_11559_));
NAND_g _18063_ (.A(_09026_), .B(_11559_), .Y(_11560_));
AND_g _18064_ (.A(_11514_), .B(_11560_), .Y(_11561_));
NAND_g _18065_ (.A(_11170_), .B(_11561_), .Y(_11562_));
NAND_g _18066_ (.A(decoded_imm[8]), .B(_10606_), .Y(_11563_));
AND_g _18067_ (.A(_10603_), .B(_11563_), .Y(_11564_));
NAND_g _18068_ (.A(_11562_), .B(_11564_), .Y(_11565_));
AND_g _18069_ (.A(_11468_), .B(_11565_), .Y(_00283_));
NAND_g _18070_ (.A(_08819_), .B(_10604_), .Y(_11566_));
NAND_g _18071_ (.A(cpuregs[14][9]), .B(_09025_), .Y(_11567_));
NAND_g _18072_ (.A(cpuregs[15][9]), .B(_00007_[0]), .Y(_11568_));
NAND_g _18073_ (.A(_11567_), .B(_11568_), .Y(_11569_));
NAND_g _18074_ (.A(_00007_[2]), .B(_11569_), .Y(_11570_));
NAND_g _18075_ (.A(cpuregs[10][9]), .B(_09025_), .Y(_11571_));
NAND_g _18076_ (.A(cpuregs[11][9]), .B(_00007_[0]), .Y(_11572_));
NAND_g _18077_ (.A(_11571_), .B(_11572_), .Y(_11573_));
NAND_g _18078_ (.A(_09027_), .B(_11573_), .Y(_11574_));
NAND_g _18079_ (.A(_11570_), .B(_11574_), .Y(_11575_));
NAND_g _18080_ (.A(_00007_[3]), .B(_11575_), .Y(_11576_));
NAND_g _18081_ (.A(cpuregs[6][9]), .B(_09025_), .Y(_11577_));
NAND_g _18082_ (.A(cpuregs[7][9]), .B(_00007_[0]), .Y(_11578_));
NAND_g _18083_ (.A(_11577_), .B(_11578_), .Y(_11579_));
NAND_g _18084_ (.A(_00007_[2]), .B(_11579_), .Y(_11580_));
NAND_g _18085_ (.A(cpuregs[2][9]), .B(_09025_), .Y(_11581_));
NAND_g _18086_ (.A(cpuregs[3][9]), .B(_00007_[0]), .Y(_11582_));
NAND_g _18087_ (.A(_11581_), .B(_11582_), .Y(_11583_));
NAND_g _18088_ (.A(_09027_), .B(_11583_), .Y(_11584_));
NAND_g _18089_ (.A(_11580_), .B(_11584_), .Y(_11585_));
NAND_g _18090_ (.A(_09028_), .B(_11585_), .Y(_11586_));
AND_g _18091_ (.A(_09029_), .B(_11586_), .Y(_11587_));
NAND_g _18092_ (.A(_11576_), .B(_11587_), .Y(_11588_));
NAND_g _18093_ (.A(cpuregs[27][9]), .B(_09027_), .Y(_11589_));
NAND_g _18094_ (.A(cpuregs[31][9]), .B(_00007_[2]), .Y(_11590_));
AND_g _18095_ (.A(_00007_[0]), .B(_11590_), .Y(_11591_));
NAND_g _18096_ (.A(_11589_), .B(_11591_), .Y(_11592_));
NAND_g _18097_ (.A(cpuregs[26][9]), .B(_09027_), .Y(_11593_));
NAND_g _18098_ (.A(cpuregs[30][9]), .B(_00007_[2]), .Y(_11594_));
AND_g _18099_ (.A(_09025_), .B(_11594_), .Y(_11595_));
NAND_g _18100_ (.A(_11593_), .B(_11595_), .Y(_11596_));
AND_g _18101_ (.A(_00007_[3]), .B(_11596_), .Y(_11597_));
NAND_g _18102_ (.A(_11592_), .B(_11597_), .Y(_11598_));
NAND_g _18103_ (.A(cpuregs[19][9]), .B(_09027_), .Y(_11599_));
NAND_g _18104_ (.A(cpuregs[23][9]), .B(_00007_[2]), .Y(_11600_));
AND_g _18105_ (.A(_00007_[0]), .B(_11600_), .Y(_11601_));
NAND_g _18106_ (.A(_11599_), .B(_11601_), .Y(_11602_));
NAND_g _18107_ (.A(cpuregs[18][9]), .B(_09027_), .Y(_11603_));
NAND_g _18108_ (.A(cpuregs[22][9]), .B(_00007_[2]), .Y(_11604_));
AND_g _18109_ (.A(_09025_), .B(_11604_), .Y(_11605_));
NAND_g _18110_ (.A(_11603_), .B(_11605_), .Y(_11606_));
AND_g _18111_ (.A(_09028_), .B(_11606_), .Y(_11607_));
NAND_g _18112_ (.A(_11602_), .B(_11607_), .Y(_11608_));
AND_g _18113_ (.A(_00007_[4]), .B(_11608_), .Y(_11609_));
NAND_g _18114_ (.A(_11598_), .B(_11609_), .Y(_11610_));
NAND_g _18115_ (.A(_11588_), .B(_11610_), .Y(_11611_));
NAND_g _18116_ (.A(_00007_[1]), .B(_11611_), .Y(_11612_));
NAND_g _18117_ (.A(cpuregs[13][9]), .B(_00007_[2]), .Y(_11613_));
NAND_g _18118_ (.A(cpuregs[9][9]), .B(_09027_), .Y(_11614_));
AND_g _18119_ (.A(_00007_[0]), .B(_11614_), .Y(_11615_));
NAND_g _18120_ (.A(_11613_), .B(_11615_), .Y(_11616_));
NAND_g _18121_ (.A(cpuregs[8][9]), .B(_09027_), .Y(_11617_));
NAND_g _18122_ (.A(cpuregs[12][9]), .B(_00007_[2]), .Y(_11618_));
AND_g _18123_ (.A(_09025_), .B(_11618_), .Y(_11619_));
NAND_g _18124_ (.A(_11617_), .B(_11619_), .Y(_11620_));
AND_g _18125_ (.A(_00007_[3]), .B(_11620_), .Y(_11621_));
NAND_g _18126_ (.A(_11616_), .B(_11621_), .Y(_11622_));
NAND_g _18127_ (.A(cpuregs[1][9]), .B(_09027_), .Y(_11623_));
NAND_g _18128_ (.A(cpuregs[5][9]), .B(_00007_[2]), .Y(_11624_));
AND_g _18129_ (.A(_00007_[0]), .B(_11624_), .Y(_11625_));
NAND_g _18130_ (.A(_11623_), .B(_11625_), .Y(_11626_));
NAND_g _18131_ (.A(cpuregs[0][9]), .B(_09027_), .Y(_11627_));
NAND_g _18132_ (.A(cpuregs[4][9]), .B(_00007_[2]), .Y(_11628_));
AND_g _18133_ (.A(_09025_), .B(_11628_), .Y(_11629_));
NAND_g _18134_ (.A(_11627_), .B(_11629_), .Y(_11630_));
AND_g _18135_ (.A(_09028_), .B(_11626_), .Y(_11631_));
NAND_g _18136_ (.A(_11630_), .B(_11631_), .Y(_11632_));
AND_g _18137_ (.A(_09029_), .B(_11632_), .Y(_11633_));
NAND_g _18138_ (.A(_11622_), .B(_11633_), .Y(_11634_));
NAND_g _18139_ (.A(cpuregs[25][9]), .B(_09027_), .Y(_11635_));
NAND_g _18140_ (.A(cpuregs[29][9]), .B(_00007_[2]), .Y(_11636_));
AND_g _18141_ (.A(_00007_[0]), .B(_11636_), .Y(_11637_));
NAND_g _18142_ (.A(_11635_), .B(_11637_), .Y(_11638_));
NAND_g _18143_ (.A(cpuregs[24][9]), .B(_09027_), .Y(_11639_));
NAND_g _18144_ (.A(cpuregs[28][9]), .B(_00007_[2]), .Y(_11640_));
AND_g _18145_ (.A(_09025_), .B(_11640_), .Y(_11641_));
NAND_g _18146_ (.A(_11639_), .B(_11641_), .Y(_11642_));
AND_g _18147_ (.A(_00007_[3]), .B(_11642_), .Y(_11643_));
NAND_g _18148_ (.A(_11638_), .B(_11643_), .Y(_11644_));
NAND_g _18149_ (.A(cpuregs[21][9]), .B(_00007_[2]), .Y(_11645_));
NAND_g _18150_ (.A(cpuregs[17][9]), .B(_09027_), .Y(_11646_));
AND_g _18151_ (.A(_00007_[0]), .B(_11646_), .Y(_11647_));
NAND_g _18152_ (.A(_11645_), .B(_11647_), .Y(_11648_));
NAND_g _18153_ (.A(cpuregs[20][9]), .B(_00007_[2]), .Y(_11649_));
NAND_g _18154_ (.A(cpuregs[16][9]), .B(_09027_), .Y(_11650_));
AND_g _18155_ (.A(_09025_), .B(_11650_), .Y(_11651_));
NAND_g _18156_ (.A(_11649_), .B(_11651_), .Y(_11652_));
AND_g _18157_ (.A(_09028_), .B(_11652_), .Y(_11653_));
NAND_g _18158_ (.A(_11648_), .B(_11653_), .Y(_11654_));
AND_g _18159_ (.A(_00007_[4]), .B(_11654_), .Y(_11655_));
NAND_g _18160_ (.A(_11644_), .B(_11655_), .Y(_11656_));
NAND_g _18161_ (.A(_11634_), .B(_11656_), .Y(_11657_));
NAND_g _18162_ (.A(_09026_), .B(_11657_), .Y(_11658_));
AND_g _18163_ (.A(_11612_), .B(_11658_), .Y(_11659_));
NAND_g _18164_ (.A(_11170_), .B(_11659_), .Y(_11660_));
NAND_g _18165_ (.A(decoded_imm[9]), .B(_10606_), .Y(_11661_));
AND_g _18166_ (.A(_10603_), .B(_11661_), .Y(_11662_));
NAND_g _18167_ (.A(_11660_), .B(_11662_), .Y(_11663_));
AND_g _18168_ (.A(_11566_), .B(_11663_), .Y(_00284_));
NAND_g _18169_ (.A(_08820_), .B(_10604_), .Y(_11664_));
NAND_g _18170_ (.A(cpuregs[9][10]), .B(_09027_), .Y(_11665_));
NAND_g _18171_ (.A(cpuregs[13][10]), .B(_00007_[2]), .Y(_11666_));
NAND_g _18172_ (.A(_11665_), .B(_11666_), .Y(_11667_));
NAND_g _18173_ (.A(_00007_[0]), .B(_11667_), .Y(_11668_));
NAND_g _18174_ (.A(cpuregs[12][10]), .B(_00007_[2]), .Y(_11669_));
NAND_g _18175_ (.A(cpuregs[8][10]), .B(_09027_), .Y(_11670_));
NAND_g _18176_ (.A(_11669_), .B(_11670_), .Y(_11671_));
NAND_g _18177_ (.A(_09025_), .B(_11671_), .Y(_11672_));
NAND_g _18178_ (.A(_11668_), .B(_11672_), .Y(_11673_));
NAND_g _18179_ (.A(_09026_), .B(_11673_), .Y(_11674_));
NAND_g _18180_ (.A(cpuregs[11][10]), .B(_09027_), .Y(_11675_));
NAND_g _18181_ (.A(cpuregs[15][10]), .B(_00007_[2]), .Y(_11676_));
NAND_g _18182_ (.A(_11675_), .B(_11676_), .Y(_11677_));
NAND_g _18183_ (.A(_00007_[0]), .B(_11677_), .Y(_11678_));
NAND_g _18184_ (.A(cpuregs[14][10]), .B(_00007_[2]), .Y(_11679_));
NAND_g _18185_ (.A(cpuregs[10][10]), .B(_09027_), .Y(_11680_));
NAND_g _18186_ (.A(_11679_), .B(_11680_), .Y(_11681_));
NAND_g _18187_ (.A(_09025_), .B(_11681_), .Y(_11682_));
NAND_g _18188_ (.A(_11678_), .B(_11682_), .Y(_11683_));
NAND_g _18189_ (.A(_00007_[1]), .B(_11683_), .Y(_11684_));
NAND_g _18190_ (.A(cpuregs[31][10]), .B(_00007_[2]), .Y(_11685_));
NAND_g _18191_ (.A(cpuregs[27][10]), .B(_09027_), .Y(_11686_));
AND_g _18192_ (.A(_00007_[0]), .B(_11686_), .Y(_11687_));
NAND_g _18193_ (.A(_11685_), .B(_11687_), .Y(_11688_));
NAND_g _18194_ (.A(cpuregs[26][10]), .B(_09027_), .Y(_11689_));
NAND_g _18195_ (.A(cpuregs[30][10]), .B(_00007_[2]), .Y(_11690_));
AND_g _18196_ (.A(_09025_), .B(_11690_), .Y(_11691_));
NAND_g _18197_ (.A(_11689_), .B(_11691_), .Y(_11692_));
AND_g _18198_ (.A(_00007_[1]), .B(_11692_), .Y(_11693_));
NAND_g _18199_ (.A(_11688_), .B(_11693_), .Y(_11694_));
NAND_g _18200_ (.A(cpuregs[29][10]), .B(_00007_[2]), .Y(_11695_));
NAND_g _18201_ (.A(cpuregs[25][10]), .B(_09027_), .Y(_11696_));
AND_g _18202_ (.A(_00007_[0]), .B(_11696_), .Y(_11697_));
NAND_g _18203_ (.A(_11695_), .B(_11697_), .Y(_11698_));
NAND_g _18204_ (.A(cpuregs[24][10]), .B(_09027_), .Y(_11699_));
NAND_g _18205_ (.A(cpuregs[28][10]), .B(_00007_[2]), .Y(_11700_));
AND_g _18206_ (.A(_09025_), .B(_11700_), .Y(_11701_));
NAND_g _18207_ (.A(_11699_), .B(_11701_), .Y(_11702_));
AND_g _18208_ (.A(_09026_), .B(_11702_), .Y(_11703_));
NAND_g _18209_ (.A(_11698_), .B(_11703_), .Y(_11704_));
NAND_g _18210_ (.A(cpuregs[1][10]), .B(_09027_), .Y(_11705_));
NAND_g _18211_ (.A(cpuregs[5][10]), .B(_00007_[2]), .Y(_11706_));
NAND_g _18212_ (.A(_11705_), .B(_11706_), .Y(_11707_));
NAND_g _18213_ (.A(_00007_[0]), .B(_11707_), .Y(_11708_));
NAND_g _18214_ (.A(cpuregs[4][10]), .B(_00007_[2]), .Y(_11709_));
NAND_g _18215_ (.A(cpuregs[0][10]), .B(_09027_), .Y(_11710_));
NAND_g _18216_ (.A(_11709_), .B(_11710_), .Y(_11711_));
NAND_g _18217_ (.A(_09025_), .B(_11711_), .Y(_11712_));
NAND_g _18218_ (.A(_11708_), .B(_11712_), .Y(_11713_));
NAND_g _18219_ (.A(_09026_), .B(_11713_), .Y(_11714_));
NAND_g _18220_ (.A(cpuregs[6][10]), .B(_00007_[2]), .Y(_11715_));
NAND_g _18221_ (.A(cpuregs[2][10]), .B(_09027_), .Y(_11716_));
NAND_g _18222_ (.A(_11715_), .B(_11716_), .Y(_11717_));
NAND_g _18223_ (.A(_09025_), .B(_11717_), .Y(_11718_));
NAND_g _18224_ (.A(cpuregs[7][10]), .B(_00007_[2]), .Y(_11719_));
NAND_g _18225_ (.A(cpuregs[3][10]), .B(_09027_), .Y(_11720_));
NAND_g _18226_ (.A(_11719_), .B(_11720_), .Y(_11721_));
NAND_g _18227_ (.A(_00007_[0]), .B(_11721_), .Y(_11722_));
NAND_g _18228_ (.A(_11718_), .B(_11722_), .Y(_11723_));
NAND_g _18229_ (.A(_00007_[1]), .B(_11723_), .Y(_11724_));
NAND_g _18230_ (.A(_08936_), .B(_09027_), .Y(_11725_));
NOR_g _18231_ (.A(cpuregs[22][10]), .B(_09027_), .Y(_11726_));
NAND_g _18232_ (.A(_08889_), .B(_00007_[2]), .Y(_11727_));
NOR_g _18233_ (.A(cpuregs[19][10]), .B(_00007_[2]), .Y(_11728_));
NOR_g _18234_ (.A(_00007_[0]), .B(_11726_), .Y(_11729_));
AND_g _18235_ (.A(_11725_), .B(_11729_), .Y(_11730_));
NAND_g _18236_ (.A(_00007_[0]), .B(_11727_), .Y(_11731_));
NOR_g _18237_ (.A(_11728_), .B(_11731_), .Y(_11732_));
NOR_g _18238_ (.A(_11730_), .B(_11732_), .Y(_11733_));
NOR_g _18239_ (.A(cpuregs[16][10]), .B(_00007_[2]), .Y(_11734_));
NOR_g _18240_ (.A(cpuregs[20][10]), .B(_09027_), .Y(_11735_));
NOR_g _18241_ (.A(_11734_), .B(_11735_), .Y(_11736_));
NOR_g _18242_ (.A(cpuregs[17][10]), .B(_00007_[2]), .Y(_11737_));
NAND_g _18243_ (.A(_08988_), .B(_00007_[2]), .Y(_11738_));
NAND_g _18244_ (.A(_00007_[0]), .B(_11738_), .Y(_11739_));
NOR_g _18245_ (.A(_11737_), .B(_11739_), .Y(_11740_));
AND_g _18246_ (.A(_09025_), .B(_11736_), .Y(_11741_));
NOR_g _18247_ (.A(_11740_), .B(_11741_), .Y(_11742_));
NAND_g _18248_ (.A(_00007_[1]), .B(_11733_), .Y(_11743_));
NAND_g _18249_ (.A(_09026_), .B(_11742_), .Y(_11744_));
AND_g _18250_ (.A(_09028_), .B(_11744_), .Y(_11745_));
NAND_g _18251_ (.A(_11743_), .B(_11745_), .Y(_11746_));
NAND_g _18252_ (.A(_11694_), .B(_11704_), .Y(_11747_));
NAND_g _18253_ (.A(_00007_[3]), .B(_11747_), .Y(_11748_));
AND_g _18254_ (.A(_00007_[4]), .B(_11748_), .Y(_11749_));
NAND_g _18255_ (.A(_11746_), .B(_11749_), .Y(_11750_));
NAND_g _18256_ (.A(_11714_), .B(_11724_), .Y(_11751_));
NAND_g _18257_ (.A(_09028_), .B(_11751_), .Y(_11752_));
NAND_g _18258_ (.A(_11674_), .B(_11684_), .Y(_11753_));
NAND_g _18259_ (.A(_00007_[3]), .B(_11753_), .Y(_11754_));
AND_g _18260_ (.A(_11752_), .B(_11754_), .Y(_11755_));
NAND_g _18261_ (.A(_09029_), .B(_11755_), .Y(_11756_));
AND_g _18262_ (.A(_11750_), .B(_11756_), .Y(_11757_));
NAND_g _18263_ (.A(_11170_), .B(_11757_), .Y(_11758_));
NAND_g _18264_ (.A(decoded_imm[10]), .B(_10606_), .Y(_11759_));
AND_g _18265_ (.A(_10603_), .B(_11759_), .Y(_11760_));
NAND_g _18266_ (.A(_11758_), .B(_11760_), .Y(_11761_));
AND_g _18267_ (.A(_11664_), .B(_11761_), .Y(_00285_));
NAND_g _18268_ (.A(_08821_), .B(_10604_), .Y(_11762_));
NAND_g _18269_ (.A(cpuregs[9][11]), .B(_09027_), .Y(_11763_));
NAND_g _18270_ (.A(cpuregs[13][11]), .B(_00007_[2]), .Y(_11764_));
NAND_g _18271_ (.A(_11763_), .B(_11764_), .Y(_11765_));
NAND_g _18272_ (.A(_00007_[0]), .B(_11765_), .Y(_11766_));
NAND_g _18273_ (.A(cpuregs[12][11]), .B(_00007_[2]), .Y(_11767_));
NAND_g _18274_ (.A(cpuregs[8][11]), .B(_09027_), .Y(_11768_));
NAND_g _18275_ (.A(_11767_), .B(_11768_), .Y(_11769_));
NAND_g _18276_ (.A(_09025_), .B(_11769_), .Y(_11770_));
NAND_g _18277_ (.A(_11766_), .B(_11770_), .Y(_11771_));
NAND_g _18278_ (.A(_09026_), .B(_11771_), .Y(_11772_));
NAND_g _18279_ (.A(cpuregs[11][11]), .B(_09027_), .Y(_11773_));
NAND_g _18280_ (.A(cpuregs[15][11]), .B(_00007_[2]), .Y(_11774_));
NAND_g _18281_ (.A(_11773_), .B(_11774_), .Y(_11775_));
NAND_g _18282_ (.A(_00007_[0]), .B(_11775_), .Y(_11776_));
NAND_g _18283_ (.A(cpuregs[14][11]), .B(_00007_[2]), .Y(_11777_));
NAND_g _18284_ (.A(cpuregs[10][11]), .B(_09027_), .Y(_11778_));
NAND_g _18285_ (.A(_11777_), .B(_11778_), .Y(_11779_));
NAND_g _18286_ (.A(_09025_), .B(_11779_), .Y(_11780_));
NAND_g _18287_ (.A(_11776_), .B(_11780_), .Y(_11781_));
NAND_g _18288_ (.A(_00007_[1]), .B(_11781_), .Y(_11782_));
NAND_g _18289_ (.A(cpuregs[31][11]), .B(_00007_[2]), .Y(_11783_));
NAND_g _18290_ (.A(cpuregs[27][11]), .B(_09027_), .Y(_11784_));
AND_g _18291_ (.A(_00007_[0]), .B(_11784_), .Y(_11785_));
NAND_g _18292_ (.A(_11783_), .B(_11785_), .Y(_11786_));
NAND_g _18293_ (.A(cpuregs[26][11]), .B(_09027_), .Y(_11787_));
NAND_g _18294_ (.A(cpuregs[30][11]), .B(_00007_[2]), .Y(_11788_));
AND_g _18295_ (.A(_09025_), .B(_11788_), .Y(_11789_));
NAND_g _18296_ (.A(_11787_), .B(_11789_), .Y(_11790_));
AND_g _18297_ (.A(_00007_[1]), .B(_11790_), .Y(_11791_));
NAND_g _18298_ (.A(_11786_), .B(_11791_), .Y(_11792_));
NAND_g _18299_ (.A(cpuregs[29][11]), .B(_00007_[2]), .Y(_11793_));
NAND_g _18300_ (.A(cpuregs[25][11]), .B(_09027_), .Y(_11794_));
AND_g _18301_ (.A(_00007_[0]), .B(_11794_), .Y(_11795_));
NAND_g _18302_ (.A(_11793_), .B(_11795_), .Y(_11796_));
NAND_g _18303_ (.A(cpuregs[24][11]), .B(_09027_), .Y(_11797_));
NAND_g _18304_ (.A(cpuregs[28][11]), .B(_00007_[2]), .Y(_11798_));
AND_g _18305_ (.A(_09025_), .B(_11798_), .Y(_11799_));
NAND_g _18306_ (.A(_11797_), .B(_11799_), .Y(_11800_));
AND_g _18307_ (.A(_09026_), .B(_11800_), .Y(_11801_));
NAND_g _18308_ (.A(_11796_), .B(_11801_), .Y(_11802_));
NAND_g _18309_ (.A(cpuregs[1][11]), .B(_09027_), .Y(_11803_));
NAND_g _18310_ (.A(cpuregs[5][11]), .B(_00007_[2]), .Y(_11804_));
NAND_g _18311_ (.A(_11803_), .B(_11804_), .Y(_11805_));
NAND_g _18312_ (.A(_00007_[0]), .B(_11805_), .Y(_11806_));
NAND_g _18313_ (.A(cpuregs[4][11]), .B(_00007_[2]), .Y(_11807_));
NAND_g _18314_ (.A(cpuregs[0][11]), .B(_09027_), .Y(_11808_));
NAND_g _18315_ (.A(_11807_), .B(_11808_), .Y(_11809_));
NAND_g _18316_ (.A(_09025_), .B(_11809_), .Y(_11810_));
NAND_g _18317_ (.A(_11806_), .B(_11810_), .Y(_11811_));
NAND_g _18318_ (.A(_09026_), .B(_11811_), .Y(_11812_));
NAND_g _18319_ (.A(cpuregs[6][11]), .B(_00007_[2]), .Y(_11813_));
NAND_g _18320_ (.A(cpuregs[2][11]), .B(_09027_), .Y(_11814_));
NAND_g _18321_ (.A(_11813_), .B(_11814_), .Y(_11815_));
NAND_g _18322_ (.A(_09025_), .B(_11815_), .Y(_11816_));
NOR_g _18323_ (.A(cpuregs[3][11]), .B(_00007_[2]), .Y(_11817_));
NAND_g _18324_ (.A(_08967_), .B(_00007_[2]), .Y(_11818_));
NOR_g _18325_ (.A(_09025_), .B(_11817_), .Y(_11819_));
NAND_g _18326_ (.A(_11818_), .B(_11819_), .Y(_11820_));
NAND_g _18327_ (.A(_11816_), .B(_11820_), .Y(_11821_));
NAND_g _18328_ (.A(_00007_[1]), .B(_11821_), .Y(_11822_));
NOR_g _18329_ (.A(cpuregs[18][11]), .B(_00007_[2]), .Y(_11823_));
NAND_g _18330_ (.A(_08919_), .B(_00007_[2]), .Y(_11824_));
NAND_g _18331_ (.A(_08890_), .B(_00007_[2]), .Y(_11825_));
NOR_g _18332_ (.A(cpuregs[19][11]), .B(_00007_[2]), .Y(_11826_));
NAND_g _18333_ (.A(_09025_), .B(_11824_), .Y(_11827_));
NOR_g _18334_ (.A(_11823_), .B(_11827_), .Y(_11828_));
NAND_g _18335_ (.A(_00007_[0]), .B(_11825_), .Y(_11829_));
NOR_g _18336_ (.A(_11826_), .B(_11829_), .Y(_11830_));
NOR_g _18337_ (.A(_11828_), .B(_11830_), .Y(_11831_));
NOR_g _18338_ (.A(cpuregs[16][11]), .B(_00007_[2]), .Y(_11832_));
AND_g _18339_ (.A(_08845_), .B(_00007_[2]), .Y(_11833_));
NOR_g _18340_ (.A(_11832_), .B(_11833_), .Y(_11834_));
NOR_g _18341_ (.A(cpuregs[17][11]), .B(_00007_[2]), .Y(_11835_));
NAND_g _18342_ (.A(_08989_), .B(_00007_[2]), .Y(_11836_));
NAND_g _18343_ (.A(_00007_[0]), .B(_11836_), .Y(_11837_));
NOR_g _18344_ (.A(_11835_), .B(_11837_), .Y(_11838_));
AND_g _18345_ (.A(_09025_), .B(_11834_), .Y(_11839_));
NOR_g _18346_ (.A(_11838_), .B(_11839_), .Y(_11840_));
NAND_g _18347_ (.A(_00007_[1]), .B(_11831_), .Y(_11841_));
NAND_g _18348_ (.A(_09026_), .B(_11840_), .Y(_11842_));
AND_g _18349_ (.A(_11841_), .B(_11842_), .Y(_11843_));
NAND_g _18350_ (.A(_09028_), .B(_11843_), .Y(_11844_));
NAND_g _18351_ (.A(_11792_), .B(_11802_), .Y(_11845_));
NAND_g _18352_ (.A(_00007_[3]), .B(_11845_), .Y(_11846_));
AND_g _18353_ (.A(_00007_[4]), .B(_11846_), .Y(_11847_));
NAND_g _18354_ (.A(_11844_), .B(_11847_), .Y(_11848_));
NAND_g _18355_ (.A(_11772_), .B(_11782_), .Y(_11849_));
NAND_g _18356_ (.A(_00007_[3]), .B(_11849_), .Y(_11850_));
NAND_g _18357_ (.A(_11812_), .B(_11822_), .Y(_11851_));
NAND_g _18358_ (.A(_09028_), .B(_11851_), .Y(_11852_));
AND_g _18359_ (.A(_11850_), .B(_11852_), .Y(_11853_));
NAND_g _18360_ (.A(_09029_), .B(_11853_), .Y(_11854_));
AND_g _18361_ (.A(_11848_), .B(_11854_), .Y(_11855_));
NAND_g _18362_ (.A(_11170_), .B(_11855_), .Y(_11856_));
NAND_g _18363_ (.A(decoded_imm[11]), .B(_10606_), .Y(_11857_));
AND_g _18364_ (.A(_10603_), .B(_11857_), .Y(_11858_));
NAND_g _18365_ (.A(_11856_), .B(_11858_), .Y(_11859_));
AND_g _18366_ (.A(_11762_), .B(_11859_), .Y(_00286_));
NAND_g _18367_ (.A(_08822_), .B(_10604_), .Y(_11860_));
NAND_g _18368_ (.A(_09008_), .B(_00007_[2]), .Y(_11861_));
NOR_g _18369_ (.A(cpuregs[2][12]), .B(_00007_[2]), .Y(_11862_));
NOR_g _18370_ (.A(_00007_[0]), .B(_11862_), .Y(_11863_));
NAND_g _18371_ (.A(_11861_), .B(_11863_), .Y(_11864_));
NAND_g _18372_ (.A(_08968_), .B(_00007_[2]), .Y(_11865_));
NOR_g _18373_ (.A(cpuregs[3][12]), .B(_00007_[2]), .Y(_11866_));
NOR_g _18374_ (.A(_09025_), .B(_11866_), .Y(_11867_));
NAND_g _18375_ (.A(_11865_), .B(_11867_), .Y(_11868_));
NAND_g _18376_ (.A(_11864_), .B(_11868_), .Y(_11869_));
NAND_g _18377_ (.A(_09028_), .B(_11869_), .Y(_11870_));
NAND_g _18378_ (.A(cpuregs[11][12]), .B(_09027_), .Y(_11871_));
NAND_g _18379_ (.A(cpuregs[15][12]), .B(_00007_[2]), .Y(_11872_));
NAND_g _18380_ (.A(_11871_), .B(_11872_), .Y(_11873_));
NAND_g _18381_ (.A(_00007_[0]), .B(_11873_), .Y(_11874_));
NAND_g _18382_ (.A(cpuregs[14][12]), .B(_00007_[2]), .Y(_11875_));
NAND_g _18383_ (.A(cpuregs[10][12]), .B(_09027_), .Y(_11876_));
NAND_g _18384_ (.A(_11875_), .B(_11876_), .Y(_11877_));
NAND_g _18385_ (.A(_09025_), .B(_11877_), .Y(_11878_));
NAND_g _18386_ (.A(_11874_), .B(_11878_), .Y(_11879_));
NAND_g _18387_ (.A(_00007_[3]), .B(_11879_), .Y(_11880_));
AND_g _18388_ (.A(_09029_), .B(_11880_), .Y(_11881_));
NAND_g _18389_ (.A(_11870_), .B(_11881_), .Y(_11882_));
NAND_g _18390_ (.A(cpuregs[31][12]), .B(_00007_[2]), .Y(_11883_));
NAND_g _18391_ (.A(cpuregs[27][12]), .B(_09027_), .Y(_11884_));
AND_g _18392_ (.A(_00007_[0]), .B(_11884_), .Y(_11885_));
NAND_g _18393_ (.A(_11883_), .B(_11885_), .Y(_11886_));
NAND_g _18394_ (.A(cpuregs[26][12]), .B(_09027_), .Y(_11887_));
NAND_g _18395_ (.A(cpuregs[30][12]), .B(_00007_[2]), .Y(_11888_));
AND_g _18396_ (.A(_09025_), .B(_11888_), .Y(_11889_));
NAND_g _18397_ (.A(_11887_), .B(_11889_), .Y(_11890_));
AND_g _18398_ (.A(_00007_[3]), .B(_11890_), .Y(_11891_));
NAND_g _18399_ (.A(_11886_), .B(_11891_), .Y(_11892_));
NOR_g _18400_ (.A(cpuregs[18][12]), .B(_00007_[2]), .Y(_11893_));
NOT_g _18401_ (.A(_11893_), .Y(_11894_));
NAND_g _18402_ (.A(_08920_), .B(_00007_[2]), .Y(_11895_));
NAND_g _18403_ (.A(_11894_), .B(_11895_), .Y(_11896_));
NAND_g _18404_ (.A(_09025_), .B(_11896_), .Y(_11897_));
NAND_g _18405_ (.A(_08891_), .B(_00007_[2]), .Y(_11898_));
NOR_g _18406_ (.A(cpuregs[19][12]), .B(_00007_[2]), .Y(_11899_));
NOT_g _18407_ (.A(_11899_), .Y(_11900_));
NAND_g _18408_ (.A(_11898_), .B(_11900_), .Y(_11901_));
NAND_g _18409_ (.A(_00007_[0]), .B(_11901_), .Y(_11902_));
AND_g _18410_ (.A(_09028_), .B(_11902_), .Y(_11903_));
NAND_g _18411_ (.A(_11897_), .B(_11903_), .Y(_11904_));
AND_g _18412_ (.A(_00007_[4]), .B(_11904_), .Y(_11905_));
NAND_g _18413_ (.A(_11892_), .B(_11905_), .Y(_11906_));
NAND_g _18414_ (.A(_11882_), .B(_11906_), .Y(_11907_));
NAND_g _18415_ (.A(_00007_[1]), .B(_11907_), .Y(_11908_));
NAND_g _18416_ (.A(_08909_), .B(_00007_[2]), .Y(_11909_));
NOR_g _18417_ (.A(cpuregs[0][12]), .B(_00007_[2]), .Y(_11910_));
NOR_g _18418_ (.A(_00007_[0]), .B(_11910_), .Y(_11911_));
NAND_g _18419_ (.A(_11909_), .B(_11911_), .Y(_11912_));
NOR_g _18420_ (.A(cpuregs[1][12]), .B(_00007_[2]), .Y(_11913_));
NOT_g _18421_ (.A(_11913_), .Y(_11914_));
NAND_g _18422_ (.A(_08951_), .B(_00007_[2]), .Y(_11915_));
AND_g _18423_ (.A(_00007_[0]), .B(_11915_), .Y(_11916_));
NAND_g _18424_ (.A(_11914_), .B(_11916_), .Y(_11917_));
NAND_g _18425_ (.A(_11912_), .B(_11917_), .Y(_11918_));
NAND_g _18426_ (.A(_09028_), .B(_11918_), .Y(_11919_));
NAND_g _18427_ (.A(cpuregs[9][12]), .B(_09027_), .Y(_11920_));
NAND_g _18428_ (.A(cpuregs[13][12]), .B(_00007_[2]), .Y(_11921_));
NAND_g _18429_ (.A(_11920_), .B(_11921_), .Y(_11922_));
NAND_g _18430_ (.A(_00007_[0]), .B(_11922_), .Y(_11923_));
NAND_g _18431_ (.A(cpuregs[12][12]), .B(_00007_[2]), .Y(_11924_));
NAND_g _18432_ (.A(cpuregs[8][12]), .B(_09027_), .Y(_11925_));
NAND_g _18433_ (.A(_11924_), .B(_11925_), .Y(_11926_));
NAND_g _18434_ (.A(_09025_), .B(_11926_), .Y(_11927_));
NAND_g _18435_ (.A(_11923_), .B(_11927_), .Y(_11928_));
NAND_g _18436_ (.A(_00007_[3]), .B(_11928_), .Y(_11929_));
AND_g _18437_ (.A(_09029_), .B(_11929_), .Y(_11930_));
NAND_g _18438_ (.A(_11919_), .B(_11930_), .Y(_11931_));
NAND_g _18439_ (.A(cpuregs[29][12]), .B(_00007_[2]), .Y(_11932_));
NAND_g _18440_ (.A(cpuregs[25][12]), .B(_09027_), .Y(_11933_));
AND_g _18441_ (.A(_00007_[0]), .B(_11933_), .Y(_11934_));
NAND_g _18442_ (.A(_11932_), .B(_11934_), .Y(_11935_));
NAND_g _18443_ (.A(cpuregs[24][12]), .B(_09027_), .Y(_11936_));
NAND_g _18444_ (.A(cpuregs[28][12]), .B(_00007_[2]), .Y(_11937_));
AND_g _18445_ (.A(_09025_), .B(_11937_), .Y(_11938_));
NAND_g _18446_ (.A(_11936_), .B(_11938_), .Y(_11939_));
AND_g _18447_ (.A(_00007_[3]), .B(_11939_), .Y(_11940_));
NAND_g _18448_ (.A(_11935_), .B(_11940_), .Y(_11941_));
NOR_g _18449_ (.A(cpuregs[16][12]), .B(_00007_[2]), .Y(_11942_));
NOT_g _18450_ (.A(_11942_), .Y(_11943_));
NAND_g _18451_ (.A(_08846_), .B(_00007_[2]), .Y(_11944_));
NAND_g _18452_ (.A(_11943_), .B(_11944_), .Y(_11945_));
NAND_g _18453_ (.A(_09025_), .B(_11945_), .Y(_11946_));
NAND_g _18454_ (.A(_08942_), .B(_09027_), .Y(_11947_));
NAND_g _18455_ (.A(_08990_), .B(_00007_[2]), .Y(_11948_));
NAND_g _18456_ (.A(_11947_), .B(_11948_), .Y(_11949_));
NAND_g _18457_ (.A(_00007_[0]), .B(_11949_), .Y(_11950_));
AND_g _18458_ (.A(_09028_), .B(_11950_), .Y(_11951_));
NAND_g _18459_ (.A(_11946_), .B(_11951_), .Y(_11952_));
AND_g _18460_ (.A(_00007_[4]), .B(_11952_), .Y(_11953_));
NAND_g _18461_ (.A(_11941_), .B(_11953_), .Y(_11954_));
NAND_g _18462_ (.A(_11931_), .B(_11954_), .Y(_11955_));
NAND_g _18463_ (.A(_09026_), .B(_11955_), .Y(_11956_));
AND_g _18464_ (.A(_11908_), .B(_11956_), .Y(_11957_));
NAND_g _18465_ (.A(_11170_), .B(_11957_), .Y(_11958_));
NAND_g _18466_ (.A(decoded_imm[12]), .B(_10606_), .Y(_11959_));
AND_g _18467_ (.A(_10603_), .B(_11959_), .Y(_11960_));
NAND_g _18468_ (.A(_11958_), .B(_11960_), .Y(_11961_));
AND_g _18469_ (.A(_11860_), .B(_11961_), .Y(_00287_));
NAND_g _18470_ (.A(_08823_), .B(_10604_), .Y(_11962_));
NAND_g _18471_ (.A(cpuregs[14][13]), .B(_09025_), .Y(_11963_));
NAND_g _18472_ (.A(cpuregs[15][13]), .B(_00007_[0]), .Y(_11964_));
NAND_g _18473_ (.A(_11963_), .B(_11964_), .Y(_11965_));
NAND_g _18474_ (.A(_00007_[2]), .B(_11965_), .Y(_11966_));
NAND_g _18475_ (.A(cpuregs[10][13]), .B(_09025_), .Y(_11967_));
NAND_g _18476_ (.A(cpuregs[11][13]), .B(_00007_[0]), .Y(_11968_));
NAND_g _18477_ (.A(_11967_), .B(_11968_), .Y(_11969_));
NAND_g _18478_ (.A(_09027_), .B(_11969_), .Y(_11970_));
NAND_g _18479_ (.A(_11966_), .B(_11970_), .Y(_11971_));
NAND_g _18480_ (.A(_00007_[3]), .B(_11971_), .Y(_11972_));
NAND_g _18481_ (.A(cpuregs[6][13]), .B(_09025_), .Y(_11973_));
NAND_g _18482_ (.A(cpuregs[7][13]), .B(_00007_[0]), .Y(_11974_));
NAND_g _18483_ (.A(_11973_), .B(_11974_), .Y(_11975_));
NAND_g _18484_ (.A(_00007_[2]), .B(_11975_), .Y(_11976_));
NAND_g _18485_ (.A(cpuregs[2][13]), .B(_09025_), .Y(_11977_));
NAND_g _18486_ (.A(cpuregs[3][13]), .B(_00007_[0]), .Y(_11978_));
NAND_g _18487_ (.A(_11977_), .B(_11978_), .Y(_11979_));
NAND_g _18488_ (.A(_09027_), .B(_11979_), .Y(_11980_));
NAND_g _18489_ (.A(_11976_), .B(_11980_), .Y(_11981_));
NAND_g _18490_ (.A(_09028_), .B(_11981_), .Y(_11982_));
AND_g _18491_ (.A(_09029_), .B(_11982_), .Y(_11983_));
NAND_g _18492_ (.A(_11972_), .B(_11983_), .Y(_11984_));
NAND_g _18493_ (.A(cpuregs[27][13]), .B(_09027_), .Y(_11985_));
NAND_g _18494_ (.A(cpuregs[31][13]), .B(_00007_[2]), .Y(_11986_));
AND_g _18495_ (.A(_00007_[0]), .B(_11986_), .Y(_11987_));
NAND_g _18496_ (.A(_11985_), .B(_11987_), .Y(_11988_));
NAND_g _18497_ (.A(cpuregs[26][13]), .B(_09027_), .Y(_11989_));
NAND_g _18498_ (.A(cpuregs[30][13]), .B(_00007_[2]), .Y(_11990_));
AND_g _18499_ (.A(_09025_), .B(_11990_), .Y(_11991_));
NAND_g _18500_ (.A(_11989_), .B(_11991_), .Y(_11992_));
AND_g _18501_ (.A(_00007_[3]), .B(_11992_), .Y(_11993_));
NAND_g _18502_ (.A(_11988_), .B(_11993_), .Y(_11994_));
NAND_g _18503_ (.A(cpuregs[19][13]), .B(_09027_), .Y(_11995_));
NAND_g _18504_ (.A(cpuregs[23][13]), .B(_00007_[2]), .Y(_11996_));
AND_g _18505_ (.A(_00007_[0]), .B(_11996_), .Y(_11997_));
NAND_g _18506_ (.A(_11995_), .B(_11997_), .Y(_11998_));
NAND_g _18507_ (.A(cpuregs[18][13]), .B(_09027_), .Y(_11999_));
NAND_g _18508_ (.A(cpuregs[22][13]), .B(_00007_[2]), .Y(_12000_));
AND_g _18509_ (.A(_09025_), .B(_12000_), .Y(_12001_));
NAND_g _18510_ (.A(_11999_), .B(_12001_), .Y(_12002_));
AND_g _18511_ (.A(_09028_), .B(_12002_), .Y(_12003_));
NAND_g _18512_ (.A(_11998_), .B(_12003_), .Y(_12004_));
AND_g _18513_ (.A(_00007_[4]), .B(_12004_), .Y(_12005_));
NAND_g _18514_ (.A(_11994_), .B(_12005_), .Y(_12006_));
NAND_g _18515_ (.A(_11984_), .B(_12006_), .Y(_12007_));
NAND_g _18516_ (.A(_00007_[1]), .B(_12007_), .Y(_12008_));
NAND_g _18517_ (.A(cpuregs[13][13]), .B(_00007_[2]), .Y(_12009_));
NAND_g _18518_ (.A(cpuregs[9][13]), .B(_09027_), .Y(_12010_));
AND_g _18519_ (.A(_00007_[0]), .B(_12010_), .Y(_12011_));
NAND_g _18520_ (.A(_12009_), .B(_12011_), .Y(_12012_));
NAND_g _18521_ (.A(cpuregs[8][13]), .B(_09027_), .Y(_12013_));
NAND_g _18522_ (.A(cpuregs[12][13]), .B(_00007_[2]), .Y(_12014_));
AND_g _18523_ (.A(_09025_), .B(_12014_), .Y(_12015_));
NAND_g _18524_ (.A(_12013_), .B(_12015_), .Y(_12016_));
AND_g _18525_ (.A(_00007_[3]), .B(_12016_), .Y(_12017_));
NAND_g _18526_ (.A(_12012_), .B(_12017_), .Y(_12018_));
NAND_g _18527_ (.A(cpuregs[1][13]), .B(_09027_), .Y(_12019_));
NAND_g _18528_ (.A(cpuregs[5][13]), .B(_00007_[2]), .Y(_12020_));
AND_g _18529_ (.A(_00007_[0]), .B(_12020_), .Y(_12021_));
NAND_g _18530_ (.A(_12019_), .B(_12021_), .Y(_12022_));
NAND_g _18531_ (.A(cpuregs[0][13]), .B(_09027_), .Y(_12023_));
NAND_g _18532_ (.A(cpuregs[4][13]), .B(_00007_[2]), .Y(_12024_));
AND_g _18533_ (.A(_09025_), .B(_12024_), .Y(_12025_));
NAND_g _18534_ (.A(_12023_), .B(_12025_), .Y(_12026_));
AND_g _18535_ (.A(_09028_), .B(_12026_), .Y(_12027_));
NAND_g _18536_ (.A(_12022_), .B(_12027_), .Y(_12028_));
AND_g _18537_ (.A(_09029_), .B(_12028_), .Y(_12029_));
NAND_g _18538_ (.A(_12018_), .B(_12029_), .Y(_12030_));
NAND_g _18539_ (.A(cpuregs[25][13]), .B(_09027_), .Y(_12031_));
NAND_g _18540_ (.A(cpuregs[29][13]), .B(_00007_[2]), .Y(_12032_));
AND_g _18541_ (.A(_00007_[0]), .B(_12032_), .Y(_12033_));
NAND_g _18542_ (.A(_12031_), .B(_12033_), .Y(_12034_));
NAND_g _18543_ (.A(cpuregs[24][13]), .B(_09027_), .Y(_12035_));
NAND_g _18544_ (.A(cpuregs[28][13]), .B(_00007_[2]), .Y(_12036_));
AND_g _18545_ (.A(_09025_), .B(_12036_), .Y(_12037_));
NAND_g _18546_ (.A(_12035_), .B(_12037_), .Y(_12038_));
AND_g _18547_ (.A(_00007_[3]), .B(_12038_), .Y(_12039_));
NAND_g _18548_ (.A(_12034_), .B(_12039_), .Y(_12040_));
NAND_g _18549_ (.A(cpuregs[21][13]), .B(_00007_[2]), .Y(_12041_));
NAND_g _18550_ (.A(cpuregs[17][13]), .B(_09027_), .Y(_12042_));
AND_g _18551_ (.A(_00007_[0]), .B(_12042_), .Y(_12043_));
NAND_g _18552_ (.A(_12041_), .B(_12043_), .Y(_12044_));
NAND_g _18553_ (.A(cpuregs[20][13]), .B(_00007_[2]), .Y(_12045_));
NAND_g _18554_ (.A(cpuregs[16][13]), .B(_09027_), .Y(_12046_));
AND_g _18555_ (.A(_09025_), .B(_12046_), .Y(_12047_));
NAND_g _18556_ (.A(_12045_), .B(_12047_), .Y(_12048_));
AND_g _18557_ (.A(_09028_), .B(_12048_), .Y(_12049_));
NAND_g _18558_ (.A(_12044_), .B(_12049_), .Y(_12050_));
AND_g _18559_ (.A(_00007_[4]), .B(_12050_), .Y(_12051_));
NAND_g _18560_ (.A(_12040_), .B(_12051_), .Y(_12052_));
NAND_g _18561_ (.A(_12030_), .B(_12052_), .Y(_12053_));
NAND_g _18562_ (.A(_09026_), .B(_12053_), .Y(_12054_));
AND_g _18563_ (.A(_12008_), .B(_12054_), .Y(_12055_));
NAND_g _18564_ (.A(_11170_), .B(_12055_), .Y(_12056_));
NAND_g _18565_ (.A(decoded_imm[13]), .B(_10606_), .Y(_12057_));
AND_g _18566_ (.A(_10603_), .B(_12057_), .Y(_12058_));
NAND_g _18567_ (.A(_12056_), .B(_12058_), .Y(_12059_));
AND_g _18568_ (.A(_11962_), .B(_12059_), .Y(_00288_));
NAND_g _18569_ (.A(_08824_), .B(_10604_), .Y(_12060_));
NAND_g _18570_ (.A(_09009_), .B(_00007_[2]), .Y(_12061_));
NOR_g _18571_ (.A(cpuregs[2][14]), .B(_00007_[2]), .Y(_12062_));
NOR_g _18572_ (.A(_00007_[0]), .B(_12062_), .Y(_12063_));
NAND_g _18573_ (.A(_12061_), .B(_12063_), .Y(_12064_));
NAND_g _18574_ (.A(_08969_), .B(_00007_[2]), .Y(_12065_));
NOR_g _18575_ (.A(cpuregs[3][14]), .B(_00007_[2]), .Y(_12066_));
NOR_g _18576_ (.A(_09025_), .B(_12066_), .Y(_12067_));
NAND_g _18577_ (.A(_12065_), .B(_12067_), .Y(_12068_));
NAND_g _18578_ (.A(_12064_), .B(_12068_), .Y(_12069_));
NAND_g _18579_ (.A(_09028_), .B(_12069_), .Y(_12070_));
NAND_g _18580_ (.A(cpuregs[11][14]), .B(_09027_), .Y(_12071_));
NAND_g _18581_ (.A(cpuregs[15][14]), .B(_00007_[2]), .Y(_12072_));
NAND_g _18582_ (.A(_12071_), .B(_12072_), .Y(_12073_));
NAND_g _18583_ (.A(_00007_[0]), .B(_12073_), .Y(_12074_));
NAND_g _18584_ (.A(cpuregs[14][14]), .B(_00007_[2]), .Y(_12075_));
NAND_g _18585_ (.A(cpuregs[10][14]), .B(_09027_), .Y(_12076_));
NAND_g _18586_ (.A(_12075_), .B(_12076_), .Y(_12077_));
NAND_g _18587_ (.A(_09025_), .B(_12077_), .Y(_12078_));
NAND_g _18588_ (.A(_12074_), .B(_12078_), .Y(_12079_));
NAND_g _18589_ (.A(_00007_[3]), .B(_12079_), .Y(_12080_));
AND_g _18590_ (.A(_09029_), .B(_12080_), .Y(_12081_));
NAND_g _18591_ (.A(_12070_), .B(_12081_), .Y(_12082_));
NAND_g _18592_ (.A(cpuregs[31][14]), .B(_00007_[2]), .Y(_12083_));
NAND_g _18593_ (.A(cpuregs[27][14]), .B(_09027_), .Y(_12084_));
AND_g _18594_ (.A(_00007_[0]), .B(_12084_), .Y(_12085_));
NAND_g _18595_ (.A(_12083_), .B(_12085_), .Y(_12086_));
NAND_g _18596_ (.A(cpuregs[26][14]), .B(_09027_), .Y(_12087_));
NAND_g _18597_ (.A(cpuregs[30][14]), .B(_00007_[2]), .Y(_12088_));
AND_g _18598_ (.A(_09025_), .B(_12088_), .Y(_12089_));
NAND_g _18599_ (.A(_12087_), .B(_12089_), .Y(_12090_));
AND_g _18600_ (.A(_00007_[3]), .B(_12090_), .Y(_12091_));
NAND_g _18601_ (.A(_12086_), .B(_12091_), .Y(_12092_));
NOR_g _18602_ (.A(cpuregs[18][14]), .B(_00007_[2]), .Y(_12093_));
NOT_g _18603_ (.A(_12093_), .Y(_12094_));
NAND_g _18604_ (.A(_08921_), .B(_00007_[2]), .Y(_12095_));
NAND_g _18605_ (.A(_12094_), .B(_12095_), .Y(_12096_));
NAND_g _18606_ (.A(_09025_), .B(_12096_), .Y(_12097_));
NAND_g _18607_ (.A(_08892_), .B(_00007_[2]), .Y(_12098_));
NOR_g _18608_ (.A(cpuregs[19][14]), .B(_00007_[2]), .Y(_12099_));
NOT_g _18609_ (.A(_12099_), .Y(_12100_));
NAND_g _18610_ (.A(_12098_), .B(_12100_), .Y(_12101_));
NAND_g _18611_ (.A(_00007_[0]), .B(_12101_), .Y(_12102_));
AND_g _18612_ (.A(_09028_), .B(_12102_), .Y(_12103_));
NAND_g _18613_ (.A(_12097_), .B(_12103_), .Y(_12104_));
AND_g _18614_ (.A(_00007_[4]), .B(_12104_), .Y(_12105_));
NAND_g _18615_ (.A(_12092_), .B(_12105_), .Y(_12106_));
NAND_g _18616_ (.A(_12082_), .B(_12106_), .Y(_12107_));
NAND_g _18617_ (.A(_00007_[1]), .B(_12107_), .Y(_12108_));
NAND_g _18618_ (.A(_08910_), .B(_00007_[2]), .Y(_12109_));
NOR_g _18619_ (.A(cpuregs[0][14]), .B(_00007_[2]), .Y(_12110_));
NOR_g _18620_ (.A(_00007_[0]), .B(_12110_), .Y(_12111_));
NAND_g _18621_ (.A(_12109_), .B(_12111_), .Y(_12112_));
NOR_g _18622_ (.A(cpuregs[1][14]), .B(_00007_[2]), .Y(_12113_));
NOT_g _18623_ (.A(_12113_), .Y(_12114_));
NAND_g _18624_ (.A(_08952_), .B(_00007_[2]), .Y(_12115_));
AND_g _18625_ (.A(_00007_[0]), .B(_12115_), .Y(_12116_));
NAND_g _18626_ (.A(_12114_), .B(_12116_), .Y(_12117_));
NAND_g _18627_ (.A(_12112_), .B(_12117_), .Y(_12118_));
NAND_g _18628_ (.A(_09028_), .B(_12118_), .Y(_12119_));
NAND_g _18629_ (.A(cpuregs[9][14]), .B(_09027_), .Y(_12120_));
NAND_g _18630_ (.A(cpuregs[13][14]), .B(_00007_[2]), .Y(_12121_));
NAND_g _18631_ (.A(_12120_), .B(_12121_), .Y(_12122_));
NAND_g _18632_ (.A(_00007_[0]), .B(_12122_), .Y(_12123_));
NAND_g _18633_ (.A(cpuregs[12][14]), .B(_00007_[2]), .Y(_12124_));
NAND_g _18634_ (.A(cpuregs[8][14]), .B(_09027_), .Y(_12125_));
NAND_g _18635_ (.A(_12124_), .B(_12125_), .Y(_12126_));
NAND_g _18636_ (.A(_09025_), .B(_12126_), .Y(_12127_));
NAND_g _18637_ (.A(_12123_), .B(_12127_), .Y(_12128_));
NAND_g _18638_ (.A(_00007_[3]), .B(_12128_), .Y(_12129_));
AND_g _18639_ (.A(_09029_), .B(_12129_), .Y(_12130_));
NAND_g _18640_ (.A(_12119_), .B(_12130_), .Y(_12131_));
NAND_g _18641_ (.A(cpuregs[29][14]), .B(_00007_[2]), .Y(_12132_));
NAND_g _18642_ (.A(cpuregs[25][14]), .B(_09027_), .Y(_12133_));
AND_g _18643_ (.A(_00007_[0]), .B(_12133_), .Y(_12134_));
NAND_g _18644_ (.A(_12132_), .B(_12134_), .Y(_12135_));
NAND_g _18645_ (.A(cpuregs[24][14]), .B(_09027_), .Y(_12136_));
NAND_g _18646_ (.A(cpuregs[28][14]), .B(_00007_[2]), .Y(_12137_));
AND_g _18647_ (.A(_09025_), .B(_12137_), .Y(_12138_));
NAND_g _18648_ (.A(_12136_), .B(_12138_), .Y(_12139_));
AND_g _18649_ (.A(_00007_[3]), .B(_12139_), .Y(_12140_));
NAND_g _18650_ (.A(_12135_), .B(_12140_), .Y(_12141_));
NOR_g _18651_ (.A(cpuregs[16][14]), .B(_00007_[2]), .Y(_12142_));
NOT_g _18652_ (.A(_12142_), .Y(_12143_));
NAND_g _18653_ (.A(_08847_), .B(_00007_[2]), .Y(_12144_));
NAND_g _18654_ (.A(_12143_), .B(_12144_), .Y(_12145_));
NAND_g _18655_ (.A(_09025_), .B(_12145_), .Y(_12146_));
NAND_g _18656_ (.A(_08943_), .B(_09027_), .Y(_12147_));
NAND_g _18657_ (.A(_08991_), .B(_00007_[2]), .Y(_12148_));
NAND_g _18658_ (.A(_12147_), .B(_12148_), .Y(_12149_));
NAND_g _18659_ (.A(_00007_[0]), .B(_12149_), .Y(_12150_));
AND_g _18660_ (.A(_09028_), .B(_12150_), .Y(_12151_));
NAND_g _18661_ (.A(_12146_), .B(_12151_), .Y(_12152_));
AND_g _18662_ (.A(_00007_[4]), .B(_12152_), .Y(_12153_));
NAND_g _18663_ (.A(_12141_), .B(_12153_), .Y(_12154_));
NAND_g _18664_ (.A(_12131_), .B(_12154_), .Y(_12155_));
NAND_g _18665_ (.A(_09026_), .B(_12155_), .Y(_12156_));
AND_g _18666_ (.A(_12108_), .B(_12156_), .Y(_12157_));
NAND_g _18667_ (.A(_11170_), .B(_12157_), .Y(_12158_));
NAND_g _18668_ (.A(decoded_imm[14]), .B(_10606_), .Y(_12159_));
AND_g _18669_ (.A(_10603_), .B(_12159_), .Y(_12160_));
NAND_g _18670_ (.A(_12158_), .B(_12160_), .Y(_12161_));
AND_g _18671_ (.A(_12060_), .B(_12161_), .Y(_00289_));
NAND_g _18672_ (.A(_08825_), .B(_10604_), .Y(_12162_));
NAND_g _18673_ (.A(cpuregs[9][15]), .B(_09027_), .Y(_12163_));
NAND_g _18674_ (.A(cpuregs[13][15]), .B(_00007_[2]), .Y(_12164_));
NAND_g _18675_ (.A(_12163_), .B(_12164_), .Y(_12165_));
NAND_g _18676_ (.A(_00007_[0]), .B(_12165_), .Y(_12166_));
NAND_g _18677_ (.A(cpuregs[12][15]), .B(_00007_[2]), .Y(_12167_));
NAND_g _18678_ (.A(cpuregs[8][15]), .B(_09027_), .Y(_12168_));
NAND_g _18679_ (.A(_12167_), .B(_12168_), .Y(_12169_));
NAND_g _18680_ (.A(_09025_), .B(_12169_), .Y(_12170_));
NAND_g _18681_ (.A(_12166_), .B(_12170_), .Y(_12171_));
NAND_g _18682_ (.A(_09026_), .B(_12171_), .Y(_12172_));
NAND_g _18683_ (.A(cpuregs[11][15]), .B(_09027_), .Y(_12173_));
NAND_g _18684_ (.A(cpuregs[15][15]), .B(_00007_[2]), .Y(_12174_));
NAND_g _18685_ (.A(_12173_), .B(_12174_), .Y(_12175_));
NAND_g _18686_ (.A(_00007_[0]), .B(_12175_), .Y(_12176_));
NAND_g _18687_ (.A(cpuregs[14][15]), .B(_00007_[2]), .Y(_12177_));
NAND_g _18688_ (.A(cpuregs[10][15]), .B(_09027_), .Y(_12178_));
NAND_g _18689_ (.A(_12177_), .B(_12178_), .Y(_12179_));
NAND_g _18690_ (.A(_09025_), .B(_12179_), .Y(_12180_));
NAND_g _18691_ (.A(_12176_), .B(_12180_), .Y(_12181_));
NAND_g _18692_ (.A(_00007_[1]), .B(_12181_), .Y(_12182_));
NAND_g _18693_ (.A(cpuregs[31][15]), .B(_00007_[2]), .Y(_12183_));
NAND_g _18694_ (.A(cpuregs[27][15]), .B(_09027_), .Y(_12184_));
AND_g _18695_ (.A(_00007_[0]), .B(_12184_), .Y(_12185_));
NAND_g _18696_ (.A(_12183_), .B(_12185_), .Y(_12186_));
NAND_g _18697_ (.A(cpuregs[26][15]), .B(_09027_), .Y(_12187_));
NAND_g _18698_ (.A(cpuregs[30][15]), .B(_00007_[2]), .Y(_12188_));
AND_g _18699_ (.A(_09025_), .B(_12188_), .Y(_12189_));
NAND_g _18700_ (.A(_12187_), .B(_12189_), .Y(_12190_));
AND_g _18701_ (.A(_00007_[1]), .B(_12190_), .Y(_12191_));
NAND_g _18702_ (.A(_12186_), .B(_12191_), .Y(_12192_));
NAND_g _18703_ (.A(cpuregs[29][15]), .B(_00007_[2]), .Y(_12193_));
NAND_g _18704_ (.A(cpuregs[25][15]), .B(_09027_), .Y(_12194_));
AND_g _18705_ (.A(_00007_[0]), .B(_12194_), .Y(_12195_));
NAND_g _18706_ (.A(_12193_), .B(_12195_), .Y(_12196_));
NAND_g _18707_ (.A(cpuregs[24][15]), .B(_09027_), .Y(_12197_));
NAND_g _18708_ (.A(cpuregs[28][15]), .B(_00007_[2]), .Y(_12198_));
AND_g _18709_ (.A(_09025_), .B(_12198_), .Y(_12199_));
NAND_g _18710_ (.A(_12197_), .B(_12199_), .Y(_12200_));
AND_g _18711_ (.A(_09026_), .B(_12200_), .Y(_12201_));
NAND_g _18712_ (.A(_12196_), .B(_12201_), .Y(_12202_));
NAND_g _18713_ (.A(cpuregs[1][15]), .B(_09027_), .Y(_12203_));
NAND_g _18714_ (.A(cpuregs[5][15]), .B(_00007_[2]), .Y(_12204_));
NAND_g _18715_ (.A(_12203_), .B(_12204_), .Y(_12205_));
NAND_g _18716_ (.A(_00007_[0]), .B(_12205_), .Y(_12206_));
NAND_g _18717_ (.A(cpuregs[4][15]), .B(_00007_[2]), .Y(_12207_));
NAND_g _18718_ (.A(cpuregs[0][15]), .B(_09027_), .Y(_12208_));
NAND_g _18719_ (.A(_12207_), .B(_12208_), .Y(_12209_));
NAND_g _18720_ (.A(_09025_), .B(_12209_), .Y(_12210_));
NAND_g _18721_ (.A(_12206_), .B(_12210_), .Y(_12211_));
NAND_g _18722_ (.A(_09026_), .B(_12211_), .Y(_12212_));
NAND_g _18723_ (.A(cpuregs[6][15]), .B(_00007_[2]), .Y(_12213_));
NAND_g _18724_ (.A(cpuregs[2][15]), .B(_09027_), .Y(_12214_));
NAND_g _18725_ (.A(_12213_), .B(_12214_), .Y(_12215_));
NAND_g _18726_ (.A(_09025_), .B(_12215_), .Y(_12216_));
NOR_g _18727_ (.A(cpuregs[3][15]), .B(_00007_[2]), .Y(_12217_));
NAND_g _18728_ (.A(_08970_), .B(_00007_[2]), .Y(_12218_));
NOR_g _18729_ (.A(_09025_), .B(_12217_), .Y(_12219_));
NAND_g _18730_ (.A(_12218_), .B(_12219_), .Y(_12220_));
NAND_g _18731_ (.A(_12216_), .B(_12220_), .Y(_12221_));
NAND_g _18732_ (.A(_00007_[1]), .B(_12221_), .Y(_12222_));
NOR_g _18733_ (.A(cpuregs[18][15]), .B(_00007_[2]), .Y(_12223_));
NAND_g _18734_ (.A(_08922_), .B(_00007_[2]), .Y(_12224_));
NAND_g _18735_ (.A(_08893_), .B(_00007_[2]), .Y(_12225_));
NOR_g _18736_ (.A(cpuregs[19][15]), .B(_00007_[2]), .Y(_12226_));
NAND_g _18737_ (.A(_09025_), .B(_12224_), .Y(_12227_));
NOR_g _18738_ (.A(_12223_), .B(_12227_), .Y(_12228_));
NAND_g _18739_ (.A(_00007_[0]), .B(_12225_), .Y(_12229_));
NOR_g _18740_ (.A(_12226_), .B(_12229_), .Y(_12230_));
NOR_g _18741_ (.A(_12228_), .B(_12230_), .Y(_12231_));
NOR_g _18742_ (.A(cpuregs[16][15]), .B(_00007_[2]), .Y(_12232_));
AND_g _18743_ (.A(_08848_), .B(_00007_[2]), .Y(_12233_));
NOR_g _18744_ (.A(_12232_), .B(_12233_), .Y(_12234_));
NOR_g _18745_ (.A(cpuregs[17][15]), .B(_00007_[2]), .Y(_12235_));
NAND_g _18746_ (.A(_08992_), .B(_00007_[2]), .Y(_12236_));
NAND_g _18747_ (.A(_00007_[0]), .B(_12236_), .Y(_12237_));
NOR_g _18748_ (.A(_12235_), .B(_12237_), .Y(_12238_));
AND_g _18749_ (.A(_09025_), .B(_12234_), .Y(_12239_));
NOR_g _18750_ (.A(_12238_), .B(_12239_), .Y(_12240_));
NAND_g _18751_ (.A(_00007_[1]), .B(_12231_), .Y(_12241_));
NAND_g _18752_ (.A(_09026_), .B(_12240_), .Y(_12242_));
AND_g _18753_ (.A(_09028_), .B(_12242_), .Y(_12243_));
NAND_g _18754_ (.A(_12241_), .B(_12243_), .Y(_12244_));
NAND_g _18755_ (.A(_12192_), .B(_12202_), .Y(_12245_));
NAND_g _18756_ (.A(_00007_[3]), .B(_12245_), .Y(_12246_));
AND_g _18757_ (.A(_00007_[4]), .B(_12246_), .Y(_12247_));
NAND_g _18758_ (.A(_12244_), .B(_12247_), .Y(_12248_));
NAND_g _18759_ (.A(_12172_), .B(_12182_), .Y(_12249_));
NAND_g _18760_ (.A(_00007_[3]), .B(_12249_), .Y(_12250_));
NAND_g _18761_ (.A(_12212_), .B(_12222_), .Y(_12251_));
NAND_g _18762_ (.A(_09028_), .B(_12251_), .Y(_12252_));
AND_g _18763_ (.A(_12250_), .B(_12252_), .Y(_12253_));
NAND_g _18764_ (.A(_09029_), .B(_12253_), .Y(_12254_));
AND_g _18765_ (.A(_12248_), .B(_12254_), .Y(_12255_));
NAND_g _18766_ (.A(_11170_), .B(_12255_), .Y(_12256_));
NAND_g _18767_ (.A(decoded_imm[15]), .B(_10606_), .Y(_12257_));
AND_g _18768_ (.A(_10603_), .B(_12257_), .Y(_12258_));
NAND_g _18769_ (.A(_12256_), .B(_12258_), .Y(_12259_));
AND_g _18770_ (.A(_12162_), .B(_12259_), .Y(_00290_));
NAND_g _18771_ (.A(_08826_), .B(_10604_), .Y(_12260_));
NAND_g _18772_ (.A(_09011_), .B(_00007_[2]), .Y(_12261_));
NOR_g _18773_ (.A(cpuregs[2][16]), .B(_00007_[2]), .Y(_12262_));
NOR_g _18774_ (.A(_00007_[0]), .B(_12262_), .Y(_12263_));
NAND_g _18775_ (.A(_12261_), .B(_12263_), .Y(_12264_));
NAND_g _18776_ (.A(_08971_), .B(_00007_[2]), .Y(_12265_));
NOR_g _18777_ (.A(cpuregs[3][16]), .B(_00007_[2]), .Y(_12266_));
NOR_g _18778_ (.A(_09025_), .B(_12266_), .Y(_12267_));
NAND_g _18779_ (.A(_12265_), .B(_12267_), .Y(_12268_));
NAND_g _18780_ (.A(_12264_), .B(_12268_), .Y(_12269_));
NAND_g _18781_ (.A(_09028_), .B(_12269_), .Y(_12270_));
NAND_g _18782_ (.A(cpuregs[11][16]), .B(_09027_), .Y(_12271_));
NAND_g _18783_ (.A(cpuregs[15][16]), .B(_00007_[2]), .Y(_12272_));
NAND_g _18784_ (.A(_12271_), .B(_12272_), .Y(_12273_));
NAND_g _18785_ (.A(_00007_[0]), .B(_12273_), .Y(_12274_));
NAND_g _18786_ (.A(cpuregs[14][16]), .B(_00007_[2]), .Y(_12275_));
NAND_g _18787_ (.A(cpuregs[10][16]), .B(_09027_), .Y(_12276_));
NAND_g _18788_ (.A(_12275_), .B(_12276_), .Y(_12277_));
NAND_g _18789_ (.A(_09025_), .B(_12277_), .Y(_12278_));
NAND_g _18790_ (.A(_12274_), .B(_12278_), .Y(_12279_));
NAND_g _18791_ (.A(_00007_[3]), .B(_12279_), .Y(_12280_));
AND_g _18792_ (.A(_09029_), .B(_12280_), .Y(_12281_));
NAND_g _18793_ (.A(_12270_), .B(_12281_), .Y(_12282_));
NAND_g _18794_ (.A(cpuregs[31][16]), .B(_00007_[2]), .Y(_12283_));
NAND_g _18795_ (.A(cpuregs[27][16]), .B(_09027_), .Y(_12284_));
AND_g _18796_ (.A(_00007_[0]), .B(_12284_), .Y(_12285_));
NAND_g _18797_ (.A(_12283_), .B(_12285_), .Y(_12286_));
NAND_g _18798_ (.A(cpuregs[26][16]), .B(_09027_), .Y(_12287_));
NAND_g _18799_ (.A(cpuregs[30][16]), .B(_00007_[2]), .Y(_12288_));
AND_g _18800_ (.A(_09025_), .B(_12288_), .Y(_12289_));
NAND_g _18801_ (.A(_12287_), .B(_12289_), .Y(_12290_));
AND_g _18802_ (.A(_00007_[3]), .B(_12290_), .Y(_12291_));
NAND_g _18803_ (.A(_12286_), .B(_12291_), .Y(_12292_));
NOR_g _18804_ (.A(cpuregs[18][16]), .B(_00007_[2]), .Y(_12293_));
NOT_g _18805_ (.A(_12293_), .Y(_12294_));
NAND_g _18806_ (.A(_08923_), .B(_00007_[2]), .Y(_12295_));
NAND_g _18807_ (.A(_12294_), .B(_12295_), .Y(_12296_));
NAND_g _18808_ (.A(_09025_), .B(_12296_), .Y(_12297_));
NAND_g _18809_ (.A(_08894_), .B(_00007_[2]), .Y(_12298_));
NOR_g _18810_ (.A(cpuregs[19][16]), .B(_00007_[2]), .Y(_12299_));
NOT_g _18811_ (.A(_12299_), .Y(_12300_));
NAND_g _18812_ (.A(_12298_), .B(_12300_), .Y(_12301_));
NAND_g _18813_ (.A(_00007_[0]), .B(_12301_), .Y(_12302_));
AND_g _18814_ (.A(_09028_), .B(_12302_), .Y(_12303_));
NAND_g _18815_ (.A(_12297_), .B(_12303_), .Y(_12304_));
AND_g _18816_ (.A(_00007_[4]), .B(_12304_), .Y(_12305_));
NAND_g _18817_ (.A(_12292_), .B(_12305_), .Y(_12306_));
NAND_g _18818_ (.A(_12282_), .B(_12306_), .Y(_12307_));
NAND_g _18819_ (.A(_00007_[1]), .B(_12307_), .Y(_12308_));
NAND_g _18820_ (.A(_08912_), .B(_00007_[2]), .Y(_12309_));
NOR_g _18821_ (.A(cpuregs[0][16]), .B(_00007_[2]), .Y(_12310_));
NOR_g _18822_ (.A(_00007_[0]), .B(_12310_), .Y(_12311_));
NAND_g _18823_ (.A(_12309_), .B(_12311_), .Y(_12312_));
NOR_g _18824_ (.A(cpuregs[1][16]), .B(_00007_[2]), .Y(_12313_));
NOT_g _18825_ (.A(_12313_), .Y(_12314_));
NAND_g _18826_ (.A(_08954_), .B(_00007_[2]), .Y(_12315_));
AND_g _18827_ (.A(_00007_[0]), .B(_12315_), .Y(_12316_));
NAND_g _18828_ (.A(_12314_), .B(_12316_), .Y(_12317_));
NAND_g _18829_ (.A(_12312_), .B(_12317_), .Y(_12318_));
NAND_g _18830_ (.A(_09028_), .B(_12318_), .Y(_12319_));
NAND_g _18831_ (.A(cpuregs[9][16]), .B(_09027_), .Y(_12320_));
NAND_g _18832_ (.A(cpuregs[13][16]), .B(_00007_[2]), .Y(_12321_));
NAND_g _18833_ (.A(_12320_), .B(_12321_), .Y(_12322_));
NAND_g _18834_ (.A(_00007_[0]), .B(_12322_), .Y(_12323_));
NAND_g _18835_ (.A(cpuregs[12][16]), .B(_00007_[2]), .Y(_12324_));
NAND_g _18836_ (.A(cpuregs[8][16]), .B(_09027_), .Y(_12325_));
NAND_g _18837_ (.A(_12324_), .B(_12325_), .Y(_12326_));
NAND_g _18838_ (.A(_09025_), .B(_12326_), .Y(_12327_));
NAND_g _18839_ (.A(_12323_), .B(_12327_), .Y(_12328_));
NAND_g _18840_ (.A(_00007_[3]), .B(_12328_), .Y(_12329_));
AND_g _18841_ (.A(_09029_), .B(_12329_), .Y(_12330_));
NAND_g _18842_ (.A(_12319_), .B(_12330_), .Y(_12331_));
NAND_g _18843_ (.A(cpuregs[29][16]), .B(_00007_[2]), .Y(_12332_));
NAND_g _18844_ (.A(cpuregs[25][16]), .B(_09027_), .Y(_12333_));
AND_g _18845_ (.A(_00007_[0]), .B(_12333_), .Y(_12334_));
NAND_g _18846_ (.A(_12332_), .B(_12334_), .Y(_12335_));
NAND_g _18847_ (.A(cpuregs[24][16]), .B(_09027_), .Y(_12336_));
NAND_g _18848_ (.A(cpuregs[28][16]), .B(_00007_[2]), .Y(_12337_));
AND_g _18849_ (.A(_09025_), .B(_12337_), .Y(_12338_));
NAND_g _18850_ (.A(_12336_), .B(_12338_), .Y(_12339_));
AND_g _18851_ (.A(_00007_[3]), .B(_12339_), .Y(_12340_));
NAND_g _18852_ (.A(_12335_), .B(_12340_), .Y(_12341_));
NOR_g _18853_ (.A(cpuregs[16][16]), .B(_00007_[2]), .Y(_12342_));
NOT_g _18854_ (.A(_12342_), .Y(_12343_));
NAND_g _18855_ (.A(_08849_), .B(_00007_[2]), .Y(_12344_));
NAND_g _18856_ (.A(_12343_), .B(_12344_), .Y(_12345_));
NAND_g _18857_ (.A(_09025_), .B(_12345_), .Y(_12346_));
NAND_g _18858_ (.A(_08944_), .B(_09027_), .Y(_12347_));
NAND_g _18859_ (.A(_08993_), .B(_00007_[2]), .Y(_12348_));
NAND_g _18860_ (.A(_12347_), .B(_12348_), .Y(_12349_));
NAND_g _18861_ (.A(_00007_[0]), .B(_12349_), .Y(_12350_));
AND_g _18862_ (.A(_09028_), .B(_12350_), .Y(_12351_));
NAND_g _18863_ (.A(_12346_), .B(_12351_), .Y(_12352_));
AND_g _18864_ (.A(_00007_[4]), .B(_12352_), .Y(_12353_));
NAND_g _18865_ (.A(_12341_), .B(_12353_), .Y(_12354_));
NAND_g _18866_ (.A(_12331_), .B(_12354_), .Y(_12355_));
NAND_g _18867_ (.A(_09026_), .B(_12355_), .Y(_12356_));
AND_g _18868_ (.A(_12308_), .B(_12356_), .Y(_12357_));
NAND_g _18869_ (.A(_11170_), .B(_12357_), .Y(_12358_));
NAND_g _18870_ (.A(decoded_imm[16]), .B(_10606_), .Y(_12359_));
AND_g _18871_ (.A(_10603_), .B(_12359_), .Y(_12360_));
NAND_g _18872_ (.A(_12358_), .B(_12360_), .Y(_12361_));
AND_g _18873_ (.A(_12260_), .B(_12361_), .Y(_00291_));
NAND_g _18874_ (.A(_08827_), .B(_10604_), .Y(_12362_));
NAND_g _18875_ (.A(cpuregs[22][17]), .B(_00007_[1]), .Y(_12363_));
NAND_g _18876_ (.A(cpuregs[20][17]), .B(_09026_), .Y(_12364_));
NAND_g _18877_ (.A(_12363_), .B(_12364_), .Y(_12365_));
NAND_g _18878_ (.A(_00007_[2]), .B(_12365_), .Y(_12366_));
NAND_g _18879_ (.A(cpuregs[18][17]), .B(_00007_[1]), .Y(_12367_));
NAND_g _18880_ (.A(cpuregs[16][17]), .B(_09026_), .Y(_12368_));
NAND_g _18881_ (.A(_12367_), .B(_12368_), .Y(_12369_));
NAND_g _18882_ (.A(_09027_), .B(_12369_), .Y(_12370_));
NAND_g _18883_ (.A(_12366_), .B(_12370_), .Y(_12371_));
AND_g _18884_ (.A(_09025_), .B(_12371_), .Y(_12372_));
NOT_g _18885_ (.A(_12372_), .Y(_12373_));
NAND_g _18886_ (.A(cpuregs[23][17]), .B(_00007_[1]), .Y(_12374_));
NAND_g _18887_ (.A(cpuregs[21][17]), .B(_09026_), .Y(_12375_));
NAND_g _18888_ (.A(_12374_), .B(_12375_), .Y(_12376_));
NAND_g _18889_ (.A(_00007_[2]), .B(_12376_), .Y(_12377_));
NAND_g _18890_ (.A(cpuregs[19][17]), .B(_00007_[1]), .Y(_12378_));
NAND_g _18891_ (.A(cpuregs[17][17]), .B(_09026_), .Y(_12379_));
NAND_g _18892_ (.A(_12378_), .B(_12379_), .Y(_12380_));
NAND_g _18893_ (.A(_09027_), .B(_12380_), .Y(_12381_));
NAND_g _18894_ (.A(_12377_), .B(_12381_), .Y(_12382_));
NAND_g _18895_ (.A(_00007_[0]), .B(_12382_), .Y(_12383_));
AND_g _18896_ (.A(_09028_), .B(_12383_), .Y(_12384_));
NAND_g _18897_ (.A(_12373_), .B(_12384_), .Y(_12385_));
NAND_g _18898_ (.A(cpuregs[31][17]), .B(_00007_[2]), .Y(_12386_));
NAND_g _18899_ (.A(cpuregs[27][17]), .B(_09027_), .Y(_12387_));
AND_g _18900_ (.A(_00007_[0]), .B(_12387_), .Y(_12388_));
NAND_g _18901_ (.A(_12386_), .B(_12388_), .Y(_12389_));
NAND_g _18902_ (.A(cpuregs[26][17]), .B(_09027_), .Y(_12390_));
NAND_g _18903_ (.A(cpuregs[30][17]), .B(_00007_[2]), .Y(_12391_));
AND_g _18904_ (.A(_09025_), .B(_12391_), .Y(_12392_));
NAND_g _18905_ (.A(_12390_), .B(_12392_), .Y(_12393_));
AND_g _18906_ (.A(_00007_[1]), .B(_12393_), .Y(_12394_));
NAND_g _18907_ (.A(_12389_), .B(_12394_), .Y(_12395_));
NAND_g _18908_ (.A(cpuregs[25][17]), .B(_09027_), .Y(_12396_));
NAND_g _18909_ (.A(cpuregs[29][17]), .B(_00007_[2]), .Y(_12397_));
AND_g _18910_ (.A(_00007_[0]), .B(_12397_), .Y(_12398_));
NAND_g _18911_ (.A(_12396_), .B(_12398_), .Y(_12399_));
NAND_g _18912_ (.A(cpuregs[24][17]), .B(_09027_), .Y(_12400_));
NAND_g _18913_ (.A(cpuregs[28][17]), .B(_00007_[2]), .Y(_12401_));
AND_g _18914_ (.A(_09025_), .B(_12401_), .Y(_12402_));
NAND_g _18915_ (.A(_12400_), .B(_12402_), .Y(_12403_));
AND_g _18916_ (.A(_09026_), .B(_12403_), .Y(_12404_));
NAND_g _18917_ (.A(_12399_), .B(_12404_), .Y(_12405_));
AND_g _18918_ (.A(_00007_[3]), .B(_12405_), .Y(_12406_));
NAND_g _18919_ (.A(_12395_), .B(_12406_), .Y(_12407_));
NAND_g _18920_ (.A(_12385_), .B(_12407_), .Y(_12408_));
NAND_g _18921_ (.A(_00007_[4]), .B(_12408_), .Y(_12409_));
NAND_g _18922_ (.A(cpuregs[3][17]), .B(_09027_), .Y(_12410_));
NAND_g _18923_ (.A(cpuregs[7][17]), .B(_00007_[2]), .Y(_12411_));
AND_g _18924_ (.A(_00007_[0]), .B(_12411_), .Y(_12412_));
NAND_g _18925_ (.A(_12410_), .B(_12412_), .Y(_12413_));
NAND_g _18926_ (.A(cpuregs[2][17]), .B(_09027_), .Y(_12414_));
NAND_g _18927_ (.A(cpuregs[6][17]), .B(_00007_[2]), .Y(_12415_));
AND_g _18928_ (.A(_09025_), .B(_12415_), .Y(_12416_));
NAND_g _18929_ (.A(_12414_), .B(_12416_), .Y(_12417_));
AND_g _18930_ (.A(_00007_[1]), .B(_12417_), .Y(_12418_));
NAND_g _18931_ (.A(_12413_), .B(_12418_), .Y(_12419_));
NAND_g _18932_ (.A(cpuregs[1][17]), .B(_09027_), .Y(_12420_));
NAND_g _18933_ (.A(cpuregs[5][17]), .B(_00007_[2]), .Y(_12421_));
AND_g _18934_ (.A(_00007_[0]), .B(_12421_), .Y(_12422_));
NAND_g _18935_ (.A(_12420_), .B(_12422_), .Y(_12423_));
NAND_g _18936_ (.A(cpuregs[0][17]), .B(_09027_), .Y(_12424_));
NAND_g _18937_ (.A(cpuregs[4][17]), .B(_00007_[2]), .Y(_12425_));
AND_g _18938_ (.A(_09025_), .B(_12425_), .Y(_12426_));
NAND_g _18939_ (.A(_12424_), .B(_12426_), .Y(_12427_));
AND_g _18940_ (.A(_09026_), .B(_12427_), .Y(_12428_));
NAND_g _18941_ (.A(_12423_), .B(_12428_), .Y(_12429_));
AND_g _18942_ (.A(_09028_), .B(_12429_), .Y(_12430_));
NAND_g _18943_ (.A(_12419_), .B(_12430_), .Y(_12431_));
NAND_g _18944_ (.A(cpuregs[12][17]), .B(_09025_), .Y(_12432_));
NAND_g _18945_ (.A(cpuregs[13][17]), .B(_00007_[0]), .Y(_12433_));
NAND_g _18946_ (.A(_12432_), .B(_12433_), .Y(_12434_));
NAND_g _18947_ (.A(_00007_[2]), .B(_12434_), .Y(_12435_));
NAND_g _18948_ (.A(cpuregs[8][17]), .B(_09025_), .Y(_12436_));
NAND_g _18949_ (.A(cpuregs[9][17]), .B(_00007_[0]), .Y(_12437_));
NAND_g _18950_ (.A(_12436_), .B(_12437_), .Y(_12438_));
NAND_g _18951_ (.A(_09027_), .B(_12438_), .Y(_12439_));
NAND_g _18952_ (.A(_12435_), .B(_12439_), .Y(_12440_));
NAND_g _18953_ (.A(_09026_), .B(_12440_), .Y(_12441_));
NAND_g _18954_ (.A(cpuregs[14][17]), .B(_09025_), .Y(_12442_));
NAND_g _18955_ (.A(cpuregs[15][17]), .B(_00007_[0]), .Y(_12443_));
NAND_g _18956_ (.A(_12442_), .B(_12443_), .Y(_12444_));
NAND_g _18957_ (.A(_00007_[2]), .B(_12444_), .Y(_12445_));
NAND_g _18958_ (.A(cpuregs[10][17]), .B(_09025_), .Y(_12446_));
NAND_g _18959_ (.A(cpuregs[11][17]), .B(_00007_[0]), .Y(_12447_));
NAND_g _18960_ (.A(_12446_), .B(_12447_), .Y(_12448_));
NAND_g _18961_ (.A(_09027_), .B(_12448_), .Y(_12449_));
NAND_g _18962_ (.A(_12445_), .B(_12449_), .Y(_12450_));
NAND_g _18963_ (.A(_00007_[1]), .B(_12450_), .Y(_12451_));
AND_g _18964_ (.A(_00007_[3]), .B(_12451_), .Y(_12452_));
NAND_g _18965_ (.A(_12441_), .B(_12452_), .Y(_12453_));
NAND_g _18966_ (.A(_12431_), .B(_12453_), .Y(_12454_));
NAND_g _18967_ (.A(_09029_), .B(_12454_), .Y(_12455_));
AND_g _18968_ (.A(_12409_), .B(_12455_), .Y(_12456_));
NAND_g _18969_ (.A(_11170_), .B(_12456_), .Y(_12457_));
NAND_g _18970_ (.A(decoded_imm[17]), .B(_10606_), .Y(_12458_));
AND_g _18971_ (.A(_10603_), .B(_12458_), .Y(_12459_));
NAND_g _18972_ (.A(_12457_), .B(_12459_), .Y(_12460_));
AND_g _18973_ (.A(_12362_), .B(_12460_), .Y(_00292_));
NAND_g _18974_ (.A(_08828_), .B(_10604_), .Y(_12461_));
NAND_g _18975_ (.A(cpuregs[22][18]), .B(_00007_[1]), .Y(_12462_));
NAND_g _18976_ (.A(cpuregs[20][18]), .B(_09026_), .Y(_12463_));
NAND_g _18977_ (.A(_12462_), .B(_12463_), .Y(_12464_));
NAND_g _18978_ (.A(_00007_[2]), .B(_12464_), .Y(_12465_));
NAND_g _18979_ (.A(cpuregs[18][18]), .B(_00007_[1]), .Y(_12466_));
NAND_g _18980_ (.A(cpuregs[16][18]), .B(_09026_), .Y(_12467_));
NAND_g _18981_ (.A(_12466_), .B(_12467_), .Y(_12468_));
NAND_g _18982_ (.A(_09027_), .B(_12468_), .Y(_12469_));
NAND_g _18983_ (.A(_12465_), .B(_12469_), .Y(_12470_));
AND_g _18984_ (.A(_09025_), .B(_12470_), .Y(_12471_));
NOT_g _18985_ (.A(_12471_), .Y(_12472_));
NAND_g _18986_ (.A(cpuregs[23][18]), .B(_00007_[1]), .Y(_12473_));
NAND_g _18987_ (.A(cpuregs[21][18]), .B(_09026_), .Y(_12474_));
NAND_g _18988_ (.A(_12473_), .B(_12474_), .Y(_12475_));
NAND_g _18989_ (.A(_00007_[2]), .B(_12475_), .Y(_12476_));
NAND_g _18990_ (.A(cpuregs[19][18]), .B(_00007_[1]), .Y(_12477_));
NAND_g _18991_ (.A(cpuregs[17][18]), .B(_09026_), .Y(_12478_));
NAND_g _18992_ (.A(_12477_), .B(_12478_), .Y(_12479_));
NAND_g _18993_ (.A(_09027_), .B(_12479_), .Y(_12480_));
NAND_g _18994_ (.A(_12476_), .B(_12480_), .Y(_12481_));
NAND_g _18995_ (.A(_00007_[0]), .B(_12481_), .Y(_12482_));
AND_g _18996_ (.A(_09028_), .B(_12482_), .Y(_12483_));
NAND_g _18997_ (.A(_12472_), .B(_12483_), .Y(_12484_));
NAND_g _18998_ (.A(cpuregs[31][18]), .B(_00007_[2]), .Y(_12485_));
NAND_g _18999_ (.A(cpuregs[27][18]), .B(_09027_), .Y(_12486_));
AND_g _19000_ (.A(_00007_[0]), .B(_12486_), .Y(_12487_));
NAND_g _19001_ (.A(_12485_), .B(_12487_), .Y(_12488_));
NAND_g _19002_ (.A(cpuregs[26][18]), .B(_09027_), .Y(_12489_));
NAND_g _19003_ (.A(cpuregs[30][18]), .B(_00007_[2]), .Y(_12490_));
AND_g _19004_ (.A(_09025_), .B(_12490_), .Y(_12491_));
NAND_g _19005_ (.A(_12489_), .B(_12491_), .Y(_12492_));
AND_g _19006_ (.A(_00007_[1]), .B(_12492_), .Y(_12493_));
NAND_g _19007_ (.A(_12488_), .B(_12493_), .Y(_12494_));
NAND_g _19008_ (.A(cpuregs[25][18]), .B(_09027_), .Y(_12495_));
NAND_g _19009_ (.A(cpuregs[29][18]), .B(_00007_[2]), .Y(_12496_));
AND_g _19010_ (.A(_00007_[0]), .B(_12496_), .Y(_12497_));
NAND_g _19011_ (.A(_12495_), .B(_12497_), .Y(_12498_));
NAND_g _19012_ (.A(cpuregs[24][18]), .B(_09027_), .Y(_12499_));
NAND_g _19013_ (.A(cpuregs[28][18]), .B(_00007_[2]), .Y(_12500_));
AND_g _19014_ (.A(_09025_), .B(_12500_), .Y(_12501_));
NAND_g _19015_ (.A(_12499_), .B(_12501_), .Y(_12502_));
AND_g _19016_ (.A(_09026_), .B(_12502_), .Y(_12503_));
NAND_g _19017_ (.A(_12498_), .B(_12503_), .Y(_12504_));
AND_g _19018_ (.A(_00007_[3]), .B(_12504_), .Y(_12505_));
NAND_g _19019_ (.A(_12494_), .B(_12505_), .Y(_12506_));
NAND_g _19020_ (.A(_12484_), .B(_12506_), .Y(_12507_));
AND_g _19021_ (.A(_00007_[4]), .B(_12507_), .Y(_12508_));
NAND_g _19022_ (.A(cpuregs[3][18]), .B(_09027_), .Y(_12509_));
NAND_g _19023_ (.A(cpuregs[7][18]), .B(_00007_[2]), .Y(_12510_));
AND_g _19024_ (.A(_00007_[0]), .B(_12510_), .Y(_12511_));
NAND_g _19025_ (.A(_12509_), .B(_12511_), .Y(_12512_));
NAND_g _19026_ (.A(cpuregs[2][18]), .B(_09027_), .Y(_12513_));
NAND_g _19027_ (.A(cpuregs[6][18]), .B(_00007_[2]), .Y(_12514_));
AND_g _19028_ (.A(_09025_), .B(_12514_), .Y(_12515_));
NAND_g _19029_ (.A(_12513_), .B(_12515_), .Y(_12516_));
AND_g _19030_ (.A(_00007_[1]), .B(_12516_), .Y(_12517_));
NAND_g _19031_ (.A(_12512_), .B(_12517_), .Y(_12518_));
NAND_g _19032_ (.A(cpuregs[1][18]), .B(_09027_), .Y(_12519_));
NAND_g _19033_ (.A(cpuregs[5][18]), .B(_00007_[2]), .Y(_12520_));
AND_g _19034_ (.A(_00007_[0]), .B(_12520_), .Y(_12521_));
NAND_g _19035_ (.A(_12519_), .B(_12521_), .Y(_12522_));
NAND_g _19036_ (.A(cpuregs[0][18]), .B(_09027_), .Y(_12523_));
NAND_g _19037_ (.A(cpuregs[4][18]), .B(_00007_[2]), .Y(_12524_));
AND_g _19038_ (.A(_09025_), .B(_12524_), .Y(_12525_));
NAND_g _19039_ (.A(_12523_), .B(_12525_), .Y(_12526_));
AND_g _19040_ (.A(_09026_), .B(_12526_), .Y(_12527_));
NAND_g _19041_ (.A(_12522_), .B(_12527_), .Y(_12528_));
AND_g _19042_ (.A(_09028_), .B(_12528_), .Y(_12529_));
NAND_g _19043_ (.A(_12518_), .B(_12529_), .Y(_12530_));
NAND_g _19044_ (.A(cpuregs[12][18]), .B(_09025_), .Y(_12531_));
NAND_g _19045_ (.A(cpuregs[13][18]), .B(_00007_[0]), .Y(_12532_));
NAND_g _19046_ (.A(_12531_), .B(_12532_), .Y(_12533_));
NAND_g _19047_ (.A(_00007_[2]), .B(_12533_), .Y(_12534_));
NAND_g _19048_ (.A(cpuregs[8][18]), .B(_09025_), .Y(_12535_));
NAND_g _19049_ (.A(cpuregs[9][18]), .B(_00007_[0]), .Y(_12536_));
NAND_g _19050_ (.A(_12535_), .B(_12536_), .Y(_12537_));
NAND_g _19051_ (.A(_09027_), .B(_12537_), .Y(_12538_));
NAND_g _19052_ (.A(_12534_), .B(_12538_), .Y(_12539_));
NAND_g _19053_ (.A(_09026_), .B(_12539_), .Y(_12540_));
NAND_g _19054_ (.A(cpuregs[14][18]), .B(_09025_), .Y(_12541_));
NAND_g _19055_ (.A(cpuregs[15][18]), .B(_00007_[0]), .Y(_12542_));
NAND_g _19056_ (.A(_12541_), .B(_12542_), .Y(_12543_));
NAND_g _19057_ (.A(_00007_[2]), .B(_12543_), .Y(_12544_));
NAND_g _19058_ (.A(cpuregs[10][18]), .B(_09025_), .Y(_12545_));
NAND_g _19059_ (.A(cpuregs[11][18]), .B(_00007_[0]), .Y(_12546_));
NAND_g _19060_ (.A(_12545_), .B(_12546_), .Y(_12547_));
NAND_g _19061_ (.A(_09027_), .B(_12547_), .Y(_12548_));
NAND_g _19062_ (.A(_12544_), .B(_12548_), .Y(_12549_));
NAND_g _19063_ (.A(_00007_[1]), .B(_12549_), .Y(_12550_));
AND_g _19064_ (.A(_00007_[3]), .B(_12550_), .Y(_12551_));
NAND_g _19065_ (.A(_12540_), .B(_12551_), .Y(_12552_));
NAND_g _19066_ (.A(_12530_), .B(_12552_), .Y(_12553_));
AND_g _19067_ (.A(_09029_), .B(_12553_), .Y(_12554_));
NOR_g _19068_ (.A(_12508_), .B(_12554_), .Y(_12555_));
NAND_g _19069_ (.A(_11170_), .B(_12555_), .Y(_12556_));
NAND_g _19070_ (.A(decoded_imm[18]), .B(_10606_), .Y(_12557_));
AND_g _19071_ (.A(_10603_), .B(_12557_), .Y(_12558_));
NAND_g _19072_ (.A(_12556_), .B(_12558_), .Y(_12559_));
AND_g _19073_ (.A(_12461_), .B(_12559_), .Y(_00293_));
NAND_g _19074_ (.A(_08829_), .B(_10604_), .Y(_12560_));
NAND_g _19075_ (.A(cpuregs[17][19]), .B(_09027_), .Y(_12561_));
NAND_g _19076_ (.A(cpuregs[21][19]), .B(_00007_[2]), .Y(_12562_));
NAND_g _19077_ (.A(_12561_), .B(_12562_), .Y(_12563_));
NAND_g _19078_ (.A(_00007_[0]), .B(_12563_), .Y(_12564_));
NAND_g _19079_ (.A(cpuregs[20][19]), .B(_00007_[2]), .Y(_12565_));
NAND_g _19080_ (.A(cpuregs[16][19]), .B(_09027_), .Y(_12566_));
NAND_g _19081_ (.A(_12565_), .B(_12566_), .Y(_12567_));
NAND_g _19082_ (.A(_09025_), .B(_12567_), .Y(_12568_));
NAND_g _19083_ (.A(_12564_), .B(_12568_), .Y(_12569_));
NAND_g _19084_ (.A(_09028_), .B(_12569_), .Y(_12570_));
NAND_g _19085_ (.A(cpuregs[25][19]), .B(_09027_), .Y(_12571_));
NAND_g _19086_ (.A(cpuregs[29][19]), .B(_00007_[2]), .Y(_12572_));
NAND_g _19087_ (.A(_12571_), .B(_12572_), .Y(_12573_));
NAND_g _19088_ (.A(_00007_[0]), .B(_12573_), .Y(_12574_));
NAND_g _19089_ (.A(cpuregs[28][19]), .B(_00007_[2]), .Y(_12575_));
NAND_g _19090_ (.A(cpuregs[24][19]), .B(_09027_), .Y(_12576_));
NAND_g _19091_ (.A(_12575_), .B(_12576_), .Y(_12577_));
NAND_g _19092_ (.A(_09025_), .B(_12577_), .Y(_12578_));
NAND_g _19093_ (.A(_12574_), .B(_12578_), .Y(_12579_));
NAND_g _19094_ (.A(_00007_[3]), .B(_12579_), .Y(_12580_));
NAND_g _19095_ (.A(cpuregs[31][19]), .B(_00007_[0]), .Y(_12581_));
NAND_g _19096_ (.A(cpuregs[30][19]), .B(_09025_), .Y(_12582_));
AND_g _19097_ (.A(_00007_[2]), .B(_12582_), .Y(_12583_));
NAND_g _19098_ (.A(_12581_), .B(_12583_), .Y(_12584_));
NAND_g _19099_ (.A(cpuregs[27][19]), .B(_00007_[0]), .Y(_12585_));
NAND_g _19100_ (.A(cpuregs[26][19]), .B(_09025_), .Y(_12586_));
AND_g _19101_ (.A(_09027_), .B(_12586_), .Y(_12587_));
NAND_g _19102_ (.A(_12585_), .B(_12587_), .Y(_12588_));
AND_g _19103_ (.A(_00007_[3]), .B(_12588_), .Y(_12589_));
NAND_g _19104_ (.A(_12584_), .B(_12589_), .Y(_12590_));
NAND_g _19105_ (.A(cpuregs[23][19]), .B(_00007_[0]), .Y(_12591_));
NAND_g _19106_ (.A(cpuregs[22][19]), .B(_09025_), .Y(_12592_));
AND_g _19107_ (.A(_00007_[2]), .B(_12592_), .Y(_12593_));
NAND_g _19108_ (.A(_12591_), .B(_12593_), .Y(_12594_));
NAND_g _19109_ (.A(cpuregs[19][19]), .B(_00007_[0]), .Y(_12595_));
NAND_g _19110_ (.A(cpuregs[18][19]), .B(_09025_), .Y(_12596_));
AND_g _19111_ (.A(_09027_), .B(_12596_), .Y(_12597_));
NAND_g _19112_ (.A(_12595_), .B(_12597_), .Y(_12598_));
AND_g _19113_ (.A(_09028_), .B(_12598_), .Y(_12599_));
NAND_g _19114_ (.A(_12594_), .B(_12599_), .Y(_12600_));
NAND_g _19115_ (.A(_12590_), .B(_12600_), .Y(_12601_));
NAND_g _19116_ (.A(_00007_[1]), .B(_12601_), .Y(_12602_));
NAND_g _19117_ (.A(_12570_), .B(_12580_), .Y(_12603_));
NAND_g _19118_ (.A(_09026_), .B(_12603_), .Y(_12604_));
AND_g _19119_ (.A(_00007_[4]), .B(_12602_), .Y(_12605_));
AND_g _19120_ (.A(_12604_), .B(_12605_), .Y(_12606_));
NOR_g _19121_ (.A(cpuregs[9][19]), .B(_00007_[2]), .Y(_12607_));
NAND_g _19122_ (.A(_08930_), .B(_00007_[2]), .Y(_12608_));
NOR_g _19123_ (.A(cpuregs[8][19]), .B(_00007_[2]), .Y(_12609_));
NOR_g _19124_ (.A(cpuregs[12][19]), .B(_09027_), .Y(_12610_));
NOR_g _19125_ (.A(_12609_), .B(_12610_), .Y(_12611_));
NAND_g _19126_ (.A(_00007_[0]), .B(_12608_), .Y(_12612_));
NOR_g _19127_ (.A(_12607_), .B(_12612_), .Y(_12613_));
AND_g _19128_ (.A(_09025_), .B(_12611_), .Y(_12614_));
NOR_g _19129_ (.A(_12613_), .B(_12614_), .Y(_12615_));
NOR_g _19130_ (.A(_09028_), .B(_12615_), .Y(_12616_));
NAND_g _19131_ (.A(cpuregs[4][19]), .B(_00007_[2]), .Y(_12617_));
NAND_g _19132_ (.A(cpuregs[0][19]), .B(_09027_), .Y(_12618_));
AND_g _19133_ (.A(_12617_), .B(_12618_), .Y(_12619_));
NAND_g _19134_ (.A(_09025_), .B(_12619_), .Y(_12620_));
NAND_g _19135_ (.A(cpuregs[5][19]), .B(_00007_[2]), .Y(_12621_));
NAND_g _19136_ (.A(cpuregs[1][19]), .B(_09027_), .Y(_12622_));
AND_g _19137_ (.A(_00007_[0]), .B(_12622_), .Y(_12623_));
NAND_g _19138_ (.A(_12621_), .B(_12623_), .Y(_12624_));
AND_g _19139_ (.A(_12620_), .B(_12624_), .Y(_12625_));
NAND_g _19140_ (.A(_09028_), .B(_12625_), .Y(_12626_));
NAND_g _19141_ (.A(_09026_), .B(_12626_), .Y(_12627_));
NOR_g _19142_ (.A(_12616_), .B(_12627_), .Y(_12628_));
NAND_g _19143_ (.A(cpuregs[6][19]), .B(_00007_[2]), .Y(_12629_));
NAND_g _19144_ (.A(cpuregs[2][19]), .B(_09027_), .Y(_12630_));
AND_g _19145_ (.A(_12629_), .B(_12630_), .Y(_12631_));
NAND_g _19146_ (.A(_09025_), .B(_12631_), .Y(_12632_));
NAND_g _19147_ (.A(cpuregs[7][19]), .B(_00007_[2]), .Y(_12633_));
NAND_g _19148_ (.A(cpuregs[3][19]), .B(_09027_), .Y(_12634_));
AND_g _19149_ (.A(_00007_[0]), .B(_12634_), .Y(_12635_));
NAND_g _19150_ (.A(_12633_), .B(_12635_), .Y(_12636_));
AND_g _19151_ (.A(_12632_), .B(_12636_), .Y(_12637_));
NAND_g _19152_ (.A(_09028_), .B(_12637_), .Y(_12638_));
NOR_g _19153_ (.A(cpuregs[10][19]), .B(_00007_[2]), .Y(_12639_));
AND_g _19154_ (.A(_08939_), .B(_00007_[2]), .Y(_12640_));
NOR_g _19155_ (.A(_12639_), .B(_12640_), .Y(_12641_));
NOR_g _19156_ (.A(cpuregs[11][19]), .B(_00007_[2]), .Y(_12642_));
NOT_g _19157_ (.A(_12642_), .Y(_12643_));
NAND_g _19158_ (.A(_08809_), .B(_00007_[2]), .Y(_12644_));
AND_g _19159_ (.A(_00007_[0]), .B(_12644_), .Y(_12645_));
NAND_g _19160_ (.A(_12643_), .B(_12645_), .Y(_12646_));
NAND_g _19161_ (.A(_09025_), .B(_12641_), .Y(_12647_));
NAND_g _19162_ (.A(_12646_), .B(_12647_), .Y(_12648_));
NAND_g _19163_ (.A(_00007_[3]), .B(_12648_), .Y(_12649_));
AND_g _19164_ (.A(_00007_[1]), .B(_12649_), .Y(_12650_));
AND_g _19165_ (.A(_12638_), .B(_12650_), .Y(_12651_));
NOR_g _19166_ (.A(_12628_), .B(_12651_), .Y(_12652_));
NOR_g _19167_ (.A(_00007_[4]), .B(_12652_), .Y(_12653_));
NOR_g _19168_ (.A(_12606_), .B(_12653_), .Y(_12654_));
NAND_g _19169_ (.A(_11170_), .B(_12654_), .Y(_12655_));
NAND_g _19170_ (.A(decoded_imm[19]), .B(_10606_), .Y(_12656_));
AND_g _19171_ (.A(_10603_), .B(_12656_), .Y(_12657_));
NAND_g _19172_ (.A(_12655_), .B(_12657_), .Y(_12658_));
AND_g _19173_ (.A(_12560_), .B(_12658_), .Y(_00294_));
NAND_g _19174_ (.A(_08830_), .B(_10604_), .Y(_12659_));
NAND_g _19175_ (.A(cpuregs[20][20]), .B(_00007_[2]), .Y(_12660_));
NAND_g _19176_ (.A(cpuregs[16][20]), .B(_09027_), .Y(_12661_));
NAND_g _19177_ (.A(_12660_), .B(_12661_), .Y(_12662_));
NAND_g _19178_ (.A(_09025_), .B(_12662_), .Y(_12663_));
NAND_g _19179_ (.A(cpuregs[17][20]), .B(_09027_), .Y(_12664_));
NAND_g _19180_ (.A(cpuregs[21][20]), .B(_00007_[2]), .Y(_12665_));
NAND_g _19181_ (.A(_12664_), .B(_12665_), .Y(_12666_));
NAND_g _19182_ (.A(_00007_[0]), .B(_12666_), .Y(_12667_));
AND_g _19183_ (.A(_12663_), .B(_12667_), .Y(_12668_));
NAND_g _19184_ (.A(_09028_), .B(_12668_), .Y(_12669_));
NAND_g _19185_ (.A(cpuregs[28][20]), .B(_00007_[2]), .Y(_12670_));
NAND_g _19186_ (.A(cpuregs[24][20]), .B(_09027_), .Y(_12671_));
NAND_g _19187_ (.A(_12670_), .B(_12671_), .Y(_12672_));
NAND_g _19188_ (.A(_09025_), .B(_12672_), .Y(_12673_));
NAND_g _19189_ (.A(cpuregs[25][20]), .B(_09027_), .Y(_12674_));
NAND_g _19190_ (.A(cpuregs[29][20]), .B(_00007_[2]), .Y(_12675_));
NAND_g _19191_ (.A(_12674_), .B(_12675_), .Y(_12676_));
NAND_g _19192_ (.A(_00007_[0]), .B(_12676_), .Y(_12677_));
AND_g _19193_ (.A(_12673_), .B(_12677_), .Y(_12678_));
NAND_g _19194_ (.A(_00007_[3]), .B(_12678_), .Y(_12679_));
AND_g _19195_ (.A(_12669_), .B(_12679_), .Y(_12680_));
NAND_g _19196_ (.A(cpuregs[27][20]), .B(_00007_[0]), .Y(_12681_));
NAND_g _19197_ (.A(cpuregs[26][20]), .B(_09025_), .Y(_12682_));
AND_g _19198_ (.A(_09027_), .B(_12682_), .Y(_12683_));
NAND_g _19199_ (.A(_12681_), .B(_12683_), .Y(_12684_));
NAND_g _19200_ (.A(cpuregs[31][20]), .B(_00007_[0]), .Y(_12685_));
NAND_g _19201_ (.A(cpuregs[30][20]), .B(_09025_), .Y(_12686_));
AND_g _19202_ (.A(_00007_[2]), .B(_12686_), .Y(_12687_));
NAND_g _19203_ (.A(_12685_), .B(_12687_), .Y(_12688_));
NAND_g _19204_ (.A(_12684_), .B(_12688_), .Y(_12689_));
NAND_g _19205_ (.A(_00007_[3]), .B(_12689_), .Y(_12690_));
NAND_g _19206_ (.A(cpuregs[19][20]), .B(_00007_[0]), .Y(_12691_));
NAND_g _19207_ (.A(cpuregs[18][20]), .B(_09025_), .Y(_12692_));
AND_g _19208_ (.A(_09027_), .B(_12692_), .Y(_12693_));
NAND_g _19209_ (.A(_12691_), .B(_12693_), .Y(_12694_));
NAND_g _19210_ (.A(cpuregs[23][20]), .B(_00007_[0]), .Y(_12695_));
NAND_g _19211_ (.A(cpuregs[22][20]), .B(_09025_), .Y(_12696_));
AND_g _19212_ (.A(_00007_[2]), .B(_12696_), .Y(_12697_));
NAND_g _19213_ (.A(_12695_), .B(_12697_), .Y(_12698_));
NAND_g _19214_ (.A(_12694_), .B(_12698_), .Y(_12699_));
NAND_g _19215_ (.A(_09028_), .B(_12699_), .Y(_12700_));
AND_g _19216_ (.A(_12690_), .B(_12700_), .Y(_12701_));
NAND_g _19217_ (.A(_00007_[1]), .B(_12701_), .Y(_12702_));
NAND_g _19218_ (.A(_09026_), .B(_12680_), .Y(_12703_));
AND_g _19219_ (.A(_00007_[4]), .B(_12703_), .Y(_12704_));
AND_g _19220_ (.A(_12702_), .B(_12704_), .Y(_12705_));
NOR_g _19221_ (.A(cpuregs[11][20]), .B(_00007_[2]), .Y(_12706_));
AND_g _19222_ (.A(_08810_), .B(_00007_[2]), .Y(_12707_));
NOR_g _19223_ (.A(_12706_), .B(_12707_), .Y(_12708_));
NOR_g _19224_ (.A(_09025_), .B(_12708_), .Y(_12709_));
NOR_g _19225_ (.A(cpuregs[10][20]), .B(_00007_[2]), .Y(_12710_));
AND_g _19226_ (.A(_08940_), .B(_00007_[2]), .Y(_12711_));
NOR_g _19227_ (.A(_12710_), .B(_12711_), .Y(_12712_));
NOR_g _19228_ (.A(_00007_[0]), .B(_12712_), .Y(_12713_));
NOR_g _19229_ (.A(_12709_), .B(_12713_), .Y(_12714_));
NAND_g _19230_ (.A(cpuregs[7][20]), .B(_00007_[2]), .Y(_12715_));
NAND_g _19231_ (.A(cpuregs[3][20]), .B(_09027_), .Y(_12716_));
AND_g _19232_ (.A(_00007_[0]), .B(_12716_), .Y(_12717_));
NAND_g _19233_ (.A(_12715_), .B(_12717_), .Y(_12718_));
NAND_g _19234_ (.A(cpuregs[6][20]), .B(_00007_[2]), .Y(_12719_));
NAND_g _19235_ (.A(cpuregs[2][20]), .B(_09027_), .Y(_12720_));
AND_g _19236_ (.A(_12719_), .B(_12720_), .Y(_12721_));
NAND_g _19237_ (.A(_09025_), .B(_12721_), .Y(_12722_));
AND_g _19238_ (.A(_12718_), .B(_12722_), .Y(_12723_));
NAND_g _19239_ (.A(_00007_[3]), .B(_12714_), .Y(_12724_));
NAND_g _19240_ (.A(_09028_), .B(_12723_), .Y(_12725_));
AND_g _19241_ (.A(_00007_[1]), .B(_12725_), .Y(_12726_));
AND_g _19242_ (.A(_12724_), .B(_12726_), .Y(_12727_));
NOR_g _19243_ (.A(cpuregs[8][20]), .B(_00007_[2]), .Y(_12728_));
NOR_g _19244_ (.A(cpuregs[12][20]), .B(_09027_), .Y(_12729_));
NOR_g _19245_ (.A(_12728_), .B(_12729_), .Y(_12730_));
NOR_g _19246_ (.A(cpuregs[9][20]), .B(_00007_[2]), .Y(_12731_));
NAND_g _19247_ (.A(_08931_), .B(_00007_[2]), .Y(_12732_));
NAND_g _19248_ (.A(_00007_[0]), .B(_12732_), .Y(_12733_));
NOR_g _19249_ (.A(_12731_), .B(_12733_), .Y(_12734_));
AND_g _19250_ (.A(_09025_), .B(_12730_), .Y(_12735_));
NOR_g _19251_ (.A(_12734_), .B(_12735_), .Y(_12736_));
NAND_g _19252_ (.A(_00007_[3]), .B(_12736_), .Y(_12737_));
NAND_g _19253_ (.A(cpuregs[5][20]), .B(_00007_[2]), .Y(_12738_));
NAND_g _19254_ (.A(cpuregs[1][20]), .B(_09027_), .Y(_12739_));
AND_g _19255_ (.A(_00007_[0]), .B(_12739_), .Y(_12740_));
NAND_g _19256_ (.A(_12738_), .B(_12740_), .Y(_12741_));
NAND_g _19257_ (.A(cpuregs[4][20]), .B(_00007_[2]), .Y(_12742_));
NAND_g _19258_ (.A(cpuregs[0][20]), .B(_09027_), .Y(_12743_));
AND_g _19259_ (.A(_12742_), .B(_12743_), .Y(_12744_));
NAND_g _19260_ (.A(_09025_), .B(_12744_), .Y(_12745_));
NAND_g _19261_ (.A(_12741_), .B(_12745_), .Y(_12746_));
NAND_g _19262_ (.A(_09028_), .B(_12746_), .Y(_12747_));
NAND_g _19263_ (.A(_12737_), .B(_12747_), .Y(_12748_));
AND_g _19264_ (.A(_09026_), .B(_12748_), .Y(_12749_));
NOR_g _19265_ (.A(_12727_), .B(_12749_), .Y(_12750_));
NOR_g _19266_ (.A(_00007_[4]), .B(_12750_), .Y(_12751_));
NOR_g _19267_ (.A(_12705_), .B(_12751_), .Y(_12752_));
NAND_g _19268_ (.A(_11170_), .B(_12752_), .Y(_12753_));
NAND_g _19269_ (.A(decoded_imm[20]), .B(_10606_), .Y(_12754_));
AND_g _19270_ (.A(_10603_), .B(_12754_), .Y(_12755_));
NAND_g _19271_ (.A(_12753_), .B(_12755_), .Y(_12756_));
AND_g _19272_ (.A(_12659_), .B(_12756_), .Y(_00295_));
NAND_g _19273_ (.A(_08831_), .B(_10604_), .Y(_12757_));
NAND_g _19274_ (.A(cpuregs[22][21]), .B(_00007_[1]), .Y(_12758_));
NAND_g _19275_ (.A(cpuregs[20][21]), .B(_09026_), .Y(_12759_));
NAND_g _19276_ (.A(_12758_), .B(_12759_), .Y(_12760_));
NAND_g _19277_ (.A(_00007_[2]), .B(_12760_), .Y(_12761_));
NAND_g _19278_ (.A(cpuregs[18][21]), .B(_00007_[1]), .Y(_12762_));
NAND_g _19279_ (.A(cpuregs[16][21]), .B(_09026_), .Y(_12763_));
NAND_g _19280_ (.A(_12762_), .B(_12763_), .Y(_12764_));
NAND_g _19281_ (.A(_09027_), .B(_12764_), .Y(_12765_));
NAND_g _19282_ (.A(_12761_), .B(_12765_), .Y(_12766_));
AND_g _19283_ (.A(_09025_), .B(_12766_), .Y(_12767_));
NOT_g _19284_ (.A(_12767_), .Y(_12768_));
NAND_g _19285_ (.A(cpuregs[23][21]), .B(_00007_[1]), .Y(_12769_));
NAND_g _19286_ (.A(cpuregs[21][21]), .B(_09026_), .Y(_12770_));
NAND_g _19287_ (.A(_12769_), .B(_12770_), .Y(_12771_));
NAND_g _19288_ (.A(_00007_[2]), .B(_12771_), .Y(_12772_));
NAND_g _19289_ (.A(cpuregs[19][21]), .B(_00007_[1]), .Y(_12773_));
NAND_g _19290_ (.A(cpuregs[17][21]), .B(_09026_), .Y(_12774_));
NAND_g _19291_ (.A(_12773_), .B(_12774_), .Y(_12775_));
NAND_g _19292_ (.A(_09027_), .B(_12775_), .Y(_12776_));
NAND_g _19293_ (.A(_12772_), .B(_12776_), .Y(_12777_));
NAND_g _19294_ (.A(_00007_[0]), .B(_12777_), .Y(_12778_));
AND_g _19295_ (.A(_09028_), .B(_12778_), .Y(_12779_));
NAND_g _19296_ (.A(_12768_), .B(_12779_), .Y(_12780_));
NAND_g _19297_ (.A(cpuregs[31][21]), .B(_00007_[2]), .Y(_12781_));
NAND_g _19298_ (.A(cpuregs[27][21]), .B(_09027_), .Y(_12782_));
AND_g _19299_ (.A(_00007_[0]), .B(_12782_), .Y(_12783_));
NAND_g _19300_ (.A(_12781_), .B(_12783_), .Y(_12784_));
NAND_g _19301_ (.A(cpuregs[26][21]), .B(_09027_), .Y(_12785_));
NAND_g _19302_ (.A(cpuregs[30][21]), .B(_00007_[2]), .Y(_12786_));
AND_g _19303_ (.A(_09025_), .B(_12786_), .Y(_12787_));
NAND_g _19304_ (.A(_12785_), .B(_12787_), .Y(_12788_));
AND_g _19305_ (.A(_00007_[1]), .B(_12788_), .Y(_12789_));
NAND_g _19306_ (.A(_12784_), .B(_12789_), .Y(_12790_));
NAND_g _19307_ (.A(cpuregs[25][21]), .B(_09027_), .Y(_12791_));
NAND_g _19308_ (.A(cpuregs[29][21]), .B(_00007_[2]), .Y(_12792_));
AND_g _19309_ (.A(_00007_[0]), .B(_12792_), .Y(_12793_));
NAND_g _19310_ (.A(_12791_), .B(_12793_), .Y(_12794_));
NAND_g _19311_ (.A(cpuregs[24][21]), .B(_09027_), .Y(_12795_));
NAND_g _19312_ (.A(cpuregs[28][21]), .B(_00007_[2]), .Y(_12796_));
AND_g _19313_ (.A(_09025_), .B(_12796_), .Y(_12797_));
NAND_g _19314_ (.A(_12795_), .B(_12797_), .Y(_12798_));
AND_g _19315_ (.A(_09026_), .B(_12798_), .Y(_12799_));
NAND_g _19316_ (.A(_12794_), .B(_12799_), .Y(_12800_));
AND_g _19317_ (.A(_00007_[3]), .B(_12800_), .Y(_12801_));
NAND_g _19318_ (.A(_12790_), .B(_12801_), .Y(_12802_));
NAND_g _19319_ (.A(_12780_), .B(_12802_), .Y(_12803_));
AND_g _19320_ (.A(_00007_[4]), .B(_12803_), .Y(_12804_));
NAND_g _19321_ (.A(cpuregs[3][21]), .B(_09027_), .Y(_12805_));
NAND_g _19322_ (.A(cpuregs[7][21]), .B(_00007_[2]), .Y(_12806_));
AND_g _19323_ (.A(_00007_[0]), .B(_12806_), .Y(_12807_));
NAND_g _19324_ (.A(_12805_), .B(_12807_), .Y(_12808_));
NAND_g _19325_ (.A(cpuregs[2][21]), .B(_09027_), .Y(_12809_));
NAND_g _19326_ (.A(cpuregs[6][21]), .B(_00007_[2]), .Y(_12810_));
AND_g _19327_ (.A(_09025_), .B(_12810_), .Y(_12811_));
NAND_g _19328_ (.A(_12809_), .B(_12811_), .Y(_12812_));
AND_g _19329_ (.A(_00007_[1]), .B(_12812_), .Y(_12813_));
NAND_g _19330_ (.A(_12808_), .B(_12813_), .Y(_12814_));
NAND_g _19331_ (.A(cpuregs[1][21]), .B(_09027_), .Y(_12815_));
NAND_g _19332_ (.A(cpuregs[5][21]), .B(_00007_[2]), .Y(_12816_));
AND_g _19333_ (.A(_00007_[0]), .B(_12816_), .Y(_12817_));
NAND_g _19334_ (.A(_12815_), .B(_12817_), .Y(_12818_));
NAND_g _19335_ (.A(cpuregs[0][21]), .B(_09027_), .Y(_12819_));
NAND_g _19336_ (.A(cpuregs[4][21]), .B(_00007_[2]), .Y(_12820_));
AND_g _19337_ (.A(_09025_), .B(_12820_), .Y(_12821_));
NAND_g _19338_ (.A(_12819_), .B(_12821_), .Y(_12822_));
AND_g _19339_ (.A(_09026_), .B(_12822_), .Y(_12823_));
NAND_g _19340_ (.A(_12818_), .B(_12823_), .Y(_12824_));
AND_g _19341_ (.A(_09028_), .B(_12824_), .Y(_12825_));
NAND_g _19342_ (.A(_12814_), .B(_12825_), .Y(_12826_));
NAND_g _19343_ (.A(cpuregs[12][21]), .B(_09025_), .Y(_12827_));
NAND_g _19344_ (.A(cpuregs[13][21]), .B(_00007_[0]), .Y(_12828_));
NAND_g _19345_ (.A(_12827_), .B(_12828_), .Y(_12829_));
NAND_g _19346_ (.A(_00007_[2]), .B(_12829_), .Y(_12830_));
NAND_g _19347_ (.A(cpuregs[8][21]), .B(_09025_), .Y(_12831_));
NAND_g _19348_ (.A(cpuregs[9][21]), .B(_00007_[0]), .Y(_12832_));
NAND_g _19349_ (.A(_12831_), .B(_12832_), .Y(_12833_));
NAND_g _19350_ (.A(_09027_), .B(_12833_), .Y(_12834_));
NAND_g _19351_ (.A(_12830_), .B(_12834_), .Y(_12835_));
NAND_g _19352_ (.A(_09026_), .B(_12835_), .Y(_12836_));
NAND_g _19353_ (.A(cpuregs[14][21]), .B(_09025_), .Y(_12837_));
NAND_g _19354_ (.A(cpuregs[15][21]), .B(_00007_[0]), .Y(_12838_));
NAND_g _19355_ (.A(_12837_), .B(_12838_), .Y(_12839_));
NAND_g _19356_ (.A(_00007_[2]), .B(_12839_), .Y(_12840_));
NAND_g _19357_ (.A(cpuregs[10][21]), .B(_09025_), .Y(_12841_));
NAND_g _19358_ (.A(cpuregs[11][21]), .B(_00007_[0]), .Y(_12842_));
NAND_g _19359_ (.A(_12841_), .B(_12842_), .Y(_12843_));
NAND_g _19360_ (.A(_09027_), .B(_12843_), .Y(_12844_));
NAND_g _19361_ (.A(_12840_), .B(_12844_), .Y(_12845_));
NAND_g _19362_ (.A(_00007_[1]), .B(_12845_), .Y(_12846_));
AND_g _19363_ (.A(_00007_[3]), .B(_12846_), .Y(_12847_));
NAND_g _19364_ (.A(_12836_), .B(_12847_), .Y(_12848_));
NAND_g _19365_ (.A(_12826_), .B(_12848_), .Y(_12849_));
AND_g _19366_ (.A(_09029_), .B(_12849_), .Y(_12850_));
NOR_g _19367_ (.A(_12804_), .B(_12850_), .Y(_12851_));
NAND_g _19368_ (.A(_11170_), .B(_12851_), .Y(_12852_));
NAND_g _19369_ (.A(decoded_imm[21]), .B(_10606_), .Y(_12853_));
AND_g _19370_ (.A(_10603_), .B(_12853_), .Y(_12854_));
NAND_g _19371_ (.A(_12852_), .B(_12854_), .Y(_12855_));
AND_g _19372_ (.A(_12757_), .B(_12855_), .Y(_00296_));
NAND_g _19373_ (.A(_08832_), .B(_10604_), .Y(_12856_));
NAND_g _19374_ (.A(cpuregs[9][22]), .B(_09027_), .Y(_12857_));
NAND_g _19375_ (.A(cpuregs[13][22]), .B(_00007_[2]), .Y(_12858_));
NAND_g _19376_ (.A(_12857_), .B(_12858_), .Y(_12859_));
NAND_g _19377_ (.A(_00007_[0]), .B(_12859_), .Y(_12860_));
NAND_g _19378_ (.A(cpuregs[12][22]), .B(_00007_[2]), .Y(_12861_));
NAND_g _19379_ (.A(cpuregs[8][22]), .B(_09027_), .Y(_12862_));
NAND_g _19380_ (.A(_12861_), .B(_12862_), .Y(_12863_));
NAND_g _19381_ (.A(_09025_), .B(_12863_), .Y(_12864_));
NAND_g _19382_ (.A(_12860_), .B(_12864_), .Y(_12865_));
NAND_g _19383_ (.A(_09026_), .B(_12865_), .Y(_12866_));
NAND_g _19384_ (.A(cpuregs[11][22]), .B(_09027_), .Y(_12867_));
NAND_g _19385_ (.A(cpuregs[15][22]), .B(_00007_[2]), .Y(_12868_));
NAND_g _19386_ (.A(_12867_), .B(_12868_), .Y(_12869_));
NAND_g _19387_ (.A(_00007_[0]), .B(_12869_), .Y(_12870_));
NAND_g _19388_ (.A(cpuregs[14][22]), .B(_00007_[2]), .Y(_12871_));
NAND_g _19389_ (.A(cpuregs[10][22]), .B(_09027_), .Y(_12872_));
NAND_g _19390_ (.A(_12871_), .B(_12872_), .Y(_12873_));
NAND_g _19391_ (.A(_09025_), .B(_12873_), .Y(_12874_));
NAND_g _19392_ (.A(_12870_), .B(_12874_), .Y(_12875_));
NAND_g _19393_ (.A(_00007_[1]), .B(_12875_), .Y(_12876_));
NAND_g _19394_ (.A(cpuregs[31][22]), .B(_00007_[2]), .Y(_12877_));
NAND_g _19395_ (.A(cpuregs[27][22]), .B(_09027_), .Y(_12878_));
AND_g _19396_ (.A(_00007_[0]), .B(_12878_), .Y(_12879_));
NAND_g _19397_ (.A(_12877_), .B(_12879_), .Y(_12880_));
NAND_g _19398_ (.A(cpuregs[26][22]), .B(_09027_), .Y(_12881_));
NAND_g _19399_ (.A(cpuregs[30][22]), .B(_00007_[2]), .Y(_12882_));
AND_g _19400_ (.A(_09025_), .B(_12882_), .Y(_12883_));
NAND_g _19401_ (.A(_12881_), .B(_12883_), .Y(_12884_));
AND_g _19402_ (.A(_00007_[1]), .B(_12884_), .Y(_12885_));
NAND_g _19403_ (.A(_12880_), .B(_12885_), .Y(_12886_));
NAND_g _19404_ (.A(cpuregs[29][22]), .B(_00007_[2]), .Y(_12887_));
NAND_g _19405_ (.A(cpuregs[25][22]), .B(_09027_), .Y(_12888_));
AND_g _19406_ (.A(_00007_[0]), .B(_12888_), .Y(_12889_));
NAND_g _19407_ (.A(_12887_), .B(_12889_), .Y(_12890_));
NAND_g _19408_ (.A(cpuregs[24][22]), .B(_09027_), .Y(_12891_));
NAND_g _19409_ (.A(cpuregs[28][22]), .B(_00007_[2]), .Y(_12892_));
AND_g _19410_ (.A(_09025_), .B(_12892_), .Y(_12893_));
NAND_g _19411_ (.A(_12891_), .B(_12893_), .Y(_12894_));
AND_g _19412_ (.A(_09026_), .B(_12894_), .Y(_12895_));
NAND_g _19413_ (.A(_12890_), .B(_12895_), .Y(_12896_));
NAND_g _19414_ (.A(cpuregs[1][22]), .B(_09027_), .Y(_12897_));
NAND_g _19415_ (.A(cpuregs[5][22]), .B(_00007_[2]), .Y(_12898_));
NAND_g _19416_ (.A(_12897_), .B(_12898_), .Y(_12899_));
NAND_g _19417_ (.A(_00007_[0]), .B(_12899_), .Y(_12900_));
NAND_g _19418_ (.A(cpuregs[4][22]), .B(_00007_[2]), .Y(_12901_));
NAND_g _19419_ (.A(cpuregs[0][22]), .B(_09027_), .Y(_12902_));
NAND_g _19420_ (.A(_12901_), .B(_12902_), .Y(_12903_));
NAND_g _19421_ (.A(_09025_), .B(_12903_), .Y(_12904_));
NAND_g _19422_ (.A(_12900_), .B(_12904_), .Y(_12905_));
NAND_g _19423_ (.A(_09026_), .B(_12905_), .Y(_12906_));
NAND_g _19424_ (.A(cpuregs[6][22]), .B(_00007_[2]), .Y(_12907_));
NAND_g _19425_ (.A(cpuregs[2][22]), .B(_09027_), .Y(_12908_));
NAND_g _19426_ (.A(_12907_), .B(_12908_), .Y(_12909_));
NAND_g _19427_ (.A(_09025_), .B(_12909_), .Y(_12910_));
NOR_g _19428_ (.A(cpuregs[3][22]), .B(_00007_[2]), .Y(_12911_));
NAND_g _19429_ (.A(_08976_), .B(_00007_[2]), .Y(_12912_));
NOR_g _19430_ (.A(_09025_), .B(_12911_), .Y(_12913_));
NAND_g _19431_ (.A(_12912_), .B(_12913_), .Y(_12914_));
NAND_g _19432_ (.A(_12910_), .B(_12914_), .Y(_12915_));
NAND_g _19433_ (.A(_00007_[1]), .B(_12915_), .Y(_12916_));
NAND_g _19434_ (.A(_08937_), .B(_09027_), .Y(_12917_));
NOR_g _19435_ (.A(cpuregs[22][22]), .B(_09027_), .Y(_12918_));
NAND_g _19436_ (.A(_08898_), .B(_00007_[2]), .Y(_12919_));
NOR_g _19437_ (.A(cpuregs[19][22]), .B(_00007_[2]), .Y(_12920_));
NOR_g _19438_ (.A(_00007_[0]), .B(_12918_), .Y(_12921_));
AND_g _19439_ (.A(_12917_), .B(_12921_), .Y(_12922_));
NAND_g _19440_ (.A(_00007_[0]), .B(_12919_), .Y(_12923_));
NOR_g _19441_ (.A(_12920_), .B(_12923_), .Y(_12924_));
NOR_g _19442_ (.A(_12922_), .B(_12924_), .Y(_12925_));
NOR_g _19443_ (.A(cpuregs[16][22]), .B(_00007_[2]), .Y(_12926_));
NOR_g _19444_ (.A(cpuregs[20][22]), .B(_09027_), .Y(_12927_));
NOR_g _19445_ (.A(_12926_), .B(_12927_), .Y(_12928_));
NOR_g _19446_ (.A(cpuregs[17][22]), .B(_00007_[2]), .Y(_12929_));
NAND_g _19447_ (.A(_08997_), .B(_00007_[2]), .Y(_12930_));
NAND_g _19448_ (.A(_00007_[0]), .B(_12930_), .Y(_12931_));
NOR_g _19449_ (.A(_12929_), .B(_12931_), .Y(_12932_));
AND_g _19450_ (.A(_09025_), .B(_12928_), .Y(_12933_));
NOR_g _19451_ (.A(_12932_), .B(_12933_), .Y(_12934_));
NAND_g _19452_ (.A(_00007_[1]), .B(_12925_), .Y(_12935_));
NAND_g _19453_ (.A(_09026_), .B(_12934_), .Y(_12936_));
AND_g _19454_ (.A(_12935_), .B(_12936_), .Y(_12937_));
NAND_g _19455_ (.A(_09028_), .B(_12937_), .Y(_12938_));
NAND_g _19456_ (.A(_12886_), .B(_12896_), .Y(_12939_));
NAND_g _19457_ (.A(_00007_[3]), .B(_12939_), .Y(_12940_));
AND_g _19458_ (.A(_00007_[4]), .B(_12940_), .Y(_12941_));
NAND_g _19459_ (.A(_12938_), .B(_12941_), .Y(_12942_));
NAND_g _19460_ (.A(_12906_), .B(_12916_), .Y(_12943_));
NAND_g _19461_ (.A(_09028_), .B(_12943_), .Y(_12944_));
NAND_g _19462_ (.A(_12866_), .B(_12876_), .Y(_12945_));
NAND_g _19463_ (.A(_00007_[3]), .B(_12945_), .Y(_12946_));
AND_g _19464_ (.A(_12944_), .B(_12946_), .Y(_12947_));
NAND_g _19465_ (.A(_09029_), .B(_12947_), .Y(_12948_));
AND_g _19466_ (.A(_12942_), .B(_12948_), .Y(_12949_));
NAND_g _19467_ (.A(_11170_), .B(_12949_), .Y(_12950_));
NAND_g _19468_ (.A(decoded_imm[22]), .B(_10606_), .Y(_12951_));
AND_g _19469_ (.A(_10603_), .B(_12951_), .Y(_12952_));
NAND_g _19470_ (.A(_12950_), .B(_12952_), .Y(_12953_));
AND_g _19471_ (.A(_12856_), .B(_12953_), .Y(_00297_));
NAND_g _19472_ (.A(_08833_), .B(_10604_), .Y(_12954_));
NAND_g _19473_ (.A(cpuregs[9][23]), .B(_09027_), .Y(_12955_));
NAND_g _19474_ (.A(cpuregs[13][23]), .B(_00007_[2]), .Y(_12956_));
NAND_g _19475_ (.A(_12955_), .B(_12956_), .Y(_12957_));
NAND_g _19476_ (.A(_00007_[0]), .B(_12957_), .Y(_12958_));
NAND_g _19477_ (.A(cpuregs[12][23]), .B(_00007_[2]), .Y(_12959_));
NAND_g _19478_ (.A(cpuregs[8][23]), .B(_09027_), .Y(_12960_));
NAND_g _19479_ (.A(_12959_), .B(_12960_), .Y(_12961_));
NAND_g _19480_ (.A(_09025_), .B(_12961_), .Y(_12962_));
NAND_g _19481_ (.A(_12958_), .B(_12962_), .Y(_12963_));
NAND_g _19482_ (.A(_09026_), .B(_12963_), .Y(_12964_));
NAND_g _19483_ (.A(cpuregs[11][23]), .B(_09027_), .Y(_12965_));
NAND_g _19484_ (.A(cpuregs[15][23]), .B(_00007_[2]), .Y(_12966_));
NAND_g _19485_ (.A(_12965_), .B(_12966_), .Y(_12967_));
NAND_g _19486_ (.A(_00007_[0]), .B(_12967_), .Y(_12968_));
NAND_g _19487_ (.A(cpuregs[14][23]), .B(_00007_[2]), .Y(_12969_));
NAND_g _19488_ (.A(cpuregs[10][23]), .B(_09027_), .Y(_12970_));
NAND_g _19489_ (.A(_12969_), .B(_12970_), .Y(_12971_));
NAND_g _19490_ (.A(_09025_), .B(_12971_), .Y(_12972_));
NAND_g _19491_ (.A(_12968_), .B(_12972_), .Y(_12973_));
NAND_g _19492_ (.A(_00007_[1]), .B(_12973_), .Y(_12974_));
NAND_g _19493_ (.A(cpuregs[31][23]), .B(_00007_[2]), .Y(_12975_));
NAND_g _19494_ (.A(cpuregs[27][23]), .B(_09027_), .Y(_12976_));
AND_g _19495_ (.A(_00007_[0]), .B(_12976_), .Y(_12977_));
NAND_g _19496_ (.A(_12975_), .B(_12977_), .Y(_12978_));
NAND_g _19497_ (.A(cpuregs[26][23]), .B(_09027_), .Y(_12979_));
NAND_g _19498_ (.A(cpuregs[30][23]), .B(_00007_[2]), .Y(_12980_));
AND_g _19499_ (.A(_09025_), .B(_12980_), .Y(_12981_));
NAND_g _19500_ (.A(_12979_), .B(_12981_), .Y(_12982_));
AND_g _19501_ (.A(_00007_[1]), .B(_12982_), .Y(_12983_));
NAND_g _19502_ (.A(_12978_), .B(_12983_), .Y(_12984_));
NAND_g _19503_ (.A(cpuregs[29][23]), .B(_00007_[2]), .Y(_12985_));
NAND_g _19504_ (.A(cpuregs[25][23]), .B(_09027_), .Y(_12986_));
AND_g _19505_ (.A(_00007_[0]), .B(_12986_), .Y(_12987_));
NAND_g _19506_ (.A(_12985_), .B(_12987_), .Y(_12988_));
NAND_g _19507_ (.A(cpuregs[24][23]), .B(_09027_), .Y(_12989_));
NAND_g _19508_ (.A(cpuregs[28][23]), .B(_00007_[2]), .Y(_12990_));
AND_g _19509_ (.A(_09025_), .B(_12990_), .Y(_12991_));
NAND_g _19510_ (.A(_12989_), .B(_12991_), .Y(_12992_));
AND_g _19511_ (.A(_09026_), .B(_12992_), .Y(_12993_));
NAND_g _19512_ (.A(_12988_), .B(_12993_), .Y(_12994_));
NAND_g _19513_ (.A(cpuregs[1][23]), .B(_09027_), .Y(_12995_));
NAND_g _19514_ (.A(cpuregs[5][23]), .B(_00007_[2]), .Y(_12996_));
NAND_g _19515_ (.A(_12995_), .B(_12996_), .Y(_12997_));
NAND_g _19516_ (.A(_00007_[0]), .B(_12997_), .Y(_12998_));
NAND_g _19517_ (.A(cpuregs[4][23]), .B(_00007_[2]), .Y(_12999_));
NAND_g _19518_ (.A(cpuregs[0][23]), .B(_09027_), .Y(_13000_));
NAND_g _19519_ (.A(_12999_), .B(_13000_), .Y(_13001_));
NAND_g _19520_ (.A(_09025_), .B(_13001_), .Y(_13002_));
NAND_g _19521_ (.A(_12998_), .B(_13002_), .Y(_13003_));
NAND_g _19522_ (.A(_09026_), .B(_13003_), .Y(_13004_));
NAND_g _19523_ (.A(cpuregs[6][23]), .B(_00007_[2]), .Y(_13005_));
NAND_g _19524_ (.A(cpuregs[2][23]), .B(_09027_), .Y(_13006_));
NAND_g _19525_ (.A(_13005_), .B(_13006_), .Y(_13007_));
NAND_g _19526_ (.A(_09025_), .B(_13007_), .Y(_13008_));
NAND_g _19527_ (.A(cpuregs[7][23]), .B(_00007_[2]), .Y(_13009_));
NAND_g _19528_ (.A(cpuregs[3][23]), .B(_09027_), .Y(_13010_));
NAND_g _19529_ (.A(_13009_), .B(_13010_), .Y(_13011_));
NAND_g _19530_ (.A(_00007_[0]), .B(_13011_), .Y(_13012_));
NAND_g _19531_ (.A(_13008_), .B(_13012_), .Y(_13013_));
NAND_g _19532_ (.A(_00007_[1]), .B(_13013_), .Y(_13014_));
NOR_g _19533_ (.A(cpuregs[18][23]), .B(_00007_[2]), .Y(_13015_));
NAND_g _19534_ (.A(_08924_), .B(_00007_[2]), .Y(_13016_));
NAND_g _19535_ (.A(_08899_), .B(_00007_[2]), .Y(_13017_));
NOR_g _19536_ (.A(cpuregs[19][23]), .B(_00007_[2]), .Y(_13018_));
NAND_g _19537_ (.A(_09025_), .B(_13016_), .Y(_13019_));
NOR_g _19538_ (.A(_13015_), .B(_13019_), .Y(_13020_));
NAND_g _19539_ (.A(_00007_[0]), .B(_13017_), .Y(_13021_));
NOR_g _19540_ (.A(_13018_), .B(_13021_), .Y(_13022_));
NOR_g _19541_ (.A(_13020_), .B(_13022_), .Y(_13023_));
NOR_g _19542_ (.A(cpuregs[16][23]), .B(_00007_[2]), .Y(_13024_));
AND_g _19543_ (.A(_08850_), .B(_00007_[2]), .Y(_13025_));
NOR_g _19544_ (.A(_13024_), .B(_13025_), .Y(_13026_));
NOR_g _19545_ (.A(cpuregs[17][23]), .B(_00007_[2]), .Y(_13027_));
NAND_g _19546_ (.A(_08998_), .B(_00007_[2]), .Y(_13028_));
NAND_g _19547_ (.A(_00007_[0]), .B(_13028_), .Y(_13029_));
NOR_g _19548_ (.A(_13027_), .B(_13029_), .Y(_13030_));
AND_g _19549_ (.A(_09025_), .B(_13026_), .Y(_13031_));
NOR_g _19550_ (.A(_13030_), .B(_13031_), .Y(_13032_));
NAND_g _19551_ (.A(_00007_[1]), .B(_13023_), .Y(_13033_));
NAND_g _19552_ (.A(_09026_), .B(_13032_), .Y(_13034_));
AND_g _19553_ (.A(_09028_), .B(_13034_), .Y(_13035_));
NAND_g _19554_ (.A(_13033_), .B(_13035_), .Y(_13036_));
NAND_g _19555_ (.A(_12984_), .B(_12994_), .Y(_13037_));
NAND_g _19556_ (.A(_00007_[3]), .B(_13037_), .Y(_13038_));
AND_g _19557_ (.A(_00007_[4]), .B(_13038_), .Y(_13039_));
NAND_g _19558_ (.A(_13036_), .B(_13039_), .Y(_13040_));
NAND_g _19559_ (.A(_12964_), .B(_12974_), .Y(_13041_));
NAND_g _19560_ (.A(_00007_[3]), .B(_13041_), .Y(_13042_));
NAND_g _19561_ (.A(_13004_), .B(_13014_), .Y(_13043_));
NAND_g _19562_ (.A(_09028_), .B(_13043_), .Y(_13044_));
AND_g _19563_ (.A(_13042_), .B(_13044_), .Y(_13045_));
NAND_g _19564_ (.A(_09029_), .B(_13045_), .Y(_13046_));
AND_g _19565_ (.A(_13040_), .B(_13046_), .Y(_13047_));
NAND_g _19566_ (.A(_11170_), .B(_13047_), .Y(_13048_));
NAND_g _19567_ (.A(decoded_imm[23]), .B(_10606_), .Y(_13049_));
AND_g _19568_ (.A(_10603_), .B(_13049_), .Y(_13050_));
NAND_g _19569_ (.A(_13048_), .B(_13050_), .Y(_13051_));
AND_g _19570_ (.A(_12954_), .B(_13051_), .Y(_00298_));
NAND_g _19571_ (.A(_08834_), .B(_10604_), .Y(_13052_));
NAND_g _19572_ (.A(cpuregs[18][24]), .B(_00007_[1]), .Y(_13053_));
NAND_g _19573_ (.A(cpuregs[16][24]), .B(_09026_), .Y(_13054_));
NAND_g _19574_ (.A(_13053_), .B(_13054_), .Y(_13055_));
NAND_g _19575_ (.A(_09027_), .B(_13055_), .Y(_13056_));
NAND_g _19576_ (.A(cpuregs[22][24]), .B(_00007_[1]), .Y(_13057_));
NAND_g _19577_ (.A(cpuregs[20][24]), .B(_09026_), .Y(_13058_));
NAND_g _19578_ (.A(_13057_), .B(_13058_), .Y(_13059_));
NAND_g _19579_ (.A(_00007_[2]), .B(_13059_), .Y(_13060_));
AND_g _19580_ (.A(_09025_), .B(_13060_), .Y(_13061_));
NAND_g _19581_ (.A(_13056_), .B(_13061_), .Y(_13062_));
NAND_g _19582_ (.A(cpuregs[19][24]), .B(_00007_[1]), .Y(_13063_));
NAND_g _19583_ (.A(cpuregs[17][24]), .B(_09026_), .Y(_13064_));
NAND_g _19584_ (.A(_13063_), .B(_13064_), .Y(_13065_));
NAND_g _19585_ (.A(_09027_), .B(_13065_), .Y(_13066_));
NAND_g _19586_ (.A(cpuregs[23][24]), .B(_00007_[1]), .Y(_13067_));
NAND_g _19587_ (.A(cpuregs[21][24]), .B(_09026_), .Y(_13068_));
NAND_g _19588_ (.A(_13067_), .B(_13068_), .Y(_13069_));
NAND_g _19589_ (.A(_00007_[2]), .B(_13069_), .Y(_13070_));
AND_g _19590_ (.A(_00007_[0]), .B(_13070_), .Y(_13071_));
NAND_g _19591_ (.A(_13066_), .B(_13071_), .Y(_13072_));
AND_g _19592_ (.A(_13062_), .B(_13072_), .Y(_13073_));
NAND_g _19593_ (.A(cpuregs[26][24]), .B(_09027_), .Y(_13074_));
NAND_g _19594_ (.A(cpuregs[30][24]), .B(_00007_[2]), .Y(_13075_));
AND_g _19595_ (.A(_09025_), .B(_13075_), .Y(_13076_));
NAND_g _19596_ (.A(_13074_), .B(_13076_), .Y(_13077_));
NAND_g _19597_ (.A(cpuregs[31][24]), .B(_00007_[2]), .Y(_13078_));
NAND_g _19598_ (.A(cpuregs[27][24]), .B(_09027_), .Y(_13079_));
AND_g _19599_ (.A(_00007_[0]), .B(_13079_), .Y(_13080_));
NAND_g _19600_ (.A(_13078_), .B(_13080_), .Y(_13081_));
NAND_g _19601_ (.A(_13077_), .B(_13081_), .Y(_13082_));
NAND_g _19602_ (.A(_00007_[1]), .B(_13082_), .Y(_13083_));
NAND_g _19603_ (.A(cpuregs[24][24]), .B(_09027_), .Y(_13084_));
NAND_g _19604_ (.A(cpuregs[28][24]), .B(_00007_[2]), .Y(_13085_));
AND_g _19605_ (.A(_09025_), .B(_13085_), .Y(_13086_));
NAND_g _19606_ (.A(_13084_), .B(_13086_), .Y(_13087_));
NAND_g _19607_ (.A(cpuregs[25][24]), .B(_09027_), .Y(_13088_));
NAND_g _19608_ (.A(cpuregs[29][24]), .B(_00007_[2]), .Y(_13089_));
AND_g _19609_ (.A(_00007_[0]), .B(_13089_), .Y(_13090_));
NAND_g _19610_ (.A(_13088_), .B(_13090_), .Y(_13091_));
NAND_g _19611_ (.A(_13087_), .B(_13091_), .Y(_13092_));
NAND_g _19612_ (.A(_09026_), .B(_13092_), .Y(_13093_));
AND_g _19613_ (.A(_00007_[3]), .B(_13093_), .Y(_13094_));
NAND_g _19614_ (.A(_13083_), .B(_13094_), .Y(_13095_));
NAND_g _19615_ (.A(_09028_), .B(_13073_), .Y(_13096_));
AND_g _19616_ (.A(_00007_[4]), .B(_13095_), .Y(_13097_));
AND_g _19617_ (.A(_13096_), .B(_13097_), .Y(_13098_));
NAND_g _19618_ (.A(_08977_), .B(_00007_[2]), .Y(_13099_));
NOR_g _19619_ (.A(cpuregs[3][24]), .B(_00007_[2]), .Y(_13100_));
NOR_g _19620_ (.A(cpuregs[2][24]), .B(_00007_[2]), .Y(_13101_));
NOR_g _19621_ (.A(cpuregs[6][24]), .B(_09027_), .Y(_13102_));
NOR_g _19622_ (.A(_13101_), .B(_13102_), .Y(_13103_));
NOR_g _19623_ (.A(_09025_), .B(_13100_), .Y(_13104_));
NAND_g _19624_ (.A(_13099_), .B(_13104_), .Y(_13105_));
NAND_g _19625_ (.A(_09025_), .B(_13103_), .Y(_13106_));
AND_g _19626_ (.A(_13105_), .B(_13106_), .Y(_13107_));
NAND_g _19627_ (.A(_00007_[1]), .B(_13107_), .Y(_13108_));
NOR_g _19628_ (.A(cpuregs[1][24]), .B(_00007_[2]), .Y(_13109_));
NAND_g _19629_ (.A(_08959_), .B(_00007_[2]), .Y(_13110_));
NOR_g _19630_ (.A(cpuregs[0][24]), .B(_00007_[2]), .Y(_13111_));
NOR_g _19631_ (.A(cpuregs[4][24]), .B(_09027_), .Y(_13112_));
NOR_g _19632_ (.A(_13111_), .B(_13112_), .Y(_13113_));
NOR_g _19633_ (.A(_09025_), .B(_13109_), .Y(_13114_));
NAND_g _19634_ (.A(_13110_), .B(_13114_), .Y(_13115_));
NAND_g _19635_ (.A(_09025_), .B(_13113_), .Y(_13116_));
AND_g _19636_ (.A(_13115_), .B(_13116_), .Y(_13117_));
NAND_g _19637_ (.A(_09026_), .B(_13117_), .Y(_13118_));
NAND_g _19638_ (.A(_13108_), .B(_13118_), .Y(_13119_));
NAND_g _19639_ (.A(_09028_), .B(_13119_), .Y(_13120_));
NAND_g _19640_ (.A(cpuregs[9][24]), .B(_09026_), .Y(_13121_));
NAND_g _19641_ (.A(cpuregs[11][24]), .B(_00007_[1]), .Y(_13122_));
AND_g _19642_ (.A(_09027_), .B(_13122_), .Y(_13123_));
NAND_g _19643_ (.A(_13121_), .B(_13123_), .Y(_13124_));
NAND_g _19644_ (.A(cpuregs[13][24]), .B(_09026_), .Y(_13125_));
NAND_g _19645_ (.A(cpuregs[15][24]), .B(_00007_[1]), .Y(_13126_));
AND_g _19646_ (.A(_00007_[2]), .B(_13126_), .Y(_13127_));
NAND_g _19647_ (.A(_13125_), .B(_13127_), .Y(_13128_));
NAND_g _19648_ (.A(_13124_), .B(_13128_), .Y(_13129_));
NAND_g _19649_ (.A(_00007_[0]), .B(_13129_), .Y(_13130_));
NAND_g _19650_ (.A(cpuregs[8][24]), .B(_09026_), .Y(_13131_));
NAND_g _19651_ (.A(cpuregs[10][24]), .B(_00007_[1]), .Y(_13132_));
AND_g _19652_ (.A(_09027_), .B(_13132_), .Y(_13133_));
NAND_g _19653_ (.A(_13131_), .B(_13133_), .Y(_13134_));
NAND_g _19654_ (.A(cpuregs[12][24]), .B(_09026_), .Y(_13135_));
NAND_g _19655_ (.A(cpuregs[14][24]), .B(_00007_[1]), .Y(_13136_));
AND_g _19656_ (.A(_00007_[2]), .B(_13136_), .Y(_13137_));
NAND_g _19657_ (.A(_13135_), .B(_13137_), .Y(_13138_));
NAND_g _19658_ (.A(_13134_), .B(_13138_), .Y(_13139_));
NAND_g _19659_ (.A(_09025_), .B(_13139_), .Y(_13140_));
NAND_g _19660_ (.A(_13130_), .B(_13140_), .Y(_13141_));
NAND_g _19661_ (.A(_00007_[3]), .B(_13141_), .Y(_13142_));
NAND_g _19662_ (.A(_13120_), .B(_13142_), .Y(_13143_));
AND_g _19663_ (.A(_09029_), .B(_13143_), .Y(_13144_));
NOR_g _19664_ (.A(_13098_), .B(_13144_), .Y(_13145_));
NAND_g _19665_ (.A(_11170_), .B(_13145_), .Y(_13146_));
NAND_g _19666_ (.A(decoded_imm[24]), .B(_10606_), .Y(_13147_));
AND_g _19667_ (.A(_10603_), .B(_13147_), .Y(_13148_));
NAND_g _19668_ (.A(_13146_), .B(_13148_), .Y(_13149_));
AND_g _19669_ (.A(_13052_), .B(_13149_), .Y(_00299_));
NAND_g _19670_ (.A(_08835_), .B(_10604_), .Y(_13150_));
NAND_g _19671_ (.A(cpuregs[14][25]), .B(_09025_), .Y(_13151_));
NAND_g _19672_ (.A(cpuregs[15][25]), .B(_00007_[0]), .Y(_13152_));
NAND_g _19673_ (.A(_13151_), .B(_13152_), .Y(_13153_));
NAND_g _19674_ (.A(_00007_[2]), .B(_13153_), .Y(_13154_));
NAND_g _19675_ (.A(cpuregs[10][25]), .B(_09025_), .Y(_13155_));
NAND_g _19676_ (.A(cpuregs[11][25]), .B(_00007_[0]), .Y(_13156_));
NAND_g _19677_ (.A(_13155_), .B(_13156_), .Y(_13157_));
NAND_g _19678_ (.A(_09027_), .B(_13157_), .Y(_13158_));
NAND_g _19679_ (.A(_13154_), .B(_13158_), .Y(_13159_));
NAND_g _19680_ (.A(_00007_[1]), .B(_13159_), .Y(_13160_));
NAND_g _19681_ (.A(_08933_), .B(_00007_[2]), .Y(_13161_));
NOR_g _19682_ (.A(cpuregs[9][25]), .B(_00007_[2]), .Y(_13162_));
NOR_g _19683_ (.A(_09025_), .B(_13162_), .Y(_13163_));
NAND_g _19684_ (.A(_13161_), .B(_13163_), .Y(_13164_));
NOR_g _19685_ (.A(cpuregs[8][25]), .B(_00007_[2]), .Y(_13165_));
AND_g _19686_ (.A(_08883_), .B(_00007_[2]), .Y(_13166_));
NOR_g _19687_ (.A(_13165_), .B(_13166_), .Y(_13167_));
NAND_g _19688_ (.A(_09025_), .B(_13167_), .Y(_13168_));
NAND_g _19689_ (.A(_13164_), .B(_13168_), .Y(_13169_));
NAND_g _19690_ (.A(_09026_), .B(_13169_), .Y(_13170_));
AND_g _19691_ (.A(_09029_), .B(_13170_), .Y(_13171_));
NAND_g _19692_ (.A(_13160_), .B(_13171_), .Y(_13172_));
NAND_g _19693_ (.A(cpuregs[27][25]), .B(_09027_), .Y(_13173_));
NAND_g _19694_ (.A(cpuregs[31][25]), .B(_00007_[2]), .Y(_13174_));
AND_g _19695_ (.A(_00007_[0]), .B(_13174_), .Y(_13175_));
NAND_g _19696_ (.A(_13173_), .B(_13175_), .Y(_13176_));
NAND_g _19697_ (.A(cpuregs[26][25]), .B(_09027_), .Y(_13177_));
NAND_g _19698_ (.A(cpuregs[30][25]), .B(_00007_[2]), .Y(_13178_));
AND_g _19699_ (.A(_09025_), .B(_13178_), .Y(_13179_));
NAND_g _19700_ (.A(_13177_), .B(_13179_), .Y(_13180_));
AND_g _19701_ (.A(_00007_[1]), .B(_13180_), .Y(_13181_));
NAND_g _19702_ (.A(_13176_), .B(_13181_), .Y(_13182_));
NAND_g _19703_ (.A(cpuregs[29][25]), .B(_00007_[2]), .Y(_13183_));
NAND_g _19704_ (.A(cpuregs[25][25]), .B(_09027_), .Y(_13184_));
AND_g _19705_ (.A(_00007_[0]), .B(_13184_), .Y(_13185_));
NAND_g _19706_ (.A(_13183_), .B(_13185_), .Y(_13186_));
NAND_g _19707_ (.A(cpuregs[28][25]), .B(_00007_[2]), .Y(_13187_));
NAND_g _19708_ (.A(cpuregs[24][25]), .B(_09027_), .Y(_13188_));
AND_g _19709_ (.A(_09025_), .B(_13188_), .Y(_13189_));
NAND_g _19710_ (.A(_13187_), .B(_13189_), .Y(_13190_));
AND_g _19711_ (.A(_09026_), .B(_13190_), .Y(_13191_));
NAND_g _19712_ (.A(_13186_), .B(_13191_), .Y(_13192_));
AND_g _19713_ (.A(_00007_[4]), .B(_13192_), .Y(_13193_));
NAND_g _19714_ (.A(_13182_), .B(_13193_), .Y(_13194_));
NAND_g _19715_ (.A(_13172_), .B(_13194_), .Y(_13195_));
AND_g _19716_ (.A(_00007_[3]), .B(_13195_), .Y(_13196_));
NAND_g _19717_ (.A(cpuregs[3][25]), .B(_09027_), .Y(_13197_));
NAND_g _19718_ (.A(cpuregs[7][25]), .B(_00007_[2]), .Y(_13198_));
AND_g _19719_ (.A(_00007_[0]), .B(_13198_), .Y(_13199_));
NAND_g _19720_ (.A(_13197_), .B(_13199_), .Y(_13200_));
NAND_g _19721_ (.A(cpuregs[2][25]), .B(_09027_), .Y(_13201_));
NAND_g _19722_ (.A(cpuregs[6][25]), .B(_00007_[2]), .Y(_13202_));
AND_g _19723_ (.A(_09025_), .B(_13202_), .Y(_13203_));
NAND_g _19724_ (.A(_13201_), .B(_13203_), .Y(_13204_));
AND_g _19725_ (.A(_00007_[1]), .B(_13204_), .Y(_13205_));
NAND_g _19726_ (.A(_13200_), .B(_13205_), .Y(_13206_));
NAND_g _19727_ (.A(cpuregs[1][25]), .B(_09027_), .Y(_13207_));
NAND_g _19728_ (.A(cpuregs[5][25]), .B(_00007_[2]), .Y(_13208_));
AND_g _19729_ (.A(_00007_[0]), .B(_13208_), .Y(_13209_));
NAND_g _19730_ (.A(_13207_), .B(_13209_), .Y(_13210_));
NAND_g _19731_ (.A(cpuregs[0][25]), .B(_09027_), .Y(_13211_));
NAND_g _19732_ (.A(cpuregs[4][25]), .B(_00007_[2]), .Y(_13212_));
AND_g _19733_ (.A(_09025_), .B(_13212_), .Y(_13213_));
NAND_g _19734_ (.A(_13211_), .B(_13213_), .Y(_13214_));
AND_g _19735_ (.A(_09026_), .B(_13214_), .Y(_13215_));
NAND_g _19736_ (.A(_13210_), .B(_13215_), .Y(_13216_));
AND_g _19737_ (.A(_09029_), .B(_13216_), .Y(_13217_));
AND_g _19738_ (.A(_13206_), .B(_13217_), .Y(_13218_));
NOR_g _19739_ (.A(cpuregs[18][25]), .B(_00007_[2]), .Y(_13219_));
AND_g _19740_ (.A(_08925_), .B(_00007_[2]), .Y(_13220_));
NOR_g _19741_ (.A(_13219_), .B(_13220_), .Y(_13221_));
NOR_g _19742_ (.A(_00007_[0]), .B(_13221_), .Y(_13222_));
NAND_g _19743_ (.A(_08900_), .B(_00007_[2]), .Y(_13223_));
NOR_g _19744_ (.A(cpuregs[19][25]), .B(_00007_[2]), .Y(_13224_));
NOT_g _19745_ (.A(_13224_), .Y(_13225_));
NAND_g _19746_ (.A(_13223_), .B(_13225_), .Y(_13226_));
NAND_g _19747_ (.A(_00007_[0]), .B(_13226_), .Y(_13227_));
NAND_g _19748_ (.A(_00007_[1]), .B(_13227_), .Y(_13228_));
NOR_g _19749_ (.A(_13222_), .B(_13228_), .Y(_13229_));
NOR_g _19750_ (.A(cpuregs[16][25]), .B(_00007_[2]), .Y(_13230_));
AND_g _19751_ (.A(_08851_), .B(_00007_[2]), .Y(_13231_));
NOR_g _19752_ (.A(_13230_), .B(_13231_), .Y(_13232_));
NOR_g _19753_ (.A(_00007_[0]), .B(_13232_), .Y(_13233_));
NOT_g _19754_ (.A(_13233_), .Y(_13234_));
NOR_g _19755_ (.A(cpuregs[17][25]), .B(_00007_[2]), .Y(_13235_));
NOT_g _19756_ (.A(_13235_), .Y(_13236_));
NAND_g _19757_ (.A(_08999_), .B(_00007_[2]), .Y(_13237_));
NAND_g _19758_ (.A(_13236_), .B(_13237_), .Y(_13238_));
NAND_g _19759_ (.A(_00007_[0]), .B(_13238_), .Y(_13239_));
AND_g _19760_ (.A(_09026_), .B(_13239_), .Y(_13240_));
NAND_g _19761_ (.A(_13234_), .B(_13240_), .Y(_13241_));
NAND_g _19762_ (.A(_00007_[4]), .B(_13241_), .Y(_13242_));
NOR_g _19763_ (.A(_13229_), .B(_13242_), .Y(_13243_));
NOR_g _19764_ (.A(_13218_), .B(_13243_), .Y(_13244_));
NOR_g _19765_ (.A(_00007_[3]), .B(_13244_), .Y(_13245_));
NOR_g _19766_ (.A(_13196_), .B(_13245_), .Y(_13246_));
NAND_g _19767_ (.A(_11170_), .B(_13246_), .Y(_13247_));
NAND_g _19768_ (.A(decoded_imm[25]), .B(_10606_), .Y(_13248_));
AND_g _19769_ (.A(_10603_), .B(_13248_), .Y(_13249_));
NAND_g _19770_ (.A(_13247_), .B(_13249_), .Y(_13250_));
AND_g _19771_ (.A(_13150_), .B(_13250_), .Y(_00300_));
NAND_g _19772_ (.A(_08836_), .B(_10604_), .Y(_13251_));
NAND_g _19773_ (.A(cpuregs[25][26]), .B(_09027_), .Y(_13252_));
NAND_g _19774_ (.A(cpuregs[29][26]), .B(_00007_[2]), .Y(_13253_));
AND_g _19775_ (.A(_00007_[0]), .B(_13253_), .Y(_13254_));
NAND_g _19776_ (.A(_13252_), .B(_13254_), .Y(_13255_));
NAND_g _19777_ (.A(cpuregs[24][26]), .B(_09027_), .Y(_13256_));
NAND_g _19778_ (.A(cpuregs[28][26]), .B(_00007_[2]), .Y(_13257_));
AND_g _19779_ (.A(_09025_), .B(_13257_), .Y(_13258_));
NAND_g _19780_ (.A(_13256_), .B(_13258_), .Y(_13259_));
AND_g _19781_ (.A(_00007_[3]), .B(_13259_), .Y(_13260_));
NAND_g _19782_ (.A(_13255_), .B(_13260_), .Y(_13261_));
NAND_g _19783_ (.A(cpuregs[21][26]), .B(_00007_[2]), .Y(_13262_));
NAND_g _19784_ (.A(cpuregs[17][26]), .B(_09027_), .Y(_13263_));
AND_g _19785_ (.A(_00007_[0]), .B(_13263_), .Y(_13264_));
NAND_g _19786_ (.A(_13262_), .B(_13264_), .Y(_13265_));
NAND_g _19787_ (.A(cpuregs[20][26]), .B(_00007_[2]), .Y(_13266_));
NAND_g _19788_ (.A(cpuregs[16][26]), .B(_09027_), .Y(_13267_));
AND_g _19789_ (.A(_09025_), .B(_13267_), .Y(_13268_));
NAND_g _19790_ (.A(_13266_), .B(_13268_), .Y(_13269_));
AND_g _19791_ (.A(_09028_), .B(_13269_), .Y(_13270_));
NAND_g _19792_ (.A(_13265_), .B(_13270_), .Y(_13271_));
AND_g _19793_ (.A(_09026_), .B(_13271_), .Y(_13272_));
NAND_g _19794_ (.A(_13261_), .B(_13272_), .Y(_13273_));
NAND_g _19795_ (.A(cpuregs[27][26]), .B(_09027_), .Y(_13274_));
NAND_g _19796_ (.A(cpuregs[31][26]), .B(_00007_[2]), .Y(_13275_));
AND_g _19797_ (.A(_00007_[0]), .B(_13275_), .Y(_13276_));
NAND_g _19798_ (.A(_13274_), .B(_13276_), .Y(_13277_));
NAND_g _19799_ (.A(cpuregs[26][26]), .B(_09027_), .Y(_13278_));
NAND_g _19800_ (.A(cpuregs[30][26]), .B(_00007_[2]), .Y(_13279_));
AND_g _19801_ (.A(_09025_), .B(_13279_), .Y(_13280_));
NAND_g _19802_ (.A(_13278_), .B(_13280_), .Y(_13281_));
AND_g _19803_ (.A(_00007_[3]), .B(_13281_), .Y(_13282_));
NAND_g _19804_ (.A(_13277_), .B(_13282_), .Y(_13283_));
NAND_g _19805_ (.A(cpuregs[19][26]), .B(_09027_), .Y(_13284_));
NAND_g _19806_ (.A(cpuregs[23][26]), .B(_00007_[2]), .Y(_13285_));
AND_g _19807_ (.A(_00007_[0]), .B(_13285_), .Y(_13286_));
NAND_g _19808_ (.A(_13284_), .B(_13286_), .Y(_13287_));
NAND_g _19809_ (.A(cpuregs[18][26]), .B(_09027_), .Y(_13288_));
NAND_g _19810_ (.A(cpuregs[22][26]), .B(_00007_[2]), .Y(_13289_));
AND_g _19811_ (.A(_09025_), .B(_13289_), .Y(_13290_));
NAND_g _19812_ (.A(_13288_), .B(_13290_), .Y(_13291_));
AND_g _19813_ (.A(_09028_), .B(_13291_), .Y(_13292_));
NAND_g _19814_ (.A(_13287_), .B(_13292_), .Y(_13293_));
AND_g _19815_ (.A(_00007_[1]), .B(_13293_), .Y(_13294_));
NAND_g _19816_ (.A(_13283_), .B(_13294_), .Y(_13295_));
NAND_g _19817_ (.A(_13273_), .B(_13295_), .Y(_13296_));
NAND_g _19818_ (.A(_00007_[4]), .B(_13296_), .Y(_13297_));
NOR_g _19819_ (.A(cpuregs[12][26]), .B(_09027_), .Y(_13298_));
NOR_g _19820_ (.A(cpuregs[8][26]), .B(_00007_[2]), .Y(_13299_));
NOR_g _19821_ (.A(_13298_), .B(_13299_), .Y(_13300_));
NOR_g _19822_ (.A(cpuregs[9][26]), .B(_00007_[2]), .Y(_13301_));
NAND_g _19823_ (.A(_08934_), .B(_00007_[2]), .Y(_13302_));
NAND_g _19824_ (.A(cpuregs[4][26]), .B(_00007_[2]), .Y(_13303_));
NAND_g _19825_ (.A(cpuregs[0][26]), .B(_09027_), .Y(_13304_));
AND_g _19826_ (.A(_09025_), .B(_13304_), .Y(_13305_));
NAND_g _19827_ (.A(_13303_), .B(_13305_), .Y(_13306_));
NAND_g _19828_ (.A(cpuregs[1][26]), .B(_09027_), .Y(_13307_));
NAND_g _19829_ (.A(cpuregs[5][26]), .B(_00007_[2]), .Y(_13308_));
AND_g _19830_ (.A(_00007_[0]), .B(_13308_), .Y(_13309_));
NAND_g _19831_ (.A(_13307_), .B(_13309_), .Y(_13310_));
NAND_g _19832_ (.A(cpuregs[3][26]), .B(_09027_), .Y(_13311_));
NAND_g _19833_ (.A(cpuregs[7][26]), .B(_00007_[2]), .Y(_13312_));
AND_g _19834_ (.A(_00007_[0]), .B(_13312_), .Y(_13313_));
NAND_g _19835_ (.A(_13311_), .B(_13313_), .Y(_13314_));
NAND_g _19836_ (.A(cpuregs[2][26]), .B(_09027_), .Y(_13315_));
NAND_g _19837_ (.A(cpuregs[6][26]), .B(_00007_[2]), .Y(_13316_));
AND_g _19838_ (.A(_09025_), .B(_13316_), .Y(_13317_));
NAND_g _19839_ (.A(_13315_), .B(_13317_), .Y(_13318_));
AND_g _19840_ (.A(_09028_), .B(_13314_), .Y(_13319_));
NAND_g _19841_ (.A(_13318_), .B(_13319_), .Y(_13320_));
NAND_g _19842_ (.A(cpuregs[15][26]), .B(_00007_[2]), .Y(_13321_));
NAND_g _19843_ (.A(cpuregs[11][26]), .B(_09027_), .Y(_13322_));
AND_g _19844_ (.A(_00007_[0]), .B(_13322_), .Y(_13323_));
NAND_g _19845_ (.A(_13321_), .B(_13323_), .Y(_13324_));
NAND_g _19846_ (.A(cpuregs[10][26]), .B(_09027_), .Y(_13325_));
NAND_g _19847_ (.A(cpuregs[14][26]), .B(_00007_[2]), .Y(_13326_));
AND_g _19848_ (.A(_09025_), .B(_13326_), .Y(_13327_));
NAND_g _19849_ (.A(_13325_), .B(_13327_), .Y(_13328_));
AND_g _19850_ (.A(_00007_[3]), .B(_13328_), .Y(_13329_));
NAND_g _19851_ (.A(_13324_), .B(_13329_), .Y(_13330_));
NAND_g _19852_ (.A(_13306_), .B(_13310_), .Y(_13331_));
NAND_g _19853_ (.A(_09028_), .B(_13331_), .Y(_13332_));
NAND_g _19854_ (.A(_09025_), .B(_13300_), .Y(_13333_));
NOR_g _19855_ (.A(_09025_), .B(_13301_), .Y(_13334_));
NAND_g _19856_ (.A(_13302_), .B(_13334_), .Y(_13335_));
AND_g _19857_ (.A(_00007_[3]), .B(_13335_), .Y(_13336_));
NAND_g _19858_ (.A(_13333_), .B(_13336_), .Y(_13337_));
AND_g _19859_ (.A(_13332_), .B(_13337_), .Y(_13338_));
NAND_g _19860_ (.A(_09026_), .B(_13338_), .Y(_13339_));
NAND_g _19861_ (.A(_13320_), .B(_13330_), .Y(_13340_));
NAND_g _19862_ (.A(_00007_[1]), .B(_13340_), .Y(_13341_));
AND_g _19863_ (.A(_09029_), .B(_13341_), .Y(_13342_));
NAND_g _19864_ (.A(_13339_), .B(_13342_), .Y(_13343_));
AND_g _19865_ (.A(_13297_), .B(_13343_), .Y(_13344_));
NAND_g _19866_ (.A(_11170_), .B(_13344_), .Y(_13345_));
NAND_g _19867_ (.A(decoded_imm[26]), .B(_10606_), .Y(_13346_));
AND_g _19868_ (.A(_10603_), .B(_13346_), .Y(_13347_));
NAND_g _19869_ (.A(_13345_), .B(_13347_), .Y(_13348_));
AND_g _19870_ (.A(_13251_), .B(_13348_), .Y(_00301_));
NAND_g _19871_ (.A(_08837_), .B(_10604_), .Y(_13349_));
NAND_g _19872_ (.A(cpuregs[9][27]), .B(_09027_), .Y(_13350_));
NAND_g _19873_ (.A(cpuregs[13][27]), .B(_00007_[2]), .Y(_13351_));
NAND_g _19874_ (.A(_13350_), .B(_13351_), .Y(_13352_));
NAND_g _19875_ (.A(_00007_[0]), .B(_13352_), .Y(_13353_));
NAND_g _19876_ (.A(cpuregs[12][27]), .B(_00007_[2]), .Y(_13354_));
NAND_g _19877_ (.A(cpuregs[8][27]), .B(_09027_), .Y(_13355_));
NAND_g _19878_ (.A(_13354_), .B(_13355_), .Y(_13356_));
NAND_g _19879_ (.A(_09025_), .B(_13356_), .Y(_13357_));
NAND_g _19880_ (.A(_13353_), .B(_13357_), .Y(_13358_));
NAND_g _19881_ (.A(_09026_), .B(_13358_), .Y(_13359_));
NAND_g _19882_ (.A(cpuregs[11][27]), .B(_09027_), .Y(_13360_));
NAND_g _19883_ (.A(cpuregs[15][27]), .B(_00007_[2]), .Y(_13361_));
NAND_g _19884_ (.A(_13360_), .B(_13361_), .Y(_13362_));
NAND_g _19885_ (.A(_00007_[0]), .B(_13362_), .Y(_13363_));
NAND_g _19886_ (.A(cpuregs[14][27]), .B(_00007_[2]), .Y(_13364_));
NAND_g _19887_ (.A(cpuregs[10][27]), .B(_09027_), .Y(_13365_));
NAND_g _19888_ (.A(_13364_), .B(_13365_), .Y(_13366_));
NAND_g _19889_ (.A(_09025_), .B(_13366_), .Y(_13367_));
NAND_g _19890_ (.A(_13363_), .B(_13367_), .Y(_13368_));
NAND_g _19891_ (.A(_00007_[1]), .B(_13368_), .Y(_13369_));
NAND_g _19892_ (.A(cpuregs[31][27]), .B(_00007_[2]), .Y(_13370_));
NAND_g _19893_ (.A(cpuregs[27][27]), .B(_09027_), .Y(_13371_));
AND_g _19894_ (.A(_00007_[0]), .B(_13371_), .Y(_13372_));
NAND_g _19895_ (.A(_13370_), .B(_13372_), .Y(_13373_));
NAND_g _19896_ (.A(cpuregs[26][27]), .B(_09027_), .Y(_13374_));
NAND_g _19897_ (.A(cpuregs[30][27]), .B(_00007_[2]), .Y(_13375_));
AND_g _19898_ (.A(_09025_), .B(_13375_), .Y(_13376_));
NAND_g _19899_ (.A(_13374_), .B(_13376_), .Y(_13377_));
AND_g _19900_ (.A(_00007_[1]), .B(_13377_), .Y(_13378_));
NAND_g _19901_ (.A(_13373_), .B(_13378_), .Y(_13379_));
NAND_g _19902_ (.A(cpuregs[29][27]), .B(_00007_[2]), .Y(_13380_));
NAND_g _19903_ (.A(cpuregs[25][27]), .B(_09027_), .Y(_13381_));
AND_g _19904_ (.A(_00007_[0]), .B(_13381_), .Y(_13382_));
NAND_g _19905_ (.A(_13380_), .B(_13382_), .Y(_13383_));
NAND_g _19906_ (.A(cpuregs[24][27]), .B(_09027_), .Y(_13384_));
NAND_g _19907_ (.A(cpuregs[28][27]), .B(_00007_[2]), .Y(_13385_));
AND_g _19908_ (.A(_09025_), .B(_13385_), .Y(_13386_));
NAND_g _19909_ (.A(_13384_), .B(_13386_), .Y(_13387_));
AND_g _19910_ (.A(_09026_), .B(_13387_), .Y(_13388_));
NAND_g _19911_ (.A(_13383_), .B(_13388_), .Y(_13389_));
NAND_g _19912_ (.A(cpuregs[1][27]), .B(_09027_), .Y(_13390_));
NAND_g _19913_ (.A(cpuregs[5][27]), .B(_00007_[2]), .Y(_13391_));
NAND_g _19914_ (.A(_13390_), .B(_13391_), .Y(_13392_));
NAND_g _19915_ (.A(_00007_[0]), .B(_13392_), .Y(_13393_));
NAND_g _19916_ (.A(cpuregs[4][27]), .B(_00007_[2]), .Y(_13394_));
NAND_g _19917_ (.A(cpuregs[0][27]), .B(_09027_), .Y(_13395_));
NAND_g _19918_ (.A(_13394_), .B(_13395_), .Y(_13396_));
NAND_g _19919_ (.A(_09025_), .B(_13396_), .Y(_13397_));
NAND_g _19920_ (.A(_13393_), .B(_13397_), .Y(_13398_));
NAND_g _19921_ (.A(_09026_), .B(_13398_), .Y(_13399_));
NAND_g _19922_ (.A(cpuregs[6][27]), .B(_00007_[2]), .Y(_13400_));
NAND_g _19923_ (.A(cpuregs[2][27]), .B(_09027_), .Y(_13401_));
NAND_g _19924_ (.A(_13400_), .B(_13401_), .Y(_13402_));
NAND_g _19925_ (.A(_09025_), .B(_13402_), .Y(_13403_));
NOR_g _19926_ (.A(cpuregs[3][27]), .B(_00007_[2]), .Y(_13404_));
NAND_g _19927_ (.A(_08978_), .B(_00007_[2]), .Y(_13405_));
NOR_g _19928_ (.A(_09025_), .B(_13404_), .Y(_13406_));
NAND_g _19929_ (.A(_13405_), .B(_13406_), .Y(_13407_));
NAND_g _19930_ (.A(_13403_), .B(_13407_), .Y(_13408_));
NAND_g _19931_ (.A(_00007_[1]), .B(_13408_), .Y(_13409_));
NAND_g _19932_ (.A(_08938_), .B(_09027_), .Y(_13410_));
NOR_g _19933_ (.A(cpuregs[22][27]), .B(_09027_), .Y(_13411_));
NAND_g _19934_ (.A(_08901_), .B(_00007_[2]), .Y(_13412_));
NOR_g _19935_ (.A(cpuregs[19][27]), .B(_00007_[2]), .Y(_13413_));
NOR_g _19936_ (.A(_00007_[0]), .B(_13411_), .Y(_13414_));
AND_g _19937_ (.A(_13410_), .B(_13414_), .Y(_13415_));
NAND_g _19938_ (.A(_00007_[0]), .B(_13412_), .Y(_13416_));
NOR_g _19939_ (.A(_13413_), .B(_13416_), .Y(_13417_));
NOR_g _19940_ (.A(_13415_), .B(_13417_), .Y(_13418_));
NOR_g _19941_ (.A(cpuregs[16][27]), .B(_00007_[2]), .Y(_13419_));
NOR_g _19942_ (.A(cpuregs[20][27]), .B(_09027_), .Y(_13420_));
NOR_g _19943_ (.A(_13419_), .B(_13420_), .Y(_13421_));
NOR_g _19944_ (.A(cpuregs[17][27]), .B(_00007_[2]), .Y(_13422_));
NAND_g _19945_ (.A(_09000_), .B(_00007_[2]), .Y(_13423_));
NAND_g _19946_ (.A(_00007_[0]), .B(_13423_), .Y(_13424_));
NOR_g _19947_ (.A(_13422_), .B(_13424_), .Y(_13425_));
AND_g _19948_ (.A(_09025_), .B(_13421_), .Y(_13426_));
NOR_g _19949_ (.A(_13425_), .B(_13426_), .Y(_13427_));
NAND_g _19950_ (.A(_00007_[1]), .B(_13418_), .Y(_13428_));
NAND_g _19951_ (.A(_09026_), .B(_13427_), .Y(_13429_));
AND_g _19952_ (.A(_09028_), .B(_13429_), .Y(_13430_));
NAND_g _19953_ (.A(_13428_), .B(_13430_), .Y(_13431_));
NAND_g _19954_ (.A(_13379_), .B(_13389_), .Y(_13432_));
NAND_g _19955_ (.A(_00007_[3]), .B(_13432_), .Y(_13433_));
AND_g _19956_ (.A(_00007_[4]), .B(_13433_), .Y(_13434_));
NAND_g _19957_ (.A(_13431_), .B(_13434_), .Y(_13435_));
NAND_g _19958_ (.A(_13359_), .B(_13369_), .Y(_13436_));
NAND_g _19959_ (.A(_00007_[3]), .B(_13436_), .Y(_13437_));
NAND_g _19960_ (.A(_13399_), .B(_13409_), .Y(_13438_));
NAND_g _19961_ (.A(_09028_), .B(_13438_), .Y(_13439_));
AND_g _19962_ (.A(_13437_), .B(_13439_), .Y(_13440_));
NAND_g _19963_ (.A(_09029_), .B(_13440_), .Y(_13441_));
AND_g _19964_ (.A(_13435_), .B(_13441_), .Y(_13442_));
NAND_g _19965_ (.A(_11170_), .B(_13442_), .Y(_13443_));
NAND_g _19966_ (.A(decoded_imm[27]), .B(_10606_), .Y(_13444_));
AND_g _19967_ (.A(_10603_), .B(_13444_), .Y(_13445_));
NAND_g _19968_ (.A(_13443_), .B(_13445_), .Y(_13446_));
AND_g _19969_ (.A(_13349_), .B(_13446_), .Y(_00302_));
NAND_g _19970_ (.A(_08838_), .B(_10604_), .Y(_13447_));
NAND_g _19971_ (.A(cpuregs[18][28]), .B(_00007_[1]), .Y(_13448_));
NAND_g _19972_ (.A(cpuregs[16][28]), .B(_09026_), .Y(_13449_));
NAND_g _19973_ (.A(_13448_), .B(_13449_), .Y(_13450_));
NAND_g _19974_ (.A(_09027_), .B(_13450_), .Y(_13451_));
NAND_g _19975_ (.A(cpuregs[22][28]), .B(_00007_[1]), .Y(_13452_));
NAND_g _19976_ (.A(cpuregs[20][28]), .B(_09026_), .Y(_13453_));
NAND_g _19977_ (.A(_13452_), .B(_13453_), .Y(_13454_));
NAND_g _19978_ (.A(_00007_[2]), .B(_13454_), .Y(_13455_));
AND_g _19979_ (.A(_09025_), .B(_13455_), .Y(_13456_));
NAND_g _19980_ (.A(_13451_), .B(_13456_), .Y(_13457_));
NAND_g _19981_ (.A(cpuregs[19][28]), .B(_00007_[1]), .Y(_13458_));
NAND_g _19982_ (.A(cpuregs[17][28]), .B(_09026_), .Y(_13459_));
NAND_g _19983_ (.A(_13458_), .B(_13459_), .Y(_13460_));
NAND_g _19984_ (.A(_09027_), .B(_13460_), .Y(_13461_));
NAND_g _19985_ (.A(cpuregs[23][28]), .B(_00007_[1]), .Y(_13462_));
NAND_g _19986_ (.A(cpuregs[21][28]), .B(_09026_), .Y(_13463_));
NAND_g _19987_ (.A(_13462_), .B(_13463_), .Y(_13464_));
NAND_g _19988_ (.A(_00007_[2]), .B(_13464_), .Y(_13465_));
AND_g _19989_ (.A(_00007_[0]), .B(_13465_), .Y(_13466_));
NAND_g _19990_ (.A(_13461_), .B(_13466_), .Y(_13467_));
AND_g _19991_ (.A(_13457_), .B(_13467_), .Y(_13468_));
NAND_g _19992_ (.A(cpuregs[26][28]), .B(_09027_), .Y(_13469_));
NAND_g _19993_ (.A(cpuregs[30][28]), .B(_00007_[2]), .Y(_13470_));
AND_g _19994_ (.A(_09025_), .B(_13470_), .Y(_13471_));
NAND_g _19995_ (.A(_13469_), .B(_13471_), .Y(_13472_));
NAND_g _19996_ (.A(cpuregs[31][28]), .B(_00007_[2]), .Y(_13473_));
NAND_g _19997_ (.A(cpuregs[27][28]), .B(_09027_), .Y(_13474_));
AND_g _19998_ (.A(_00007_[0]), .B(_13474_), .Y(_13475_));
NAND_g _19999_ (.A(_13473_), .B(_13475_), .Y(_13476_));
NAND_g _20000_ (.A(_13472_), .B(_13476_), .Y(_13477_));
NAND_g _20001_ (.A(_00007_[1]), .B(_13477_), .Y(_13478_));
NAND_g _20002_ (.A(cpuregs[24][28]), .B(_09027_), .Y(_13479_));
NAND_g _20003_ (.A(cpuregs[28][28]), .B(_00007_[2]), .Y(_13480_));
AND_g _20004_ (.A(_09025_), .B(_13480_), .Y(_13481_));
NAND_g _20005_ (.A(_13479_), .B(_13481_), .Y(_13482_));
NAND_g _20006_ (.A(cpuregs[25][28]), .B(_09027_), .Y(_13483_));
NAND_g _20007_ (.A(cpuregs[29][28]), .B(_00007_[2]), .Y(_13484_));
AND_g _20008_ (.A(_00007_[0]), .B(_13484_), .Y(_13485_));
NAND_g _20009_ (.A(_13483_), .B(_13485_), .Y(_13486_));
NAND_g _20010_ (.A(_13482_), .B(_13486_), .Y(_13487_));
NAND_g _20011_ (.A(_09026_), .B(_13487_), .Y(_13488_));
AND_g _20012_ (.A(_00007_[3]), .B(_13488_), .Y(_13489_));
NAND_g _20013_ (.A(_13478_), .B(_13489_), .Y(_13490_));
NAND_g _20014_ (.A(_09028_), .B(_13468_), .Y(_13491_));
AND_g _20015_ (.A(_00007_[4]), .B(_13490_), .Y(_13492_));
AND_g _20016_ (.A(_13491_), .B(_13492_), .Y(_13493_));
NAND_g _20017_ (.A(_08979_), .B(_00007_[2]), .Y(_13494_));
NOR_g _20018_ (.A(cpuregs[3][28]), .B(_00007_[2]), .Y(_13495_));
NOR_g _20019_ (.A(cpuregs[2][28]), .B(_00007_[2]), .Y(_13496_));
AND_g _20020_ (.A(_09016_), .B(_00007_[2]), .Y(_13497_));
NOR_g _20021_ (.A(_13496_), .B(_13497_), .Y(_13498_));
NOR_g _20022_ (.A(_09025_), .B(_13495_), .Y(_13499_));
NAND_g _20023_ (.A(_13494_), .B(_13499_), .Y(_13500_));
NAND_g _20024_ (.A(_09025_), .B(_13498_), .Y(_13501_));
AND_g _20025_ (.A(_13500_), .B(_13501_), .Y(_13502_));
NAND_g _20026_ (.A(_00007_[1]), .B(_13502_), .Y(_13503_));
NOR_g _20027_ (.A(cpuregs[1][28]), .B(_00007_[2]), .Y(_13504_));
NAND_g _20028_ (.A(_08960_), .B(_00007_[2]), .Y(_13505_));
NOR_g _20029_ (.A(cpuregs[0][28]), .B(_00007_[2]), .Y(_13506_));
AND_g _20030_ (.A(_08917_), .B(_00007_[2]), .Y(_13507_));
NOR_g _20031_ (.A(_13506_), .B(_13507_), .Y(_13508_));
NOR_g _20032_ (.A(_09025_), .B(_13504_), .Y(_13509_));
NAND_g _20033_ (.A(_13505_), .B(_13509_), .Y(_13510_));
NAND_g _20034_ (.A(_09025_), .B(_13508_), .Y(_13511_));
AND_g _20035_ (.A(_13510_), .B(_13511_), .Y(_13512_));
NAND_g _20036_ (.A(_09026_), .B(_13512_), .Y(_13513_));
NAND_g _20037_ (.A(_13503_), .B(_13513_), .Y(_13514_));
NAND_g _20038_ (.A(_09028_), .B(_13514_), .Y(_13515_));
NAND_g _20039_ (.A(cpuregs[9][28]), .B(_09026_), .Y(_13516_));
NAND_g _20040_ (.A(cpuregs[11][28]), .B(_00007_[1]), .Y(_13517_));
AND_g _20041_ (.A(_09027_), .B(_13517_), .Y(_13518_));
NAND_g _20042_ (.A(_13516_), .B(_13518_), .Y(_13519_));
NAND_g _20043_ (.A(cpuregs[13][28]), .B(_09026_), .Y(_13520_));
NAND_g _20044_ (.A(cpuregs[15][28]), .B(_00007_[1]), .Y(_13521_));
AND_g _20045_ (.A(_00007_[2]), .B(_13521_), .Y(_13522_));
NAND_g _20046_ (.A(_13520_), .B(_13522_), .Y(_13523_));
NAND_g _20047_ (.A(_13519_), .B(_13523_), .Y(_13524_));
NAND_g _20048_ (.A(_00007_[0]), .B(_13524_), .Y(_13525_));
NAND_g _20049_ (.A(cpuregs[8][28]), .B(_09026_), .Y(_13526_));
NAND_g _20050_ (.A(cpuregs[10][28]), .B(_00007_[1]), .Y(_13527_));
AND_g _20051_ (.A(_09027_), .B(_13527_), .Y(_13528_));
NAND_g _20052_ (.A(_13526_), .B(_13528_), .Y(_13529_));
NAND_g _20053_ (.A(cpuregs[12][28]), .B(_09026_), .Y(_13530_));
NAND_g _20054_ (.A(cpuregs[14][28]), .B(_00007_[1]), .Y(_13531_));
AND_g _20055_ (.A(_00007_[2]), .B(_13531_), .Y(_13532_));
NAND_g _20056_ (.A(_13530_), .B(_13532_), .Y(_13533_));
NAND_g _20057_ (.A(_13529_), .B(_13533_), .Y(_13534_));
NAND_g _20058_ (.A(_09025_), .B(_13534_), .Y(_13535_));
NAND_g _20059_ (.A(_13525_), .B(_13535_), .Y(_13536_));
NAND_g _20060_ (.A(_00007_[3]), .B(_13536_), .Y(_13537_));
NAND_g _20061_ (.A(_13515_), .B(_13537_), .Y(_13538_));
AND_g _20062_ (.A(_09029_), .B(_13538_), .Y(_13539_));
NOR_g _20063_ (.A(_13493_), .B(_13539_), .Y(_13540_));
NAND_g _20064_ (.A(_11170_), .B(_13540_), .Y(_13541_));
NAND_g _20065_ (.A(decoded_imm[28]), .B(_10606_), .Y(_13542_));
AND_g _20066_ (.A(_10603_), .B(_13542_), .Y(_13543_));
NAND_g _20067_ (.A(_13541_), .B(_13543_), .Y(_13544_));
AND_g _20068_ (.A(_13447_), .B(_13544_), .Y(_00303_));
NAND_g _20069_ (.A(_08839_), .B(_10604_), .Y(_13545_));
NAND_g _20070_ (.A(cpuregs[13][29]), .B(_00007_[2]), .Y(_13546_));
NAND_g _20071_ (.A(cpuregs[9][29]), .B(_09027_), .Y(_13547_));
AND_g _20072_ (.A(_00007_[0]), .B(_13547_), .Y(_13548_));
NAND_g _20073_ (.A(_13546_), .B(_13548_), .Y(_13549_));
NAND_g _20074_ (.A(cpuregs[8][29]), .B(_09027_), .Y(_13550_));
NAND_g _20075_ (.A(cpuregs[12][29]), .B(_00007_[2]), .Y(_13551_));
AND_g _20076_ (.A(_09025_), .B(_13551_), .Y(_13552_));
NAND_g _20077_ (.A(_13550_), .B(_13552_), .Y(_13553_));
AND_g _20078_ (.A(_00007_[3]), .B(_13553_), .Y(_13554_));
NAND_g _20079_ (.A(_13549_), .B(_13554_), .Y(_13555_));
NAND_g _20080_ (.A(cpuregs[1][29]), .B(_09027_), .Y(_13556_));
NAND_g _20081_ (.A(cpuregs[5][29]), .B(_00007_[2]), .Y(_13557_));
AND_g _20082_ (.A(_00007_[0]), .B(_13557_), .Y(_13558_));
NAND_g _20083_ (.A(_13556_), .B(_13558_), .Y(_13559_));
NAND_g _20084_ (.A(cpuregs[0][29]), .B(_09027_), .Y(_13560_));
NAND_g _20085_ (.A(cpuregs[4][29]), .B(_00007_[2]), .Y(_13561_));
AND_g _20086_ (.A(_09025_), .B(_13561_), .Y(_13562_));
NAND_g _20087_ (.A(_13560_), .B(_13562_), .Y(_13563_));
AND_g _20088_ (.A(_09028_), .B(_13559_), .Y(_13564_));
NAND_g _20089_ (.A(_13563_), .B(_13564_), .Y(_13565_));
NAND_g _20090_ (.A(cpuregs[3][29]), .B(_09027_), .Y(_13566_));
NAND_g _20091_ (.A(cpuregs[7][29]), .B(_00007_[2]), .Y(_13567_));
AND_g _20092_ (.A(_00007_[0]), .B(_13567_), .Y(_13568_));
NAND_g _20093_ (.A(_13566_), .B(_13568_), .Y(_13569_));
NAND_g _20094_ (.A(cpuregs[2][29]), .B(_09027_), .Y(_13570_));
NAND_g _20095_ (.A(cpuregs[6][29]), .B(_00007_[2]), .Y(_13571_));
AND_g _20096_ (.A(_09025_), .B(_13571_), .Y(_13572_));
NAND_g _20097_ (.A(_13570_), .B(_13572_), .Y(_13573_));
AND_g _20098_ (.A(_09028_), .B(_13569_), .Y(_13574_));
NAND_g _20099_ (.A(_13573_), .B(_13574_), .Y(_13575_));
NAND_g _20100_ (.A(cpuregs[15][29]), .B(_00007_[2]), .Y(_13576_));
NAND_g _20101_ (.A(cpuregs[11][29]), .B(_09027_), .Y(_13577_));
AND_g _20102_ (.A(_00007_[0]), .B(_13577_), .Y(_13578_));
NAND_g _20103_ (.A(_13576_), .B(_13578_), .Y(_13579_));
NAND_g _20104_ (.A(cpuregs[10][29]), .B(_09027_), .Y(_13580_));
NAND_g _20105_ (.A(cpuregs[14][29]), .B(_00007_[2]), .Y(_13581_));
AND_g _20106_ (.A(_09025_), .B(_13581_), .Y(_13582_));
NAND_g _20107_ (.A(_13580_), .B(_13582_), .Y(_13583_));
AND_g _20108_ (.A(_00007_[3]), .B(_13583_), .Y(_13584_));
NAND_g _20109_ (.A(_13579_), .B(_13584_), .Y(_13585_));
NAND_g _20110_ (.A(_13575_), .B(_13585_), .Y(_13586_));
NAND_g _20111_ (.A(_00007_[1]), .B(_13586_), .Y(_13587_));
NAND_g _20112_ (.A(_13555_), .B(_13565_), .Y(_13588_));
NAND_g _20113_ (.A(_09026_), .B(_13588_), .Y(_13589_));
AND_g _20114_ (.A(_13587_), .B(_13589_), .Y(_13590_));
NAND_g _20115_ (.A(_09029_), .B(_13590_), .Y(_13591_));
NAND_g _20116_ (.A(cpuregs[25][29]), .B(_09027_), .Y(_13592_));
NAND_g _20117_ (.A(cpuregs[29][29]), .B(_00007_[2]), .Y(_13593_));
AND_g _20118_ (.A(_00007_[0]), .B(_13593_), .Y(_13594_));
NAND_g _20119_ (.A(_13592_), .B(_13594_), .Y(_13595_));
NAND_g _20120_ (.A(cpuregs[24][29]), .B(_09027_), .Y(_13596_));
NAND_g _20121_ (.A(cpuregs[28][29]), .B(_00007_[2]), .Y(_13597_));
AND_g _20122_ (.A(_09025_), .B(_13597_), .Y(_13598_));
NAND_g _20123_ (.A(_13596_), .B(_13598_), .Y(_13599_));
AND_g _20124_ (.A(_00007_[3]), .B(_13599_), .Y(_13600_));
NAND_g _20125_ (.A(_13595_), .B(_13600_), .Y(_13601_));
NAND_g _20126_ (.A(cpuregs[21][29]), .B(_00007_[2]), .Y(_13602_));
NAND_g _20127_ (.A(cpuregs[17][29]), .B(_09027_), .Y(_13603_));
AND_g _20128_ (.A(_00007_[0]), .B(_13603_), .Y(_13604_));
NAND_g _20129_ (.A(_13602_), .B(_13604_), .Y(_13605_));
NAND_g _20130_ (.A(cpuregs[20][29]), .B(_00007_[2]), .Y(_13606_));
NAND_g _20131_ (.A(cpuregs[16][29]), .B(_09027_), .Y(_13607_));
AND_g _20132_ (.A(_09025_), .B(_13607_), .Y(_13608_));
NAND_g _20133_ (.A(_13606_), .B(_13608_), .Y(_13609_));
AND_g _20134_ (.A(_09028_), .B(_13609_), .Y(_13610_));
NAND_g _20135_ (.A(_13605_), .B(_13610_), .Y(_13611_));
AND_g _20136_ (.A(_09026_), .B(_13611_), .Y(_13612_));
NAND_g _20137_ (.A(_13601_), .B(_13612_), .Y(_13613_));
NAND_g _20138_ (.A(cpuregs[27][29]), .B(_09027_), .Y(_13614_));
NAND_g _20139_ (.A(cpuregs[31][29]), .B(_00007_[2]), .Y(_13615_));
AND_g _20140_ (.A(_00007_[0]), .B(_13615_), .Y(_13616_));
NAND_g _20141_ (.A(_13614_), .B(_13616_), .Y(_13617_));
NAND_g _20142_ (.A(cpuregs[26][29]), .B(_09027_), .Y(_13618_));
NAND_g _20143_ (.A(cpuregs[30][29]), .B(_00007_[2]), .Y(_13619_));
AND_g _20144_ (.A(_09025_), .B(_13619_), .Y(_13620_));
NAND_g _20145_ (.A(_13618_), .B(_13620_), .Y(_13621_));
AND_g _20146_ (.A(_00007_[3]), .B(_13621_), .Y(_13622_));
NAND_g _20147_ (.A(_13617_), .B(_13622_), .Y(_13623_));
NAND_g _20148_ (.A(cpuregs[19][29]), .B(_09027_), .Y(_13624_));
NAND_g _20149_ (.A(cpuregs[23][29]), .B(_00007_[2]), .Y(_13625_));
AND_g _20150_ (.A(_00007_[0]), .B(_13625_), .Y(_13626_));
NAND_g _20151_ (.A(_13624_), .B(_13626_), .Y(_13627_));
NAND_g _20152_ (.A(cpuregs[18][29]), .B(_09027_), .Y(_13628_));
NAND_g _20153_ (.A(cpuregs[22][29]), .B(_00007_[2]), .Y(_13629_));
AND_g _20154_ (.A(_09025_), .B(_13629_), .Y(_13630_));
NAND_g _20155_ (.A(_13628_), .B(_13630_), .Y(_13631_));
AND_g _20156_ (.A(_09028_), .B(_13631_), .Y(_13632_));
NAND_g _20157_ (.A(_13627_), .B(_13632_), .Y(_13633_));
AND_g _20158_ (.A(_00007_[1]), .B(_13633_), .Y(_13634_));
NAND_g _20159_ (.A(_13623_), .B(_13634_), .Y(_13635_));
NAND_g _20160_ (.A(_13613_), .B(_13635_), .Y(_13636_));
NAND_g _20161_ (.A(_00007_[4]), .B(_13636_), .Y(_13637_));
AND_g _20162_ (.A(_13591_), .B(_13637_), .Y(_13638_));
NAND_g _20163_ (.A(_11170_), .B(_13638_), .Y(_13639_));
NAND_g _20164_ (.A(decoded_imm[29]), .B(_10606_), .Y(_13640_));
AND_g _20165_ (.A(_10603_), .B(_13640_), .Y(_13641_));
NAND_g _20166_ (.A(_13639_), .B(_13641_), .Y(_13642_));
AND_g _20167_ (.A(_13545_), .B(_13642_), .Y(_00304_));
NAND_g _20168_ (.A(_08840_), .B(_10604_), .Y(_13643_));
NAND_g _20169_ (.A(cpuregs[22][30]), .B(_00007_[1]), .Y(_13644_));
NAND_g _20170_ (.A(cpuregs[20][30]), .B(_09026_), .Y(_13645_));
NAND_g _20171_ (.A(_13644_), .B(_13645_), .Y(_13646_));
NAND_g _20172_ (.A(_00007_[2]), .B(_13646_), .Y(_13647_));
NAND_g _20173_ (.A(cpuregs[18][30]), .B(_00007_[1]), .Y(_13648_));
NAND_g _20174_ (.A(cpuregs[16][30]), .B(_09026_), .Y(_13649_));
NAND_g _20175_ (.A(_13648_), .B(_13649_), .Y(_13650_));
NAND_g _20176_ (.A(_09027_), .B(_13650_), .Y(_13651_));
NAND_g _20177_ (.A(_13647_), .B(_13651_), .Y(_13652_));
AND_g _20178_ (.A(_09025_), .B(_13652_), .Y(_13653_));
NOT_g _20179_ (.A(_13653_), .Y(_13654_));
NAND_g _20180_ (.A(cpuregs[23][30]), .B(_00007_[1]), .Y(_13655_));
NAND_g _20181_ (.A(cpuregs[21][30]), .B(_09026_), .Y(_13656_));
NAND_g _20182_ (.A(_13655_), .B(_13656_), .Y(_13657_));
NAND_g _20183_ (.A(_00007_[2]), .B(_13657_), .Y(_13658_));
NAND_g _20184_ (.A(cpuregs[19][30]), .B(_00007_[1]), .Y(_13659_));
NAND_g _20185_ (.A(cpuregs[17][30]), .B(_09026_), .Y(_13660_));
NAND_g _20186_ (.A(_13659_), .B(_13660_), .Y(_13661_));
NAND_g _20187_ (.A(_09027_), .B(_13661_), .Y(_13662_));
NAND_g _20188_ (.A(_13658_), .B(_13662_), .Y(_13663_));
NAND_g _20189_ (.A(_00007_[0]), .B(_13663_), .Y(_13664_));
AND_g _20190_ (.A(_09028_), .B(_13664_), .Y(_13665_));
NAND_g _20191_ (.A(_13654_), .B(_13665_), .Y(_13666_));
NAND_g _20192_ (.A(cpuregs[31][30]), .B(_00007_[2]), .Y(_13667_));
NAND_g _20193_ (.A(cpuregs[27][30]), .B(_09027_), .Y(_13668_));
AND_g _20194_ (.A(_00007_[0]), .B(_13668_), .Y(_13669_));
NAND_g _20195_ (.A(_13667_), .B(_13669_), .Y(_13670_));
NAND_g _20196_ (.A(cpuregs[26][30]), .B(_09027_), .Y(_13671_));
NAND_g _20197_ (.A(cpuregs[30][30]), .B(_00007_[2]), .Y(_13672_));
AND_g _20198_ (.A(_09025_), .B(_13672_), .Y(_13673_));
NAND_g _20199_ (.A(_13671_), .B(_13673_), .Y(_13674_));
AND_g _20200_ (.A(_00007_[1]), .B(_13674_), .Y(_13675_));
NAND_g _20201_ (.A(_13670_), .B(_13675_), .Y(_13676_));
NAND_g _20202_ (.A(cpuregs[25][30]), .B(_09027_), .Y(_13677_));
NAND_g _20203_ (.A(cpuregs[29][30]), .B(_00007_[2]), .Y(_13678_));
AND_g _20204_ (.A(_00007_[0]), .B(_13678_), .Y(_13679_));
NAND_g _20205_ (.A(_13677_), .B(_13679_), .Y(_13680_));
NAND_g _20206_ (.A(cpuregs[24][30]), .B(_09027_), .Y(_13681_));
NAND_g _20207_ (.A(cpuregs[28][30]), .B(_00007_[2]), .Y(_13682_));
AND_g _20208_ (.A(_09025_), .B(_13682_), .Y(_13683_));
NAND_g _20209_ (.A(_13681_), .B(_13683_), .Y(_13684_));
AND_g _20210_ (.A(_09026_), .B(_13684_), .Y(_13685_));
NAND_g _20211_ (.A(_13680_), .B(_13685_), .Y(_13686_));
AND_g _20212_ (.A(_00007_[3]), .B(_13686_), .Y(_13687_));
NAND_g _20213_ (.A(_13676_), .B(_13687_), .Y(_13688_));
NAND_g _20214_ (.A(_13666_), .B(_13688_), .Y(_13689_));
AND_g _20215_ (.A(_00007_[4]), .B(_13689_), .Y(_13690_));
NAND_g _20216_ (.A(cpuregs[3][30]), .B(_09027_), .Y(_13691_));
NAND_g _20217_ (.A(cpuregs[7][30]), .B(_00007_[2]), .Y(_13692_));
AND_g _20218_ (.A(_00007_[0]), .B(_13692_), .Y(_13693_));
NAND_g _20219_ (.A(_13691_), .B(_13693_), .Y(_13694_));
NAND_g _20220_ (.A(cpuregs[2][30]), .B(_09027_), .Y(_13695_));
NAND_g _20221_ (.A(cpuregs[6][30]), .B(_00007_[2]), .Y(_13696_));
AND_g _20222_ (.A(_09025_), .B(_13696_), .Y(_13697_));
NAND_g _20223_ (.A(_13695_), .B(_13697_), .Y(_13698_));
AND_g _20224_ (.A(_00007_[1]), .B(_13698_), .Y(_13699_));
NAND_g _20225_ (.A(_13694_), .B(_13699_), .Y(_13700_));
NAND_g _20226_ (.A(cpuregs[1][30]), .B(_09027_), .Y(_13701_));
NAND_g _20227_ (.A(cpuregs[5][30]), .B(_00007_[2]), .Y(_13702_));
AND_g _20228_ (.A(_00007_[0]), .B(_13702_), .Y(_13703_));
NAND_g _20229_ (.A(_13701_), .B(_13703_), .Y(_13704_));
NAND_g _20230_ (.A(cpuregs[0][30]), .B(_09027_), .Y(_13705_));
NAND_g _20231_ (.A(cpuregs[4][30]), .B(_00007_[2]), .Y(_13706_));
AND_g _20232_ (.A(_09025_), .B(_13706_), .Y(_13707_));
NAND_g _20233_ (.A(_13705_), .B(_13707_), .Y(_13708_));
AND_g _20234_ (.A(_09026_), .B(_13708_), .Y(_13709_));
NAND_g _20235_ (.A(_13704_), .B(_13709_), .Y(_13710_));
AND_g _20236_ (.A(_09028_), .B(_13710_), .Y(_13711_));
NAND_g _20237_ (.A(_13700_), .B(_13711_), .Y(_13712_));
NAND_g _20238_ (.A(cpuregs[12][30]), .B(_09025_), .Y(_13713_));
NAND_g _20239_ (.A(cpuregs[13][30]), .B(_00007_[0]), .Y(_13714_));
NAND_g _20240_ (.A(_13713_), .B(_13714_), .Y(_13715_));
NAND_g _20241_ (.A(_00007_[2]), .B(_13715_), .Y(_13716_));
NAND_g _20242_ (.A(cpuregs[8][30]), .B(_09025_), .Y(_13717_));
NAND_g _20243_ (.A(cpuregs[9][30]), .B(_00007_[0]), .Y(_13718_));
NAND_g _20244_ (.A(_13717_), .B(_13718_), .Y(_13719_));
NAND_g _20245_ (.A(_09027_), .B(_13719_), .Y(_13720_));
NAND_g _20246_ (.A(_13716_), .B(_13720_), .Y(_13721_));
NAND_g _20247_ (.A(_09026_), .B(_13721_), .Y(_13722_));
NAND_g _20248_ (.A(cpuregs[14][30]), .B(_09025_), .Y(_13723_));
NAND_g _20249_ (.A(cpuregs[15][30]), .B(_00007_[0]), .Y(_13724_));
NAND_g _20250_ (.A(_13723_), .B(_13724_), .Y(_13725_));
NAND_g _20251_ (.A(_00007_[2]), .B(_13725_), .Y(_13726_));
NAND_g _20252_ (.A(cpuregs[10][30]), .B(_09025_), .Y(_13727_));
NAND_g _20253_ (.A(cpuregs[11][30]), .B(_00007_[0]), .Y(_13728_));
NAND_g _20254_ (.A(_13727_), .B(_13728_), .Y(_13729_));
NAND_g _20255_ (.A(_09027_), .B(_13729_), .Y(_13730_));
NAND_g _20256_ (.A(_13726_), .B(_13730_), .Y(_13731_));
NAND_g _20257_ (.A(_00007_[1]), .B(_13731_), .Y(_13732_));
AND_g _20258_ (.A(_00007_[3]), .B(_13732_), .Y(_13733_));
NAND_g _20259_ (.A(_13722_), .B(_13733_), .Y(_13734_));
NAND_g _20260_ (.A(_13712_), .B(_13734_), .Y(_13735_));
AND_g _20261_ (.A(_09029_), .B(_13735_), .Y(_13736_));
NOR_g _20262_ (.A(_13690_), .B(_13736_), .Y(_13737_));
NAND_g _20263_ (.A(_11170_), .B(_13737_), .Y(_13738_));
NAND_g _20264_ (.A(decoded_imm[30]), .B(_10606_), .Y(_13739_));
AND_g _20265_ (.A(_10603_), .B(_13739_), .Y(_13740_));
NAND_g _20266_ (.A(_13738_), .B(_13740_), .Y(_13741_));
AND_g _20267_ (.A(_13643_), .B(_13741_), .Y(_00305_));
NAND_g _20268_ (.A(_08841_), .B(_10604_), .Y(_13742_));
NAND_g _20269_ (.A(cpuregs[25][31]), .B(_09027_), .Y(_13743_));
NAND_g _20270_ (.A(cpuregs[29][31]), .B(_00007_[2]), .Y(_13744_));
AND_g _20271_ (.A(_00007_[0]), .B(_13744_), .Y(_13745_));
NAND_g _20272_ (.A(_13743_), .B(_13745_), .Y(_13746_));
NAND_g _20273_ (.A(cpuregs[24][31]), .B(_09027_), .Y(_13747_));
NAND_g _20274_ (.A(cpuregs[28][31]), .B(_00007_[2]), .Y(_13748_));
AND_g _20275_ (.A(_09025_), .B(_13748_), .Y(_13749_));
NAND_g _20276_ (.A(_13747_), .B(_13749_), .Y(_13750_));
AND_g _20277_ (.A(_00007_[3]), .B(_13750_), .Y(_13751_));
NAND_g _20278_ (.A(_13746_), .B(_13751_), .Y(_13752_));
NAND_g _20279_ (.A(cpuregs[21][31]), .B(_00007_[2]), .Y(_13753_));
NAND_g _20280_ (.A(cpuregs[17][31]), .B(_09027_), .Y(_13754_));
AND_g _20281_ (.A(_00007_[0]), .B(_13754_), .Y(_13755_));
NAND_g _20282_ (.A(_13753_), .B(_13755_), .Y(_13756_));
NAND_g _20283_ (.A(cpuregs[20][31]), .B(_00007_[2]), .Y(_13757_));
NAND_g _20284_ (.A(cpuregs[16][31]), .B(_09027_), .Y(_13758_));
AND_g _20285_ (.A(_09025_), .B(_13758_), .Y(_13759_));
NAND_g _20286_ (.A(_13757_), .B(_13759_), .Y(_13760_));
AND_g _20287_ (.A(_09028_), .B(_13760_), .Y(_13761_));
NAND_g _20288_ (.A(_13756_), .B(_13761_), .Y(_13762_));
AND_g _20289_ (.A(_09026_), .B(_13762_), .Y(_13763_));
NAND_g _20290_ (.A(_13752_), .B(_13763_), .Y(_13764_));
NAND_g _20291_ (.A(cpuregs[27][31]), .B(_09027_), .Y(_13765_));
NAND_g _20292_ (.A(cpuregs[31][31]), .B(_00007_[2]), .Y(_13766_));
AND_g _20293_ (.A(_00007_[0]), .B(_13766_), .Y(_13767_));
NAND_g _20294_ (.A(_13765_), .B(_13767_), .Y(_13768_));
NAND_g _20295_ (.A(cpuregs[26][31]), .B(_09027_), .Y(_13769_));
NAND_g _20296_ (.A(cpuregs[30][31]), .B(_00007_[2]), .Y(_13770_));
AND_g _20297_ (.A(_09025_), .B(_13770_), .Y(_13771_));
NAND_g _20298_ (.A(_13769_), .B(_13771_), .Y(_13772_));
AND_g _20299_ (.A(_00007_[3]), .B(_13772_), .Y(_13773_));
NAND_g _20300_ (.A(_13768_), .B(_13773_), .Y(_13774_));
NAND_g _20301_ (.A(cpuregs[19][31]), .B(_09027_), .Y(_13775_));
NAND_g _20302_ (.A(cpuregs[23][31]), .B(_00007_[2]), .Y(_13776_));
AND_g _20303_ (.A(_00007_[0]), .B(_13776_), .Y(_13777_));
NAND_g _20304_ (.A(_13775_), .B(_13777_), .Y(_13778_));
NAND_g _20305_ (.A(cpuregs[18][31]), .B(_09027_), .Y(_13779_));
NAND_g _20306_ (.A(cpuregs[22][31]), .B(_00007_[2]), .Y(_13780_));
AND_g _20307_ (.A(_09025_), .B(_13780_), .Y(_13781_));
NAND_g _20308_ (.A(_13779_), .B(_13781_), .Y(_13782_));
AND_g _20309_ (.A(_09028_), .B(_13782_), .Y(_13783_));
NAND_g _20310_ (.A(_13778_), .B(_13783_), .Y(_13784_));
AND_g _20311_ (.A(_00007_[1]), .B(_13784_), .Y(_13785_));
NAND_g _20312_ (.A(_13774_), .B(_13785_), .Y(_13786_));
NAND_g _20313_ (.A(_13764_), .B(_13786_), .Y(_13787_));
NAND_g _20314_ (.A(_00007_[4]), .B(_13787_), .Y(_13788_));
NAND_g _20315_ (.A(cpuregs[13][31]), .B(_00007_[2]), .Y(_13789_));
NAND_g _20316_ (.A(cpuregs[9][31]), .B(_09027_), .Y(_13790_));
AND_g _20317_ (.A(_00007_[0]), .B(_13790_), .Y(_13791_));
NAND_g _20318_ (.A(_13789_), .B(_13791_), .Y(_13792_));
NAND_g _20319_ (.A(cpuregs[8][31]), .B(_09027_), .Y(_13793_));
NAND_g _20320_ (.A(cpuregs[12][31]), .B(_00007_[2]), .Y(_13794_));
AND_g _20321_ (.A(_09025_), .B(_13794_), .Y(_13795_));
NAND_g _20322_ (.A(_13793_), .B(_13795_), .Y(_13796_));
AND_g _20323_ (.A(_00007_[3]), .B(_13796_), .Y(_13797_));
NAND_g _20324_ (.A(_13792_), .B(_13797_), .Y(_13798_));
NAND_g _20325_ (.A(cpuregs[1][31]), .B(_09027_), .Y(_13799_));
NAND_g _20326_ (.A(cpuregs[5][31]), .B(_00007_[2]), .Y(_13800_));
AND_g _20327_ (.A(_00007_[0]), .B(_13800_), .Y(_13801_));
NAND_g _20328_ (.A(_13799_), .B(_13801_), .Y(_13802_));
NAND_g _20329_ (.A(cpuregs[0][31]), .B(_09027_), .Y(_13803_));
NAND_g _20330_ (.A(cpuregs[4][31]), .B(_00007_[2]), .Y(_13804_));
AND_g _20331_ (.A(_09025_), .B(_13804_), .Y(_13805_));
NAND_g _20332_ (.A(_13803_), .B(_13805_), .Y(_13806_));
AND_g _20333_ (.A(_09028_), .B(_13802_), .Y(_13807_));
NAND_g _20334_ (.A(_13806_), .B(_13807_), .Y(_13808_));
NAND_g _20335_ (.A(cpuregs[3][31]), .B(_09027_), .Y(_13809_));
NAND_g _20336_ (.A(cpuregs[7][31]), .B(_00007_[2]), .Y(_13810_));
AND_g _20337_ (.A(_00007_[0]), .B(_13810_), .Y(_13811_));
NAND_g _20338_ (.A(_13809_), .B(_13811_), .Y(_13812_));
NAND_g _20339_ (.A(cpuregs[2][31]), .B(_09027_), .Y(_13813_));
NAND_g _20340_ (.A(cpuregs[6][31]), .B(_00007_[2]), .Y(_13814_));
AND_g _20341_ (.A(_09025_), .B(_13814_), .Y(_13815_));
NAND_g _20342_ (.A(_13813_), .B(_13815_), .Y(_13816_));
AND_g _20343_ (.A(_09028_), .B(_13812_), .Y(_13817_));
NAND_g _20344_ (.A(_13816_), .B(_13817_), .Y(_13818_));
NAND_g _20345_ (.A(cpuregs[15][31]), .B(_00007_[2]), .Y(_13819_));
NAND_g _20346_ (.A(cpuregs[11][31]), .B(_09027_), .Y(_13820_));
AND_g _20347_ (.A(_00007_[0]), .B(_13820_), .Y(_13821_));
NAND_g _20348_ (.A(_13819_), .B(_13821_), .Y(_13822_));
NAND_g _20349_ (.A(cpuregs[10][31]), .B(_09027_), .Y(_13823_));
NAND_g _20350_ (.A(cpuregs[14][31]), .B(_00007_[2]), .Y(_13824_));
AND_g _20351_ (.A(_09025_), .B(_13824_), .Y(_13825_));
NAND_g _20352_ (.A(_13823_), .B(_13825_), .Y(_13826_));
AND_g _20353_ (.A(_00007_[3]), .B(_13826_), .Y(_13827_));
NAND_g _20354_ (.A(_13822_), .B(_13827_), .Y(_13828_));
NAND_g _20355_ (.A(_13818_), .B(_13828_), .Y(_13829_));
NAND_g _20356_ (.A(_00007_[1]), .B(_13829_), .Y(_13830_));
NAND_g _20357_ (.A(_13798_), .B(_13808_), .Y(_13831_));
NAND_g _20358_ (.A(_09026_), .B(_13831_), .Y(_13832_));
AND_g _20359_ (.A(_13830_), .B(_13832_), .Y(_13833_));
NAND_g _20360_ (.A(_09029_), .B(_13833_), .Y(_13834_));
AND_g _20361_ (.A(_13788_), .B(_13834_), .Y(_13835_));
NAND_g _20362_ (.A(_11170_), .B(_13835_), .Y(_13836_));
NAND_g _20363_ (.A(decoded_imm[31]), .B(_10606_), .Y(_13837_));
AND_g _20364_ (.A(_10603_), .B(_13837_), .Y(_13838_));
NAND_g _20365_ (.A(_13836_), .B(_13838_), .Y(_13839_));
AND_g _20366_ (.A(_13742_), .B(_13839_), .Y(_00306_));
AND_g _20367_ (.A(decoder_trigger), .B(_09024_), .Y(_13840_));
NAND_g _20368_ (.A(decoder_trigger), .B(_09024_), .Y(_13841_));
NAND_g _20369_ (.A(instr_sw), .B(_13841_), .Y(_13842_));
NAND_g _20370_ (.A(_08865_), .B(mem_rdata_q[13]), .Y(_13843_));
NOR_g _20371_ (.A(mem_rdata_q[14]), .B(_13843_), .Y(_13844_));
AND_g _20372_ (.A(is_sb_sh_sw), .B(_13840_), .Y(_13845_));
NAND_g _20373_ (.A(_13844_), .B(_13845_), .Y(_13846_));
NAND_g _20374_ (.A(_13842_), .B(_13846_), .Y(_00307_));
AND_g _20375_ (.A(resetn), .B(_09908_), .Y(_13847_));
NAND_g _20376_ (.A(resetn), .B(_09908_), .Y(_13848_));
AND_g _20377_ (.A(_08807_), .B(_13847_), .Y(_13849_));
NOT_g _20378_ (.A(_13849_), .Y(_13850_));
AND_g _20379_ (.A(_09070_), .B(_10592_), .Y(_13851_));
AND_g _20380_ (.A(_09068_), .B(_13851_), .Y(_13852_));
NAND_g _20381_ (.A(cpu_state[0]), .B(_13852_), .Y(_13853_));
NOR_g _20382_ (.A(cpu_state[1]), .B(_13853_), .Y(_13854_));
NOT_g _20383_ (.A(_13854_), .Y(_13855_));
NAND_g _20384_ (.A(cpu_state[1]), .B(_13852_), .Y(_13856_));
NOR_g _20385_ (.A(cpu_state[0]), .B(_13856_), .Y(_13857_));
NOT_g _20386_ (.A(_13857_), .Y(_13858_));
NOR_g _20387_ (.A(_13854_), .B(_13857_), .Y(_13859_));
NAND_g _20388_ (.A(_13855_), .B(_13858_), .Y(_13860_));
NAND_g _20389_ (.A(_13849_), .B(_13860_), .Y(_13861_));
NOT_g _20390_ (.A(_13861_), .Y(_00308_));
NOR_g _20391_ (.A(_08807_), .B(_10605_), .Y(_13862_));
AND_g _20392_ (.A(is_lb_lh_lw_lbu_lhu), .B(_10748_), .Y(_13863_));
NOR_g _20393_ (.A(_13862_), .B(_13863_), .Y(_13864_));
NAND_g _20394_ (.A(_08804_), .B(is_sll_srl_sra), .Y(_13865_));
NAND_g _20395_ (.A(_08807_), .B(_08862_), .Y(_13866_));
NAND_g _20396_ (.A(_13865_), .B(_13866_), .Y(_13867_));
NAND_g _20397_ (.A(_08864_), .B(_13867_), .Y(_13868_));
AND_g _20398_ (.A(_10605_), .B(_13868_), .Y(_13869_));
NAND_g _20399_ (.A(_10752_), .B(_13869_), .Y(_13870_));
NAND_g _20400_ (.A(_13864_), .B(_13870_), .Y(_13871_));
NAND_g _20401_ (.A(_10595_), .B(_13871_), .Y(_13872_));
NAND_g _20402_ (.A(_10595_), .B(_10751_), .Y(_13873_));
AND_g _20403_ (.A(_09067_), .B(_13851_), .Y(_13874_));
NOR_g _20404_ (.A(_09019_), .B(cpu_state[3]), .Y(_13875_));
AND_g _20405_ (.A(_13874_), .B(_13875_), .Y(_13876_));
NAND_g _20406_ (.A(_13874_), .B(_13875_), .Y(_13877_));
NOR_g _20407_ (.A(reg_sh[3]), .B(reg_sh[2]), .Y(_13878_));
AND_g _20408_ (.A(_09022_), .B(_13878_), .Y(_13879_));
NAND_g _20409_ (.A(_09022_), .B(_13878_), .Y(_13880_));
NAND_g _20410_ (.A(_09021_), .B(_13879_), .Y(_13881_));
NOR_g _20411_ (.A(reg_sh[1]), .B(_13881_), .Y(_13882_));
NOR_g _20412_ (.A(_13877_), .B(_13882_), .Y(_13883_));
NOT_g _20413_ (.A(_13883_), .Y(_13884_));
AND_g _20414_ (.A(_09074_), .B(_10601_), .Y(_13885_));
NAND_g _20415_ (.A(_13877_), .B(_13885_), .Y(_13886_));
AND_g _20416_ (.A(_13884_), .B(_13886_), .Y(_13887_));
AND_g _20417_ (.A(_13873_), .B(_13887_), .Y(_13888_));
AND_g _20418_ (.A(_13876_), .B(_13882_), .Y(_13889_));
NAND_g _20419_ (.A(mem_do_prefetch), .B(_13889_), .Y(_13890_));
NAND_g _20420_ (.A(_09073_), .B(_09892_), .Y(_13891_));
NAND_g _20421_ (.A(_10599_), .B(_13868_), .Y(_13892_));
AND_g _20422_ (.A(_13891_), .B(_13892_), .Y(_13893_));
AND_g _20423_ (.A(_13890_), .B(_13893_), .Y(_13894_));
AND_g _20424_ (.A(_13888_), .B(_13894_), .Y(_13895_));
NAND_g _20425_ (.A(_13872_), .B(_13895_), .Y(_13896_));
NOR_g _20426_ (.A(mem_do_rinst), .B(_13888_), .Y(_13897_));
NOR_g _20427_ (.A(_09910_), .B(_13897_), .Y(_13898_));
NAND_g _20428_ (.A(_13896_), .B(_13898_), .Y(_13899_));
AND_g _20429_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(resetn), .Y(_13900_));
NOR_g _20430_ (.A(pcpi_rs2[31]), .B(pcpi_rs1[31]), .Y(_13901_));
NAND_g _20431_ (.A(pcpi_rs2[31]), .B(pcpi_rs1[31]), .Y(_13902_));
XOR_g _20432_ (.A(pcpi_rs2[31]), .B(pcpi_rs1[31]), .Y(_13903_));
XNOR_g _20433_ (.A(pcpi_rs2[31]), .B(pcpi_rs1[31]), .Y(_13904_));
NAND_g _20434_ (.A(_08840_), .B(pcpi_rs1[30]), .Y(_13905_));
NOT_g _20435_ (.A(_13905_), .Y(_13906_));
NOR_g _20436_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_13907_));
NAND_g _20437_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_13908_));
XOR_g _20438_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_13909_));
XNOR_g _20439_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_13910_));
NAND_g _20440_ (.A(_08839_), .B(pcpi_rs1[29]), .Y(_13911_));
NOR_g _20441_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_13912_));
NOT_g _20442_ (.A(_13912_), .Y(_13913_));
NAND_g _20443_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_13914_));
XOR_g _20444_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_13915_));
XNOR_g _20445_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_13916_));
AND_g _20446_ (.A(_08838_), .B(pcpi_rs1[28]), .Y(_13917_));
NAND_g _20447_ (.A(_13916_), .B(_13917_), .Y(_13918_));
AND_g _20448_ (.A(_13911_), .B(_13918_), .Y(_13919_));
NAND_g _20449_ (.A(_13911_), .B(_13918_), .Y(_13920_));
NOR_g _20450_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_13921_));
NAND_g _20451_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_13922_));
XOR_g _20452_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_13923_));
XNOR_g _20453_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_13924_));
NOR_g _20454_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_13925_));
NOT_g _20455_ (.A(_13925_), .Y(_13926_));
NAND_g _20456_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_13927_));
XOR_g _20457_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_13928_));
XNOR_g _20458_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_13929_));
NOR_g _20459_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_13930_));
NAND_g _20460_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_13931_));
XOR_g _20461_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_13932_));
XNOR_g _20462_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_13933_));
AND_g _20463_ (.A(_13929_), .B(_13933_), .Y(_13934_));
NAND_g _20464_ (.A(_08835_), .B(pcpi_rs1[25]), .Y(_13935_));
NOR_g _20465_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_13936_));
NAND_g _20466_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_13937_));
XOR_g _20467_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_13938_));
XNOR_g _20468_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_13939_));
AND_g _20469_ (.A(_08834_), .B(pcpi_rs1[24]), .Y(_13940_));
NAND_g _20470_ (.A(_13939_), .B(_13940_), .Y(_13941_));
AND_g _20471_ (.A(_13935_), .B(_13941_), .Y(_13942_));
NAND_g _20472_ (.A(_13935_), .B(_13941_), .Y(_13943_));
NAND_g _20473_ (.A(_13934_), .B(_13943_), .Y(_13944_));
AND_g _20474_ (.A(_08836_), .B(pcpi_rs1[26]), .Y(_13945_));
NAND_g _20475_ (.A(_08836_), .B(pcpi_rs1[26]), .Y(_13946_));
NAND_g _20476_ (.A(_13929_), .B(_13945_), .Y(_13947_));
NAND_g _20477_ (.A(_08837_), .B(pcpi_rs1[27]), .Y(_13948_));
AND_g _20478_ (.A(_13944_), .B(_13948_), .Y(_13949_));
AND_g _20479_ (.A(_13947_), .B(_13949_), .Y(_13950_));
NAND_g _20480_ (.A(_13947_), .B(_13949_), .Y(_13951_));
NOR_g _20481_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_13952_));
NAND_g _20482_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_13953_));
XOR_g _20483_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_13954_));
XNOR_g _20484_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_13955_));
NOR_g _20485_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_13956_));
NOT_g _20486_ (.A(_13956_), .Y(_13957_));
NAND_g _20487_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_13958_));
XOR_g _20488_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_13959_));
XNOR_g _20489_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_13960_));
AND_g _20490_ (.A(_13955_), .B(_13960_), .Y(_13961_));
NAND_g _20491_ (.A(_08831_), .B(pcpi_rs1[21]), .Y(_13962_));
NOR_g _20492_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_13963_));
NOT_g _20493_ (.A(_13963_), .Y(_13964_));
NAND_g _20494_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_13965_));
XOR_g _20495_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_13966_));
XNOR_g _20496_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_13967_));
AND_g _20497_ (.A(_08830_), .B(pcpi_rs1[20]), .Y(_13968_));
NAND_g _20498_ (.A(_08830_), .B(pcpi_rs1[20]), .Y(_13969_));
NAND_g _20499_ (.A(_13967_), .B(_13968_), .Y(_13970_));
AND_g _20500_ (.A(_13962_), .B(_13970_), .Y(_13971_));
NAND_g _20501_ (.A(_13962_), .B(_13970_), .Y(_13972_));
NAND_g _20502_ (.A(_13961_), .B(_13972_), .Y(_13973_));
AND_g _20503_ (.A(_08832_), .B(pcpi_rs1[22]), .Y(_13974_));
NAND_g _20504_ (.A(_08832_), .B(pcpi_rs1[22]), .Y(_13975_));
NAND_g _20505_ (.A(_13955_), .B(_13974_), .Y(_13976_));
NAND_g _20506_ (.A(_08833_), .B(pcpi_rs1[23]), .Y(_13977_));
AND_g _20507_ (.A(_13976_), .B(_13977_), .Y(_13978_));
AND_g _20508_ (.A(_13973_), .B(_13978_), .Y(_13979_));
NAND_g _20509_ (.A(_08829_), .B(pcpi_rs1[19]), .Y(_13980_));
NOR_g _20510_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_13981_));
NOT_g _20511_ (.A(_13981_), .Y(_13982_));
NAND_g _20512_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_13983_));
XOR_g _20513_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_13984_));
XNOR_g _20514_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_13985_));
NAND_g _20515_ (.A(_08828_), .B(pcpi_rs1[18]), .Y(_13986_));
NOR_g _20516_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_13987_));
NOT_g _20517_ (.A(_13987_), .Y(_13988_));
NAND_g _20518_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_13989_));
XOR_g _20519_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_13990_));
XNOR_g _20520_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_13991_));
NAND_g _20521_ (.A(_08827_), .B(pcpi_rs1[17]), .Y(_13992_));
NOR_g _20522_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_13993_));
NAND_g _20523_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_13994_));
XOR_g _20524_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_13995_));
XNOR_g _20525_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_13996_));
AND_g _20526_ (.A(_08826_), .B(pcpi_rs1[16]), .Y(_13997_));
NAND_g _20527_ (.A(_13996_), .B(_13997_), .Y(_13998_));
AND_g _20528_ (.A(_13992_), .B(_13998_), .Y(_13999_));
NAND_g _20529_ (.A(_13992_), .B(_13998_), .Y(_14000_));
NAND_g _20530_ (.A(_13991_), .B(_14000_), .Y(_14001_));
NAND_g _20531_ (.A(_13986_), .B(_14001_), .Y(_14002_));
NAND_g _20532_ (.A(_13985_), .B(_14002_), .Y(_14003_));
AND_g _20533_ (.A(_13980_), .B(_14003_), .Y(_14004_));
NAND_g _20534_ (.A(_13980_), .B(_14003_), .Y(_14005_));
NOR_g _20535_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_14006_));
AND_g _20536_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_14007_));
NAND_g _20537_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_14008_));
XOR_g _20538_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_14009_));
XNOR_g _20539_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_14010_));
NOR_g _20540_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_14011_));
AND_g _20541_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_14012_));
NAND_g _20542_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_14013_));
XNOR_g _20543_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_14014_));
AND_g _20544_ (.A(_14010_), .B(_14014_), .Y(_14015_));
NOR_g _20545_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_14016_));
NAND_g _20546_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_14017_));
XOR_g _20547_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_14018_));
XNOR_g _20548_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_14019_));
NOR_g _20549_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_14020_));
NAND_g _20550_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_14021_));
XOR_g _20551_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_14022_));
XNOR_g _20552_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_14023_));
AND_g _20553_ (.A(_14019_), .B(_14023_), .Y(_14024_));
AND_g _20554_ (.A(_14015_), .B(_14024_), .Y(_14025_));
NOR_g _20555_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_14026_));
NAND_g _20556_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_14027_));
XOR_g _20557_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_14028_));
XNOR_g _20558_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_14029_));
NOR_g _20559_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_14030_));
NAND_g _20560_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_14031_));
XOR_g _20561_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_14032_));
XNOR_g _20562_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_14033_));
AND_g _20563_ (.A(_14029_), .B(_14033_), .Y(_14034_));
NOR_g _20564_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_14035_));
NAND_g _20565_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_14036_));
XOR_g _20566_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_14037_));
XNOR_g _20567_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_14038_));
NOR_g _20568_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_14039_));
NAND_g _20569_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_14040_));
XOR_g _20570_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_14041_));
XNOR_g _20571_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_14042_));
AND_g _20572_ (.A(_14038_), .B(_14042_), .Y(_14043_));
AND_g _20573_ (.A(_14034_), .B(_14043_), .Y(_14044_));
AND_g _20574_ (.A(_14025_), .B(_14044_), .Y(_14045_));
NAND_g _20575_ (.A(pcpi_rs2[7]), .B(_08962_), .Y(_14046_));
NOR_g _20576_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_14047_));
AND_g _20577_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_14048_));
NAND_g _20578_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_14049_));
XOR_g _20579_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_14050_));
XNOR_g _20580_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_14051_));
NAND_g _20581_ (.A(_08815_), .B(pcpi_rs1[5]), .Y(_14052_));
NOR_g _20582_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_14053_));
AND_g _20583_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_14054_));
NAND_g _20584_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_14055_));
XNOR_g _20585_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_14056_));
NOR_g _20586_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_14057_));
AND_g _20587_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_14058_));
NAND_g _20588_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_14059_));
XOR_g _20589_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_14060_));
XNOR_g _20590_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_14061_));
NAND_g _20591_ (.A(_08813_), .B(pcpi_rs1[2]), .Y(_14062_));
NOR_g _20592_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_14063_));
AND_g _20593_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_14064_));
NAND_g _20594_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_14065_));
XOR_g _20595_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_14066_));
XNOR_g _20596_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_14067_));
NAND_g _20597_ (.A(_08812_), .B(pcpi_rs1[1]), .Y(_14068_));
NOR_g _20598_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_14069_));
AND_g _20599_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_14070_));
NAND_g _20600_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_14071_));
XOR_g _20601_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_14072_));
XNOR_g _20602_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_14073_));
NOR_g _20603_ (.A(pcpi_rs2[0]), .B(pcpi_rs1[0]), .Y(_14074_));
NAND_g _20604_ (.A(pcpi_rs2[0]), .B(pcpi_rs1[0]), .Y(_14075_));
XNOR_g _20605_ (.A(pcpi_rs2[0]), .B(pcpi_rs1[0]), .Y(_14076_));
NAND_g _20606_ (.A(pcpi_rs2[0]), .B(_08961_), .Y(_14077_));
NAND_g _20607_ (.A(_14073_), .B(_14077_), .Y(_14078_));
NAND_g _20608_ (.A(_14068_), .B(_14078_), .Y(_14079_));
NAND_g _20609_ (.A(_14067_), .B(_14079_), .Y(_14080_));
NAND_g _20610_ (.A(_14062_), .B(_14080_), .Y(_14081_));
NAND_g _20611_ (.A(pcpi_rs1[3]), .B(_14081_), .Y(_14082_));
AND_g _20612_ (.A(pcpi_rs2[3]), .B(_14082_), .Y(_14083_));
NOR_g _20613_ (.A(pcpi_rs1[3]), .B(_14081_), .Y(_14084_));
NOR_g _20614_ (.A(_14083_), .B(_14084_), .Y(_14085_));
NAND_g _20615_ (.A(_14061_), .B(_14085_), .Y(_14086_));
NAND_g _20616_ (.A(_08814_), .B(pcpi_rs1[4]), .Y(_14087_));
NAND_g _20617_ (.A(_14086_), .B(_14087_), .Y(_14088_));
NAND_g _20618_ (.A(_14056_), .B(_14088_), .Y(_14089_));
NAND_g _20619_ (.A(_14052_), .B(_14089_), .Y(_14090_));
NAND_g _20620_ (.A(_14051_), .B(_14090_), .Y(_14091_));
NAND_g _20621_ (.A(_08816_), .B(pcpi_rs1[6]), .Y(_14092_));
NAND_g _20622_ (.A(_08817_), .B(pcpi_rs1[7]), .Y(_14093_));
AND_g _20623_ (.A(_14092_), .B(_14093_), .Y(_14094_));
NAND_g _20624_ (.A(_14091_), .B(_14094_), .Y(_14095_));
AND_g _20625_ (.A(_14046_), .B(_14095_), .Y(_14096_));
NAND_g _20626_ (.A(_14045_), .B(_14096_), .Y(_14097_));
NAND_g _20627_ (.A(_08823_), .B(pcpi_rs1[13]), .Y(_14098_));
AND_g _20628_ (.A(_08822_), .B(pcpi_rs1[12]), .Y(_14099_));
NAND_g _20629_ (.A(_08822_), .B(pcpi_rs1[12]), .Y(_14100_));
NAND_g _20630_ (.A(_14029_), .B(_14099_), .Y(_14101_));
AND_g _20631_ (.A(_14098_), .B(_14101_), .Y(_14102_));
NAND_g _20632_ (.A(_08819_), .B(pcpi_rs1[9]), .Y(_14103_));
NAND_g _20633_ (.A(_08818_), .B(pcpi_rs1[8]), .Y(_14104_));
NOT_g _20634_ (.A(_14104_), .Y(_14105_));
NAND_g _20635_ (.A(_14019_), .B(_14105_), .Y(_14106_));
NAND_g _20636_ (.A(_14103_), .B(_14106_), .Y(_14107_));
NAND_g _20637_ (.A(_14015_), .B(_14107_), .Y(_14108_));
AND_g _20638_ (.A(_08820_), .B(pcpi_rs1[10]), .Y(_14109_));
NAND_g _20639_ (.A(_14010_), .B(_14109_), .Y(_14110_));
NAND_g _20640_ (.A(_08821_), .B(pcpi_rs1[11]), .Y(_14111_));
AND_g _20641_ (.A(_14110_), .B(_14111_), .Y(_14112_));
AND_g _20642_ (.A(_14108_), .B(_14112_), .Y(_14113_));
NOT_g _20643_ (.A(_14113_), .Y(_14114_));
NAND_g _20644_ (.A(_14034_), .B(_14114_), .Y(_14115_));
NAND_g _20645_ (.A(_14102_), .B(_14115_), .Y(_14116_));
NAND_g _20646_ (.A(_14043_), .B(_14116_), .Y(_14117_));
NAND_g _20647_ (.A(_08825_), .B(pcpi_rs1[15]), .Y(_14118_));
AND_g _20648_ (.A(_08824_), .B(pcpi_rs1[14]), .Y(_14119_));
NAND_g _20649_ (.A(_08824_), .B(pcpi_rs1[14]), .Y(_14120_));
NAND_g _20650_ (.A(_14038_), .B(_14119_), .Y(_14121_));
AND_g _20651_ (.A(_14118_), .B(_14121_), .Y(_14122_));
AND_g _20652_ (.A(_14117_), .B(_14122_), .Y(_14123_));
NAND_g _20653_ (.A(_14097_), .B(_14123_), .Y(_14124_));
AND_g _20654_ (.A(_13985_), .B(_13991_), .Y(_14125_));
NOR_g _20655_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_14126_));
NAND_g _20656_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_14127_));
XOR_g _20657_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_14128_));
NOR_g _20658_ (.A(_13995_), .B(_14128_), .Y(_14129_));
AND_g _20659_ (.A(_14125_), .B(_14129_), .Y(_14130_));
NAND_g _20660_ (.A(_14124_), .B(_14129_), .Y(_14131_));
NAND_g _20661_ (.A(_14124_), .B(_14130_), .Y(_14132_));
NAND_g _20662_ (.A(_14004_), .B(_14132_), .Y(_14133_));
NOR_g _20663_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_14134_));
NAND_g _20664_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_14135_));
XOR_g _20665_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_14136_));
XNOR_g _20666_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_14137_));
AND_g _20667_ (.A(_14133_), .B(_14137_), .Y(_14138_));
NAND_g _20668_ (.A(_13967_), .B(_14138_), .Y(_14139_));
AND_g _20669_ (.A(_13967_), .B(_14137_), .Y(_14140_));
AND_g _20670_ (.A(_13961_), .B(_14140_), .Y(_14141_));
NAND_g _20671_ (.A(_14133_), .B(_14141_), .Y(_14142_));
NAND_g _20672_ (.A(_13979_), .B(_14142_), .Y(_14143_));
NOR_g _20673_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_14144_));
NAND_g _20674_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_14145_));
XOR_g _20675_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_14146_));
XNOR_g _20676_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_14147_));
AND_g _20677_ (.A(_13939_), .B(_14147_), .Y(_14148_));
AND_g _20678_ (.A(_14143_), .B(_14148_), .Y(_14149_));
NAND_g _20679_ (.A(_14143_), .B(_14148_), .Y(_14150_));
NAND_g _20680_ (.A(_13934_), .B(_14149_), .Y(_14151_));
NAND_g _20681_ (.A(_13950_), .B(_14151_), .Y(_14152_));
AND_g _20682_ (.A(_13924_), .B(_14152_), .Y(_14153_));
NAND_g _20683_ (.A(_13924_), .B(_14152_), .Y(_14154_));
NAND_g _20684_ (.A(_13916_), .B(_14153_), .Y(_14155_));
NAND_g _20685_ (.A(_13919_), .B(_14155_), .Y(_14156_));
NAND_g _20686_ (.A(_13910_), .B(_14156_), .Y(_14157_));
AND_g _20687_ (.A(_13905_), .B(_14157_), .Y(_14158_));
NAND_g _20688_ (.A(_13905_), .B(_14157_), .Y(_14159_));
AND_g _20689_ (.A(_13904_), .B(_13910_), .Y(_14160_));
AND_g _20690_ (.A(_13916_), .B(_13924_), .Y(_14161_));
AND_g _20691_ (.A(_14160_), .B(_14161_), .Y(_14162_));
AND_g _20692_ (.A(_13934_), .B(_14148_), .Y(_14163_));
AND_g _20693_ (.A(_14162_), .B(_14163_), .Y(_14164_));
AND_g _20694_ (.A(_14130_), .B(_14141_), .Y(_14165_));
AND_g _20695_ (.A(_14164_), .B(_14165_), .Y(_14166_));
NAND_g _20696_ (.A(_14124_), .B(_14166_), .Y(_14167_));
NAND_g _20697_ (.A(_14005_), .B(_14141_), .Y(_14168_));
NAND_g _20698_ (.A(_13979_), .B(_14168_), .Y(_14169_));
NAND_g _20699_ (.A(_14164_), .B(_14169_), .Y(_14170_));
NAND_g _20700_ (.A(_13951_), .B(_14162_), .Y(_14171_));
NAND_g _20701_ (.A(_08841_), .B(pcpi_rs1[31]), .Y(_14172_));
NAND_g _20702_ (.A(_13920_), .B(_14160_), .Y(_14173_));
AND_g _20703_ (.A(_14172_), .B(_14173_), .Y(_14174_));
AND_g _20704_ (.A(_14171_), .B(_14174_), .Y(_14175_));
AND_g _20705_ (.A(_14170_), .B(_14175_), .Y(_14176_));
AND_g _20706_ (.A(_14167_), .B(_14176_), .Y(_14177_));
NAND_g _20707_ (.A(_13904_), .B(_14158_), .Y(_14178_));
NAND_g _20708_ (.A(_14172_), .B(_14178_), .Y(_14179_));
AND_g _20709_ (.A(_14172_), .B(_14178_), .Y(_14180_));
NAND_g _20710_ (.A(instr_bge), .B(_14180_), .Y(_14181_));
NAND_g _20711_ (.A(is_slti_blt_slt), .B(_14179_), .Y(_14182_));
NAND_g _20712_ (.A(_13904_), .B(_13906_), .Y(_14183_));
NAND_g _20713_ (.A(_14177_), .B(_14183_), .Y(_14184_));
AND_g _20714_ (.A(_14177_), .B(_14183_), .Y(_14185_));
NAND_g _20715_ (.A(is_sltiu_bltu_sltu), .B(_14185_), .Y(_14186_));
AND_g _20716_ (.A(_14073_), .B(_14076_), .Y(_14187_));
NOR_g _20717_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_14188_));
AND_g _20718_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_14189_));
NAND_g _20719_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_14190_));
XOR_g _20720_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_14191_));
XNOR_g _20721_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_14192_));
NOR_g _20722_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_14193_));
NAND_g _20723_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_14194_));
XOR_g _20724_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_14195_));
NOR_g _20725_ (.A(_14191_), .B(_14195_), .Y(_14196_));
AND_g _20726_ (.A(_14187_), .B(_14196_), .Y(_14197_));
AND_g _20727_ (.A(_14051_), .B(_14056_), .Y(_14198_));
AND_g _20728_ (.A(_14061_), .B(_14067_), .Y(_14199_));
AND_g _20729_ (.A(_14198_), .B(_14199_), .Y(_14200_));
AND_g _20730_ (.A(_14197_), .B(_14200_), .Y(_14201_));
AND_g _20731_ (.A(_14045_), .B(_14201_), .Y(_14202_));
AND_g _20732_ (.A(_14166_), .B(_14202_), .Y(_14203_));
NAND_g _20733_ (.A(_14166_), .B(_14202_), .Y(_14204_));
NAND_g _20734_ (.A(instr_beq), .B(_14203_), .Y(_14205_));
NAND_g _20735_ (.A(instr_bne), .B(_14204_), .Y(_14206_));
AND_g _20736_ (.A(_14205_), .B(_14206_), .Y(_14207_));
NAND_g _20737_ (.A(instr_bgeu), .B(_14184_), .Y(_14208_));
AND_g _20738_ (.A(_14207_), .B(_14208_), .Y(_14209_));
AND_g _20739_ (.A(_14186_), .B(_14209_), .Y(_14210_));
AND_g _20740_ (.A(_14182_), .B(_14210_), .Y(_14211_));
NAND_g _20741_ (.A(_14181_), .B(_14211_), .Y(_14212_));
AND_g _20742_ (.A(_09019_), .B(cpu_state[3]), .Y(_14213_));
AND_g _20743_ (.A(_13874_), .B(_14213_), .Y(_14214_));
NAND_g _20744_ (.A(_13874_), .B(_14213_), .Y(_14215_));
AND_g _20745_ (.A(cpu_state[3]), .B(_13874_), .Y(_14216_));
AND_g _20746_ (.A(_09019_), .B(_14216_), .Y(_14217_));
NOT_g _20747_ (.A(_14217_), .Y(_14218_));
AND_g _20748_ (.A(_14212_), .B(_14217_), .Y(_14219_));
NAND_g _20749_ (.A(_13900_), .B(_14219_), .Y(_14220_));
AND_g _20750_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(_14217_), .Y(_14221_));
NAND_g _20751_ (.A(_13899_), .B(_14220_), .Y(_00309_));
NAND_g _20752_ (.A(mem_do_prefetch), .B(_13848_), .Y(_14222_));
AND_g _20753_ (.A(_13854_), .B(_14222_), .Y(_14223_));
AND_g _20754_ (.A(_08803_), .B(_14223_), .Y(_14224_));
NAND_g _20755_ (.A(_08803_), .B(_14223_), .Y(_14225_));
AND_g _20756_ (.A(resetn), .B(_14224_), .Y(_14226_));
NOT_g _20757_ (.A(_14226_), .Y(_14227_));
NAND_g _20758_ (.A(mem_do_rdata), .B(_09909_), .Y(_14228_));
NAND_g _20759_ (.A(_14227_), .B(_14228_), .Y(_00310_));
AND_g _20760_ (.A(_13857_), .B(_14222_), .Y(_14229_));
AND_g _20761_ (.A(_08789_), .B(_14229_), .Y(_14230_));
NOT_g _20762_ (.A(_14230_), .Y(_14231_));
AND_g _20763_ (.A(mem_do_wdata), .B(_09907_), .Y(_14232_));
NOR_g _20764_ (.A(_14230_), .B(_14232_), .Y(_14233_));
NOR_g _20765_ (.A(_08811_), .B(_14233_), .Y(_00311_));
NAND_g _20766_ (.A(mem_do_wdata), .B(_14229_), .Y(_14234_));
NOR_g _20767_ (.A(_13859_), .B(_14222_), .Y(_14235_));
NOR_g _20768_ (.A(_08811_), .B(_14235_), .Y(_14236_));
AND_g _20769_ (.A(_14234_), .B(_14236_), .Y(_14237_));
NAND_g _20770_ (.A(_09074_), .B(_13859_), .Y(_14238_));
NAND_g _20771_ (.A(mem_do_rdata), .B(_14223_), .Y(_14239_));
AND_g _20772_ (.A(_14238_), .B(_14239_), .Y(_14240_));
AND_g _20773_ (.A(_14237_), .B(_14240_), .Y(_14241_));
NOR_g _20774_ (.A(instr_lb), .B(instr_lbu), .Y(_14242_));
NAND_g _20775_ (.A(_10726_), .B(_14230_), .Y(_14243_));
NOR_g _20776_ (.A(instr_sb), .B(_14243_), .Y(_14244_));
AND_g _20777_ (.A(_10740_), .B(_14242_), .Y(_14245_));
NAND_g _20778_ (.A(_14224_), .B(_14245_), .Y(_14246_));
NOR_g _20779_ (.A(instr_lw), .B(_14246_), .Y(_14247_));
NOR_g _20780_ (.A(_14244_), .B(_14247_), .Y(_14248_));
AND_g _20781_ (.A(_14241_), .B(_14248_), .Y(_14249_));
NOR_g _20782_ (.A(_10740_), .B(_14225_), .Y(_14250_));
AND_g _20783_ (.A(instr_sh), .B(_14230_), .Y(_14251_));
NOR_g _20784_ (.A(_14250_), .B(_14251_), .Y(_14252_));
AND_g _20785_ (.A(_14249_), .B(_14252_), .Y(_14253_));
NOR_g _20786_ (.A(mem_wordsize[0]), .B(_14249_), .Y(_14254_));
NOR_g _20787_ (.A(_14253_), .B(_14254_), .Y(_00312_));
NOR_g _20788_ (.A(_14225_), .B(_14242_), .Y(_14255_));
AND_g _20789_ (.A(instr_sb), .B(_14230_), .Y(_14256_));
NOR_g _20790_ (.A(_14255_), .B(_14256_), .Y(_14257_));
AND_g _20791_ (.A(_14249_), .B(_14257_), .Y(_14258_));
NOR_g _20792_ (.A(mem_wordsize[1]), .B(_14249_), .Y(_14259_));
NOR_g _20793_ (.A(_14258_), .B(_14259_), .Y(_00313_));
NOR_g _20794_ (.A(_08811_), .B(trap), .Y(_14260_));
AND_g _20795_ (.A(_09901_), .B(_14260_), .Y(_14261_));
NOR_g _20796_ (.A(mem_do_rinst), .B(mem_do_prefetch), .Y(_14262_));
NAND_g _20797_ (.A(_08804_), .B(_08807_), .Y(_14263_));
NOR_g _20798_ (.A(mem_do_wdata), .B(mem_do_rdata), .Y(_14264_));
NAND_g _20799_ (.A(_08803_), .B(_14262_), .Y(_14265_));
AND_g _20800_ (.A(_14262_), .B(_14264_), .Y(_14266_));
NAND_g _20801_ (.A(_14262_), .B(_14264_), .Y(_14267_));
AND_g _20802_ (.A(mem_do_wdata), .B(_09901_), .Y(_14268_));
AND_g _20803_ (.A(resetn), .B(_14268_), .Y(mem_la_write));
AND_g _20804_ (.A(_09901_), .B(_14265_), .Y(_14269_));
AND_g _20805_ (.A(resetn), .B(_14269_), .Y(mem_la_read));
AND_g _20806_ (.A(_14261_), .B(_14267_), .Y(_14270_));
NAND_g _20807_ (.A(_14261_), .B(_14267_), .Y(_14271_));
AND_g _20808_ (.A(_09897_), .B(_14260_), .Y(_14272_));
NAND_g _20809_ (.A(resetn), .B(trap), .Y(_14273_));
NOR_g _20810_ (.A(mem_ready), .B(_14273_), .Y(_14274_));
NOR_g _20811_ (.A(_14272_), .B(_14274_), .Y(_14275_));
NOR_g _20812_ (.A(_09897_), .B(_09903_), .Y(_14276_));
AND_g _20813_ (.A(_09902_), .B(_14260_), .Y(_14277_));
NAND_g _20814_ (.A(_14276_), .B(_14277_), .Y(_14278_));
NAND_g _20815_ (.A(_14261_), .B(_14266_), .Y(_14279_));
AND_g _20816_ (.A(_14278_), .B(_14279_), .Y(_14280_));
AND_g _20817_ (.A(_08789_), .B(_14261_), .Y(_14281_));
NAND_g _20818_ (.A(_14275_), .B(_14280_), .Y(_14282_));
NAND_g _20819_ (.A(mem_valid), .B(_14282_), .Y(_14283_));
NAND_g _20820_ (.A(_14271_), .B(_14283_), .Y(_00314_));
AND_g _20821_ (.A(_08854_), .B(_09497_), .Y(_14284_));
AND_g _20822_ (.A(latched_rd[2]), .B(_14284_), .Y(_14285_));
AND_g _20823_ (.A(_09083_), .B(_09084_), .Y(_14286_));
AND_g _20824_ (.A(_14285_), .B(_14286_), .Y(_14287_));
NAND_g _20825_ (.A(_14285_), .B(_14286_), .Y(_14288_));
NAND_g _20826_ (.A(_09098_), .B(_14287_), .Y(_14289_));
NAND_g _20827_ (.A(cpuregs[20][0]), .B(_14288_), .Y(_14290_));
NAND_g _20828_ (.A(_14289_), .B(_14290_), .Y(_00315_));
NAND_g _20829_ (.A(_09109_), .B(_14287_), .Y(_14291_));
NAND_g _20830_ (.A(cpuregs[20][1]), .B(_14288_), .Y(_14292_));
NAND_g _20831_ (.A(_14291_), .B(_14292_), .Y(_00316_));
NAND_g _20832_ (.A(_09118_), .B(_14287_), .Y(_14293_));
NAND_g _20833_ (.A(cpuregs[20][2]), .B(_14288_), .Y(_14294_));
NAND_g _20834_ (.A(_14293_), .B(_14294_), .Y(_00317_));
NAND_g _20835_ (.A(_09131_), .B(_14287_), .Y(_14295_));
NAND_g _20836_ (.A(cpuregs[20][3]), .B(_14288_), .Y(_14296_));
NAND_g _20837_ (.A(_14295_), .B(_14296_), .Y(_00318_));
NAND_g _20838_ (.A(_09144_), .B(_14287_), .Y(_14297_));
NAND_g _20839_ (.A(cpuregs[20][4]), .B(_14288_), .Y(_14298_));
NAND_g _20840_ (.A(_14297_), .B(_14298_), .Y(_00319_));
NAND_g _20841_ (.A(_09157_), .B(_14287_), .Y(_14299_));
NAND_g _20842_ (.A(cpuregs[20][5]), .B(_14288_), .Y(_14300_));
NAND_g _20843_ (.A(_14299_), .B(_14300_), .Y(_00320_));
NAND_g _20844_ (.A(_09170_), .B(_14287_), .Y(_14301_));
NAND_g _20845_ (.A(cpuregs[20][6]), .B(_14288_), .Y(_14302_));
NAND_g _20846_ (.A(_14301_), .B(_14302_), .Y(_00321_));
NAND_g _20847_ (.A(_09183_), .B(_14287_), .Y(_14303_));
NAND_g _20848_ (.A(cpuregs[20][7]), .B(_14288_), .Y(_14304_));
NAND_g _20849_ (.A(_14303_), .B(_14304_), .Y(_00322_));
NAND_g _20850_ (.A(_09196_), .B(_14287_), .Y(_14305_));
NAND_g _20851_ (.A(cpuregs[20][8]), .B(_14288_), .Y(_14306_));
NAND_g _20852_ (.A(_14305_), .B(_14306_), .Y(_00323_));
NAND_g _20853_ (.A(_09209_), .B(_14287_), .Y(_14307_));
NAND_g _20854_ (.A(cpuregs[20][9]), .B(_14288_), .Y(_14308_));
NAND_g _20855_ (.A(_14307_), .B(_14308_), .Y(_00324_));
NAND_g _20856_ (.A(_09222_), .B(_14287_), .Y(_14309_));
NAND_g _20857_ (.A(cpuregs[20][10]), .B(_14288_), .Y(_14310_));
NAND_g _20858_ (.A(_14309_), .B(_14310_), .Y(_00325_));
NAND_g _20859_ (.A(_09235_), .B(_14287_), .Y(_14311_));
NAND_g _20860_ (.A(cpuregs[20][11]), .B(_14288_), .Y(_14312_));
NAND_g _20861_ (.A(_14311_), .B(_14312_), .Y(_00326_));
NAND_g _20862_ (.A(_09248_), .B(_14287_), .Y(_14313_));
NAND_g _20863_ (.A(cpuregs[20][12]), .B(_14288_), .Y(_14314_));
NAND_g _20864_ (.A(_14313_), .B(_14314_), .Y(_00327_));
NAND_g _20865_ (.A(_09261_), .B(_14287_), .Y(_14315_));
NAND_g _20866_ (.A(cpuregs[20][13]), .B(_14288_), .Y(_14316_));
NAND_g _20867_ (.A(_14315_), .B(_14316_), .Y(_00328_));
NAND_g _20868_ (.A(_09274_), .B(_14287_), .Y(_14317_));
NAND_g _20869_ (.A(cpuregs[20][14]), .B(_14288_), .Y(_14318_));
NAND_g _20870_ (.A(_14317_), .B(_14318_), .Y(_00329_));
NAND_g _20871_ (.A(_09287_), .B(_14287_), .Y(_14319_));
NAND_g _20872_ (.A(cpuregs[20][15]), .B(_14288_), .Y(_14320_));
NAND_g _20873_ (.A(_14319_), .B(_14320_), .Y(_00330_));
NAND_g _20874_ (.A(_09300_), .B(_14287_), .Y(_14321_));
NAND_g _20875_ (.A(cpuregs[20][16]), .B(_14288_), .Y(_14322_));
NAND_g _20876_ (.A(_14321_), .B(_14322_), .Y(_00331_));
NOR_g _20877_ (.A(cpuregs[20][17]), .B(_14287_), .Y(_14323_));
NOR_g _20878_ (.A(_09313_), .B(_14288_), .Y(_14324_));
NOR_g _20879_ (.A(_14323_), .B(_14324_), .Y(_00332_));
NOR_g _20880_ (.A(cpuregs[20][18]), .B(_14287_), .Y(_14325_));
NOR_g _20881_ (.A(_09325_), .B(_14288_), .Y(_14326_));
NOR_g _20882_ (.A(_14325_), .B(_14326_), .Y(_00333_));
NAND_g _20883_ (.A(_09338_), .B(_14287_), .Y(_14327_));
NAND_g _20884_ (.A(cpuregs[20][19]), .B(_14288_), .Y(_14328_));
NAND_g _20885_ (.A(_14327_), .B(_14328_), .Y(_00334_));
NAND_g _20886_ (.A(_09351_), .B(_14287_), .Y(_14329_));
NAND_g _20887_ (.A(cpuregs[20][20]), .B(_14288_), .Y(_14330_));
NAND_g _20888_ (.A(_14329_), .B(_14330_), .Y(_00335_));
NAND_g _20889_ (.A(_09364_), .B(_14287_), .Y(_14331_));
NAND_g _20890_ (.A(cpuregs[20][21]), .B(_14288_), .Y(_14332_));
NAND_g _20891_ (.A(_14331_), .B(_14332_), .Y(_00336_));
NAND_g _20892_ (.A(_09377_), .B(_14287_), .Y(_14333_));
NAND_g _20893_ (.A(cpuregs[20][22]), .B(_14288_), .Y(_14334_));
NAND_g _20894_ (.A(_14333_), .B(_14334_), .Y(_00337_));
NAND_g _20895_ (.A(_09390_), .B(_14287_), .Y(_14335_));
NAND_g _20896_ (.A(cpuregs[20][23]), .B(_14288_), .Y(_14336_));
NAND_g _20897_ (.A(_14335_), .B(_14336_), .Y(_00338_));
NAND_g _20898_ (.A(_09403_), .B(_14287_), .Y(_14337_));
NAND_g _20899_ (.A(cpuregs[20][24]), .B(_14288_), .Y(_14338_));
NAND_g _20900_ (.A(_14337_), .B(_14338_), .Y(_00339_));
NAND_g _20901_ (.A(_09416_), .B(_14287_), .Y(_14339_));
NAND_g _20902_ (.A(cpuregs[20][25]), .B(_14288_), .Y(_14340_));
NAND_g _20903_ (.A(_14339_), .B(_14340_), .Y(_00340_));
NAND_g _20904_ (.A(_09429_), .B(_14287_), .Y(_14341_));
NAND_g _20905_ (.A(cpuregs[20][26]), .B(_14288_), .Y(_14342_));
NAND_g _20906_ (.A(_14341_), .B(_14342_), .Y(_00341_));
NAND_g _20907_ (.A(_09442_), .B(_14287_), .Y(_14343_));
NAND_g _20908_ (.A(cpuregs[20][27]), .B(_14288_), .Y(_14344_));
NAND_g _20909_ (.A(_14343_), .B(_14344_), .Y(_00342_));
NAND_g _20910_ (.A(_09455_), .B(_14287_), .Y(_14345_));
NAND_g _20911_ (.A(cpuregs[20][28]), .B(_14288_), .Y(_14346_));
NAND_g _20912_ (.A(_14345_), .B(_14346_), .Y(_00343_));
NAND_g _20913_ (.A(_09468_), .B(_14287_), .Y(_14347_));
NAND_g _20914_ (.A(cpuregs[20][29]), .B(_14288_), .Y(_14348_));
NAND_g _20915_ (.A(_14347_), .B(_14348_), .Y(_00344_));
NAND_g _20916_ (.A(_09481_), .B(_14287_), .Y(_14349_));
NAND_g _20917_ (.A(cpuregs[20][30]), .B(_14288_), .Y(_14350_));
NAND_g _20918_ (.A(_14349_), .B(_14350_), .Y(_00345_));
NAND_g _20919_ (.A(_09493_), .B(_14287_), .Y(_14351_));
NAND_g _20920_ (.A(cpuregs[20][31]), .B(_14288_), .Y(_14352_));
NAND_g _20921_ (.A(_14351_), .B(_14352_), .Y(_00346_));
AND_g _20922_ (.A(_09074_), .B(_14215_), .Y(_14353_));
NAND_g _20923_ (.A(latched_store), .B(_14353_), .Y(_14354_));
NAND_g _20924_ (.A(_10595_), .B(_10710_), .Y(_14355_));
NOR_g _20925_ (.A(_13854_), .B(_13876_), .Y(_14356_));
AND_g _20926_ (.A(_08790_), .B(_14217_), .Y(_14357_));
NOT_g _20927_ (.A(_14357_), .Y(_14358_));
NAND_g _20928_ (.A(_14356_), .B(_14358_), .Y(_14359_));
AND_g _20929_ (.A(_14354_), .B(_14355_), .Y(_14360_));
NOR_g _20930_ (.A(_14219_), .B(_14359_), .Y(_14361_));
NAND_g _20931_ (.A(_14360_), .B(_14361_), .Y(_14362_));
AND_g _20932_ (.A(resetn), .B(_14362_), .Y(_00347_));
NOR_g _20933_ (.A(latched_stalu), .B(_14357_), .Y(_14363_));
NOT_g _20934_ (.A(_14363_), .Y(_14364_));
AND_g _20935_ (.A(_09920_), .B(_14364_), .Y(_00348_));
NAND_g _20936_ (.A(latched_branch), .B(_14353_), .Y(_14365_));
NAND_g _20937_ (.A(instr_jal), .B(_09893_), .Y(_14366_));
NAND_g _20938_ (.A(instr_jalr), .B(_14357_), .Y(_14367_));
AND_g _20939_ (.A(_14365_), .B(_14366_), .Y(_14368_));
NAND_g _20940_ (.A(_14367_), .B(_14368_), .Y(_14369_));
NAND_g _20941_ (.A(resetn), .B(_14369_), .Y(_14370_));
NAND_g _20942_ (.A(_14220_), .B(_14370_), .Y(_00349_));
NAND_g _20943_ (.A(is_lbu_lhu_lw), .B(_14226_), .Y(_14371_));
AND_g _20944_ (.A(_09074_), .B(_14225_), .Y(_14372_));
AND_g _20945_ (.A(latched_is_lu), .B(resetn), .Y(_14373_));
NAND_g _20946_ (.A(_14372_), .B(_14373_), .Y(_14374_));
NAND_g _20947_ (.A(_14371_), .B(_14374_), .Y(_00350_));
NAND_g _20948_ (.A(instr_lh), .B(_14226_), .Y(_14375_));
AND_g _20949_ (.A(latched_is_lh), .B(resetn), .Y(_14376_));
NAND_g _20950_ (.A(_14372_), .B(_14376_), .Y(_14377_));
NAND_g _20951_ (.A(_14375_), .B(_14377_), .Y(_00351_));
NAND_g _20952_ (.A(instr_lb), .B(_14226_), .Y(_14378_));
AND_g _20953_ (.A(latched_is_lb), .B(resetn), .Y(_14379_));
NAND_g _20954_ (.A(_14372_), .B(_14379_), .Y(_14380_));
NAND_g _20955_ (.A(_14378_), .B(_14380_), .Y(_00352_));
NOR_g _20956_ (.A(_08811_), .B(_14353_), .Y(_14381_));
NAND_g _20957_ (.A(_14358_), .B(_14381_), .Y(_14382_));
NAND_g _20958_ (.A(latched_rd[0]), .B(_14382_), .Y(_14383_));
NAND_g _20959_ (.A(decoded_rd[0]), .B(_09075_), .Y(_14384_));
NAND_g _20960_ (.A(_14383_), .B(_14384_), .Y(_00353_));
NAND_g _20961_ (.A(latched_rd[1]), .B(_14382_), .Y(_14385_));
NAND_g _20962_ (.A(decoded_rd[1]), .B(_09075_), .Y(_14386_));
NAND_g _20963_ (.A(_14385_), .B(_14386_), .Y(_00354_));
NAND_g _20964_ (.A(latched_rd[2]), .B(_14382_), .Y(_14387_));
NAND_g _20965_ (.A(decoded_rd[2]), .B(_09075_), .Y(_14388_));
NAND_g _20966_ (.A(_14387_), .B(_14388_), .Y(_00355_));
NAND_g _20967_ (.A(latched_rd[3]), .B(_14382_), .Y(_14389_));
NAND_g _20968_ (.A(decoded_rd[3]), .B(_09075_), .Y(_14390_));
NAND_g _20969_ (.A(_14389_), .B(_14390_), .Y(_00356_));
NAND_g _20970_ (.A(latched_rd[4]), .B(_14382_), .Y(_14391_));
NAND_g _20971_ (.A(decoded_rd[4]), .B(_09075_), .Y(_14392_));
NAND_g _20972_ (.A(_14391_), .B(_14392_), .Y(_00357_));
AND_g _20973_ (.A(mem_do_rinst), .B(_13847_), .Y(_14393_));
NAND_g _20974_ (.A(mem_do_rinst), .B(_13847_), .Y(_14394_));
NAND_g _20975_ (.A(mem_rdata[0]), .B(_09903_), .Y(_14395_));
NAND_g _20976_ (.A(mem_rdata_q[0]), .B(_09904_), .Y(_14396_));
NAND_g _20977_ (.A(_14395_), .B(_14396_), .Y(_00514_));
NAND_g _20978_ (.A(mem_rdata[1]), .B(_09903_), .Y(_14397_));
NAND_g _20979_ (.A(mem_rdata_q[1]), .B(_09904_), .Y(_14398_));
NAND_g _20980_ (.A(_14397_), .B(_14398_), .Y(_00515_));
AND_g _20981_ (.A(_00514_), .B(_00515_), .Y(_14399_));
NAND_g _20982_ (.A(mem_rdata[2]), .B(_09903_), .Y(_14400_));
NAND_g _20983_ (.A(mem_rdata_q[2]), .B(_09904_), .Y(_14401_));
NAND_g _20984_ (.A(_14400_), .B(_14401_), .Y(_00516_));
AND_g _20985_ (.A(_14399_), .B(_00516_), .Y(_14402_));
NAND_g _20986_ (.A(mem_rdata[3]), .B(_09903_), .Y(_14403_));
NAND_g _20987_ (.A(mem_rdata_q[3]), .B(_09904_), .Y(_14404_));
AND_g _20988_ (.A(_14403_), .B(_14404_), .Y(_14405_));
NOT_g _20989_ (.A(_14405_), .Y(_00517_));
AND_g _20990_ (.A(_14402_), .B(_14405_), .Y(_14406_));
NAND_g _20991_ (.A(mem_rdata[6]), .B(_09903_), .Y(_14407_));
NAND_g _20992_ (.A(mem_rdata_q[6]), .B(_09904_), .Y(_14408_));
AND_g _20993_ (.A(_14407_), .B(_14408_), .Y(_14409_));
NOT_g _20994_ (.A(_14409_), .Y(_00520_));
NAND_g _20995_ (.A(mem_rdata[4]), .B(_09903_), .Y(_14410_));
NAND_g _20996_ (.A(mem_rdata_q[4]), .B(_09904_), .Y(_14411_));
AND_g _20997_ (.A(_14410_), .B(_14411_), .Y(_14412_));
NOT_g _20998_ (.A(_14412_), .Y(_00518_));
AND_g _20999_ (.A(_14409_), .B(_00518_), .Y(_14413_));
NAND_g _21000_ (.A(mem_rdata[5]), .B(_09903_), .Y(_14414_));
NAND_g _21001_ (.A(mem_rdata_q[5]), .B(_09904_), .Y(_14415_));
AND_g _21002_ (.A(_14414_), .B(_14415_), .Y(_14416_));
NOT_g _21003_ (.A(_14416_), .Y(_00519_));
AND_g _21004_ (.A(_14413_), .B(_00519_), .Y(_14417_));
NAND_g _21005_ (.A(_14406_), .B(_14417_), .Y(_14418_));
NAND_g _21006_ (.A(_14393_), .B(_14418_), .Y(_14419_));
NAND_g _21007_ (.A(_08855_), .B(_14394_), .Y(_14420_));
AND_g _21008_ (.A(_14419_), .B(_14420_), .Y(_00358_));
AND_g _21009_ (.A(_14413_), .B(_14416_), .Y(_14421_));
NAND_g _21010_ (.A(_14406_), .B(_14421_), .Y(_14422_));
NAND_g _21011_ (.A(_14393_), .B(_14422_), .Y(_14423_));
NAND_g _21012_ (.A(_08856_), .B(_14394_), .Y(_14424_));
AND_g _21013_ (.A(_14423_), .B(_14424_), .Y(_00359_));
AND_g _21014_ (.A(_00520_), .B(_14412_), .Y(_14425_));
AND_g _21015_ (.A(_00519_), .B(_14425_), .Y(_14426_));
AND_g _21016_ (.A(_14402_), .B(_00517_), .Y(_14427_));
NAND_g _21017_ (.A(_14426_), .B(_14427_), .Y(_14428_));
NAND_g _21018_ (.A(_14393_), .B(_14428_), .Y(_14429_));
NAND_g _21019_ (.A(_08857_), .B(_14394_), .Y(_14430_));
AND_g _21020_ (.A(_14429_), .B(_14430_), .Y(_00360_));
AND_g _21021_ (.A(resetn), .B(_13841_), .Y(_14431_));
NAND_g _21022_ (.A(instr_beq), .B(_14431_), .Y(_14432_));
NOR_g _21023_ (.A(mem_rdata_q[12]), .B(mem_rdata_q[13]), .Y(_14433_));
AND_g _21024_ (.A(_08867_), .B(_14433_), .Y(_14434_));
AND_g _21025_ (.A(_13840_), .B(_13900_), .Y(_14435_));
NAND_g _21026_ (.A(_14434_), .B(_14435_), .Y(_14436_));
NAND_g _21027_ (.A(_14432_), .B(_14436_), .Y(_00361_));
NAND_g _21028_ (.A(mem_rdata_q[12]), .B(_08866_), .Y(_14437_));
NOR_g _21029_ (.A(mem_rdata_q[14]), .B(_14437_), .Y(_14438_));
NAND_g _21030_ (.A(_14435_), .B(_14438_), .Y(_14439_));
NAND_g _21031_ (.A(instr_bne), .B(_14431_), .Y(_14440_));
NAND_g _21032_ (.A(_14439_), .B(_14440_), .Y(_00362_));
AND_g _21033_ (.A(mem_rdata_q[14]), .B(_14433_), .Y(_14441_));
NAND_g _21034_ (.A(_14435_), .B(_14441_), .Y(_14442_));
NAND_g _21035_ (.A(instr_blt), .B(_14431_), .Y(_14443_));
NAND_g _21036_ (.A(_14442_), .B(_14443_), .Y(_00363_));
NOR_g _21037_ (.A(_08867_), .B(_14437_), .Y(_14444_));
NAND_g _21038_ (.A(_14435_), .B(_14444_), .Y(_14445_));
NAND_g _21039_ (.A(instr_bge), .B(_14431_), .Y(_14446_));
NAND_g _21040_ (.A(_14445_), .B(_14446_), .Y(_00364_));
NOR_g _21041_ (.A(_08867_), .B(_13843_), .Y(_14447_));
NAND_g _21042_ (.A(_14435_), .B(_14447_), .Y(_14448_));
NAND_g _21043_ (.A(instr_bltu), .B(_14431_), .Y(_14449_));
NAND_g _21044_ (.A(_14448_), .B(_14449_), .Y(_00365_));
AND_g _21045_ (.A(mem_rdata_q[12]), .B(mem_rdata_q[13]), .Y(_14450_));
AND_g _21046_ (.A(mem_rdata_q[14]), .B(_14450_), .Y(_14451_));
NAND_g _21047_ (.A(_14435_), .B(_14451_), .Y(_14452_));
NAND_g _21048_ (.A(instr_bgeu), .B(_14431_), .Y(_14453_));
NAND_g _21049_ (.A(_14452_), .B(_14453_), .Y(_00366_));
NAND_g _21050_ (.A(instr_jalr), .B(_14394_), .Y(_14454_));
NAND_g _21051_ (.A(mem_rdata[14]), .B(_09903_), .Y(_14455_));
NAND_g _21052_ (.A(mem_rdata_q[14]), .B(_09904_), .Y(_14456_));
NAND_g _21053_ (.A(_14455_), .B(_14456_), .Y(_00428_));
NOR_g _21054_ (.A(_14394_), .B(_00428_), .Y(_14457_));
NAND_g _21055_ (.A(mem_rdata[13]), .B(_09903_), .Y(_14458_));
NAND_g _21056_ (.A(mem_rdata_q[13]), .B(_09904_), .Y(_14459_));
NAND_g _21057_ (.A(_14458_), .B(_14459_), .Y(_00427_));
NAND_g _21058_ (.A(mem_rdata[12]), .B(_09903_), .Y(_14460_));
NAND_g _21059_ (.A(mem_rdata_q[12]), .B(_09904_), .Y(_14461_));
NAND_g _21060_ (.A(_14460_), .B(_14461_), .Y(_00426_));
NOR_g _21061_ (.A(_00427_), .B(_00426_), .Y(_14462_));
AND_g _21062_ (.A(_14426_), .B(_14462_), .Y(_14463_));
AND_g _21063_ (.A(_14406_), .B(_14463_), .Y(_14464_));
NAND_g _21064_ (.A(_14457_), .B(_14464_), .Y(_14465_));
NAND_g _21065_ (.A(_14454_), .B(_14465_), .Y(_00367_));
NAND_g _21066_ (.A(instr_lb), .B(_13841_), .Y(_14466_));
AND_g _21067_ (.A(is_lb_lh_lw_lbu_lhu), .B(_13840_), .Y(_14467_));
NAND_g _21068_ (.A(_14434_), .B(_14467_), .Y(_14468_));
NAND_g _21069_ (.A(_14466_), .B(_14468_), .Y(_00368_));
NAND_g _21070_ (.A(instr_lh), .B(_13841_), .Y(_14469_));
NAND_g _21071_ (.A(_14438_), .B(_14467_), .Y(_14470_));
NAND_g _21072_ (.A(_14469_), .B(_14470_), .Y(_00369_));
NAND_g _21073_ (.A(instr_lw), .B(_13841_), .Y(_14471_));
NAND_g _21074_ (.A(_13844_), .B(_14467_), .Y(_14472_));
NAND_g _21075_ (.A(_14471_), .B(_14472_), .Y(_00370_));
NAND_g _21076_ (.A(instr_lbu), .B(_13841_), .Y(_14473_));
NAND_g _21077_ (.A(_14441_), .B(_14467_), .Y(_14474_));
NAND_g _21078_ (.A(_14473_), .B(_14474_), .Y(_00371_));
NAND_g _21079_ (.A(instr_lhu), .B(_13841_), .Y(_14475_));
NAND_g _21080_ (.A(_14444_), .B(_14467_), .Y(_14476_));
NAND_g _21081_ (.A(_14475_), .B(_14476_), .Y(_00372_));
NAND_g _21082_ (.A(_08791_), .B(_08860_), .Y(_14477_));
NAND_g _21083_ (.A(_13883_), .B(_14477_), .Y(_14478_));
AND_g _21084_ (.A(_13859_), .B(_13877_), .Y(_14479_));
NAND_g _21085_ (.A(_10596_), .B(_14479_), .Y(_14480_));
NAND_g _21086_ (.A(_08793_), .B(_08859_), .Y(_14481_));
NAND_g _21087_ (.A(_10723_), .B(_10741_), .Y(_14482_));
NOR_g _21088_ (.A(_14481_), .B(_14482_), .Y(_14483_));
AND_g _21089_ (.A(_13876_), .B(_14483_), .Y(_14484_));
NOR_g _21090_ (.A(_13889_), .B(_14484_), .Y(_14485_));
AND_g _21091_ (.A(_14480_), .B(_14485_), .Y(_14486_));
AND_g _21092_ (.A(_14239_), .B(_14486_), .Y(_14487_));
AND_g _21093_ (.A(_14237_), .B(_14487_), .Y(_14488_));
AND_g _21094_ (.A(_14478_), .B(_14488_), .Y(_14489_));
NOR_g _21095_ (.A(pcpi_rs1[31]), .B(_14489_), .Y(_14490_));
NAND_g _21096_ (.A(decoded_imm[30]), .B(pcpi_rs1[30]), .Y(_14491_));
XOR_g _21097_ (.A(decoded_imm[30]), .B(pcpi_rs1[30]), .Y(_14492_));
NAND_g _21098_ (.A(decoded_imm[29]), .B(pcpi_rs1[29]), .Y(_14493_));
NOR_g _21099_ (.A(decoded_imm[29]), .B(pcpi_rs1[29]), .Y(_14494_));
NAND_g _21100_ (.A(decoded_imm[28]), .B(pcpi_rs1[28]), .Y(_14495_));
XOR_g _21101_ (.A(decoded_imm[28]), .B(pcpi_rs1[28]), .Y(_14496_));
NOR_g _21102_ (.A(decoded_imm[27]), .B(pcpi_rs1[27]), .Y(_14497_));
NAND_g _21103_ (.A(decoded_imm[27]), .B(pcpi_rs1[27]), .Y(_14498_));
NAND_g _21104_ (.A(decoded_imm[26]), .B(pcpi_rs1[26]), .Y(_14499_));
XOR_g _21105_ (.A(decoded_imm[26]), .B(pcpi_rs1[26]), .Y(_14500_));
NAND_g _21106_ (.A(decoded_imm[25]), .B(pcpi_rs1[25]), .Y(_14501_));
NOR_g _21107_ (.A(decoded_imm[25]), .B(pcpi_rs1[25]), .Y(_14502_));
NAND_g _21108_ (.A(decoded_imm[24]), .B(pcpi_rs1[24]), .Y(_14503_));
XOR_g _21109_ (.A(decoded_imm[24]), .B(pcpi_rs1[24]), .Y(_14504_));
NAND_g _21110_ (.A(decoded_imm[23]), .B(pcpi_rs1[23]), .Y(_14505_));
NOR_g _21111_ (.A(decoded_imm[23]), .B(pcpi_rs1[23]), .Y(_14506_));
NAND_g _21112_ (.A(decoded_imm[22]), .B(pcpi_rs1[22]), .Y(_14507_));
XOR_g _21113_ (.A(decoded_imm[22]), .B(pcpi_rs1[22]), .Y(_14508_));
NAND_g _21114_ (.A(decoded_imm[21]), .B(pcpi_rs1[21]), .Y(_14509_));
NOR_g _21115_ (.A(decoded_imm[21]), .B(pcpi_rs1[21]), .Y(_14510_));
NAND_g _21116_ (.A(decoded_imm[20]), .B(pcpi_rs1[20]), .Y(_14511_));
XOR_g _21117_ (.A(decoded_imm[20]), .B(pcpi_rs1[20]), .Y(_14512_));
NOR_g _21118_ (.A(decoded_imm[19]), .B(pcpi_rs1[19]), .Y(_14513_));
NAND_g _21119_ (.A(decoded_imm[19]), .B(pcpi_rs1[19]), .Y(_14514_));
NAND_g _21120_ (.A(decoded_imm[18]), .B(pcpi_rs1[18]), .Y(_14515_));
XOR_g _21121_ (.A(decoded_imm[18]), .B(pcpi_rs1[18]), .Y(_14516_));
NAND_g _21122_ (.A(decoded_imm[17]), .B(pcpi_rs1[17]), .Y(_14517_));
NOR_g _21123_ (.A(decoded_imm[17]), .B(pcpi_rs1[17]), .Y(_14518_));
NAND_g _21124_ (.A(decoded_imm[16]), .B(pcpi_rs1[16]), .Y(_14519_));
XOR_g _21125_ (.A(decoded_imm[16]), .B(pcpi_rs1[16]), .Y(_14520_));
NAND_g _21126_ (.A(decoded_imm[15]), .B(pcpi_rs1[15]), .Y(_14521_));
NOR_g _21127_ (.A(decoded_imm[15]), .B(pcpi_rs1[15]), .Y(_14522_));
NAND_g _21128_ (.A(decoded_imm[14]), .B(pcpi_rs1[14]), .Y(_14523_));
XOR_g _21129_ (.A(decoded_imm[14]), .B(pcpi_rs1[14]), .Y(_14524_));
NAND_g _21130_ (.A(decoded_imm[13]), .B(pcpi_rs1[13]), .Y(_14525_));
NOR_g _21131_ (.A(decoded_imm[13]), .B(pcpi_rs1[13]), .Y(_14526_));
NAND_g _21132_ (.A(decoded_imm[12]), .B(pcpi_rs1[12]), .Y(_14527_));
XOR_g _21133_ (.A(decoded_imm[12]), .B(pcpi_rs1[12]), .Y(_14528_));
NAND_g _21134_ (.A(decoded_imm[11]), .B(pcpi_rs1[11]), .Y(_14529_));
NOR_g _21135_ (.A(decoded_imm[11]), .B(pcpi_rs1[11]), .Y(_14530_));
NAND_g _21136_ (.A(decoded_imm[10]), .B(pcpi_rs1[10]), .Y(_14531_));
XOR_g _21137_ (.A(decoded_imm[10]), .B(pcpi_rs1[10]), .Y(_14532_));
NAND_g _21138_ (.A(decoded_imm[9]), .B(pcpi_rs1[9]), .Y(_14533_));
NOR_g _21139_ (.A(decoded_imm[9]), .B(pcpi_rs1[9]), .Y(_14534_));
NAND_g _21140_ (.A(decoded_imm[8]), .B(pcpi_rs1[8]), .Y(_14535_));
XOR_g _21141_ (.A(decoded_imm[8]), .B(pcpi_rs1[8]), .Y(_14536_));
NAND_g _21142_ (.A(decoded_imm[7]), .B(pcpi_rs1[7]), .Y(_14537_));
NOR_g _21143_ (.A(decoded_imm[7]), .B(pcpi_rs1[7]), .Y(_14538_));
NAND_g _21144_ (.A(decoded_imm[6]), .B(pcpi_rs1[6]), .Y(_14539_));
XOR_g _21145_ (.A(decoded_imm[6]), .B(pcpi_rs1[6]), .Y(_14540_));
NAND_g _21146_ (.A(decoded_imm[5]), .B(pcpi_rs1[5]), .Y(_14541_));
NAND_g _21147_ (.A(decoded_imm[4]), .B(pcpi_rs1[4]), .Y(_14542_));
XOR_g _21148_ (.A(decoded_imm[4]), .B(pcpi_rs1[4]), .Y(_14543_));
NAND_g _21149_ (.A(decoded_imm[3]), .B(pcpi_rs1[3]), .Y(_14544_));
NOR_g _21150_ (.A(decoded_imm[3]), .B(pcpi_rs1[3]), .Y(_14545_));
NAND_g _21151_ (.A(decoded_imm[2]), .B(pcpi_rs1[2]), .Y(_14546_));
NAND_g _21152_ (.A(decoded_imm[1]), .B(pcpi_rs1[1]), .Y(_14547_));
AND_g _21153_ (.A(decoded_imm[0]), .B(pcpi_rs1[0]), .Y(_14548_));
NAND_g _21154_ (.A(decoded_imm[0]), .B(pcpi_rs1[0]), .Y(_14549_));
XOR_g _21155_ (.A(decoded_imm[1]), .B(pcpi_rs1[1]), .Y(_14550_));
NAND_g _21156_ (.A(_14548_), .B(_14550_), .Y(_14551_));
NAND_g _21157_ (.A(_14547_), .B(_14551_), .Y(_14552_));
XOR_g _21158_ (.A(decoded_imm[2]), .B(pcpi_rs1[2]), .Y(_14553_));
NAND_g _21159_ (.A(_14552_), .B(_14553_), .Y(_14554_));
AND_g _21160_ (.A(_14546_), .B(_14554_), .Y(_14555_));
AND_g _21161_ (.A(_14544_), .B(_14555_), .Y(_14556_));
NOR_g _21162_ (.A(_14545_), .B(_14556_), .Y(_14557_));
NAND_g _21163_ (.A(_14543_), .B(_14557_), .Y(_14558_));
NAND_g _21164_ (.A(_14542_), .B(_14558_), .Y(_14559_));
XOR_g _21165_ (.A(decoded_imm[5]), .B(pcpi_rs1[5]), .Y(_14560_));
NAND_g _21166_ (.A(_14559_), .B(_14560_), .Y(_14561_));
NAND_g _21167_ (.A(_14541_), .B(_14561_), .Y(_14562_));
NAND_g _21168_ (.A(_14540_), .B(_14562_), .Y(_14563_));
AND_g _21169_ (.A(_14539_), .B(_14563_), .Y(_14564_));
AND_g _21170_ (.A(_14537_), .B(_14564_), .Y(_14565_));
NOR_g _21171_ (.A(_14538_), .B(_14565_), .Y(_14566_));
NAND_g _21172_ (.A(_14536_), .B(_14566_), .Y(_14567_));
AND_g _21173_ (.A(_14535_), .B(_14567_), .Y(_14568_));
AND_g _21174_ (.A(_14533_), .B(_14568_), .Y(_14569_));
NOR_g _21175_ (.A(_14534_), .B(_14569_), .Y(_14570_));
NAND_g _21176_ (.A(_14532_), .B(_14570_), .Y(_14571_));
AND_g _21177_ (.A(_14531_), .B(_14571_), .Y(_14572_));
AND_g _21178_ (.A(_14529_), .B(_14572_), .Y(_14573_));
NOR_g _21179_ (.A(_14530_), .B(_14573_), .Y(_14574_));
NAND_g _21180_ (.A(_14528_), .B(_14574_), .Y(_14575_));
AND_g _21181_ (.A(_14527_), .B(_14575_), .Y(_14576_));
AND_g _21182_ (.A(_14525_), .B(_14576_), .Y(_14577_));
NOR_g _21183_ (.A(_14526_), .B(_14577_), .Y(_14578_));
NAND_g _21184_ (.A(_14524_), .B(_14578_), .Y(_14579_));
AND_g _21185_ (.A(_14523_), .B(_14579_), .Y(_14580_));
AND_g _21186_ (.A(_14521_), .B(_14580_), .Y(_14581_));
NOR_g _21187_ (.A(_14522_), .B(_14581_), .Y(_14582_));
NAND_g _21188_ (.A(_14520_), .B(_14582_), .Y(_14583_));
AND_g _21189_ (.A(_14519_), .B(_14583_), .Y(_14584_));
AND_g _21190_ (.A(_14517_), .B(_14584_), .Y(_14585_));
NOR_g _21191_ (.A(_14518_), .B(_14585_), .Y(_14586_));
NAND_g _21192_ (.A(_14516_), .B(_14586_), .Y(_14587_));
AND_g _21193_ (.A(_14515_), .B(_14587_), .Y(_14588_));
AND_g _21194_ (.A(_14514_), .B(_14588_), .Y(_14589_));
NOR_g _21195_ (.A(_14513_), .B(_14589_), .Y(_14590_));
NAND_g _21196_ (.A(_14512_), .B(_14590_), .Y(_14591_));
AND_g _21197_ (.A(_14511_), .B(_14591_), .Y(_14592_));
AND_g _21198_ (.A(_14509_), .B(_14592_), .Y(_14593_));
NOR_g _21199_ (.A(_14510_), .B(_14593_), .Y(_14594_));
NAND_g _21200_ (.A(_14508_), .B(_14594_), .Y(_14595_));
AND_g _21201_ (.A(_14507_), .B(_14595_), .Y(_14596_));
AND_g _21202_ (.A(_14505_), .B(_14596_), .Y(_14597_));
NOR_g _21203_ (.A(_14506_), .B(_14597_), .Y(_14598_));
NAND_g _21204_ (.A(_14504_), .B(_14598_), .Y(_14599_));
AND_g _21205_ (.A(_14503_), .B(_14599_), .Y(_14600_));
AND_g _21206_ (.A(_14501_), .B(_14600_), .Y(_14601_));
NOR_g _21207_ (.A(_14502_), .B(_14601_), .Y(_14602_));
NAND_g _21208_ (.A(_14500_), .B(_14602_), .Y(_14603_));
AND_g _21209_ (.A(_14499_), .B(_14603_), .Y(_14604_));
AND_g _21210_ (.A(_14498_), .B(_14604_), .Y(_14605_));
NOR_g _21211_ (.A(_14497_), .B(_14605_), .Y(_14606_));
NAND_g _21212_ (.A(_14496_), .B(_14606_), .Y(_14607_));
AND_g _21213_ (.A(_14495_), .B(_14607_), .Y(_14608_));
AND_g _21214_ (.A(_14493_), .B(_14608_), .Y(_14609_));
NOR_g _21215_ (.A(_14494_), .B(_14609_), .Y(_14610_));
NAND_g _21216_ (.A(_14492_), .B(_14610_), .Y(_14611_));
NAND_g _21217_ (.A(_14491_), .B(_14611_), .Y(_14612_));
XNOR_g _21218_ (.A(pcpi_rs1[31]), .B(decoded_imm[31]), .Y(_14613_));
NAND_g _21219_ (.A(_14225_), .B(_14231_), .Y(_14614_));
XNOR_g _21220_ (.A(_14612_), .B(_14613_), .Y(_14615_));
NAND_g _21221_ (.A(_14614_), .B(_14615_), .Y(_14616_));
AND_g _21222_ (.A(_08855_), .B(is_lui_auipc_jal), .Y(_14617_));
NAND_g _21223_ (.A(reg_pc[31]), .B(_14617_), .Y(_14618_));
NOR_g _21224_ (.A(decoded_imm_j[15]), .B(decoded_imm_j[16]), .Y(_14619_));
NOR_g _21225_ (.A(decoded_imm_j[17]), .B(decoded_imm_j[19]), .Y(_14620_));
NAND_g _21226_ (.A(_14619_), .B(_14620_), .Y(_14621_));
NOR_g _21227_ (.A(decoded_imm_j[18]), .B(_14621_), .Y(_14622_));
NOR_g _21228_ (.A(is_lui_auipc_jal), .B(_14622_), .Y(_14623_));
AND_g _21229_ (.A(_10750_), .B(_14623_), .Y(_14624_));
NAND_g _21230_ (.A(cpuregs[24][31]), .B(_09032_), .Y(_14625_));
NAND_g _21231_ (.A(cpuregs[28][31]), .B(_00008_[2]), .Y(_14626_));
AND_g _21232_ (.A(_09030_), .B(_14626_), .Y(_14627_));
NAND_g _21233_ (.A(_14625_), .B(_14627_), .Y(_14628_));
NAND_g _21234_ (.A(cpuregs[29][31]), .B(_00008_[2]), .Y(_14629_));
NAND_g _21235_ (.A(cpuregs[25][31]), .B(_09032_), .Y(_14630_));
AND_g _21236_ (.A(_00008_[0]), .B(_14630_), .Y(_14631_));
NAND_g _21237_ (.A(_14629_), .B(_14631_), .Y(_14632_));
AND_g _21238_ (.A(_14628_), .B(_14632_), .Y(_14633_));
NAND_g _21239_ (.A(cpuregs[26][31]), .B(_09032_), .Y(_14634_));
NAND_g _21240_ (.A(cpuregs[30][31]), .B(_00008_[2]), .Y(_14635_));
AND_g _21241_ (.A(_09030_), .B(_14635_), .Y(_14636_));
NAND_g _21242_ (.A(_14634_), .B(_14636_), .Y(_14637_));
NAND_g _21243_ (.A(cpuregs[31][31]), .B(_00008_[2]), .Y(_14638_));
NAND_g _21244_ (.A(cpuregs[27][31]), .B(_09032_), .Y(_14639_));
AND_g _21245_ (.A(_00008_[0]), .B(_14639_), .Y(_14640_));
NAND_g _21246_ (.A(_14638_), .B(_14640_), .Y(_14641_));
AND_g _21247_ (.A(_14637_), .B(_14641_), .Y(_14642_));
NAND_g _21248_ (.A(_00008_[1]), .B(_14642_), .Y(_14643_));
NAND_g _21249_ (.A(_09031_), .B(_14633_), .Y(_14644_));
NAND_g _21250_ (.A(_14643_), .B(_14644_), .Y(_14645_));
NAND_g _21251_ (.A(_00008_[4]), .B(_14645_), .Y(_14646_));
NAND_g _21252_ (.A(cpuregs[8][31]), .B(_09032_), .Y(_14647_));
NAND_g _21253_ (.A(cpuregs[12][31]), .B(_00008_[2]), .Y(_14648_));
AND_g _21254_ (.A(_09030_), .B(_14648_), .Y(_14649_));
NAND_g _21255_ (.A(_14647_), .B(_14649_), .Y(_14650_));
NAND_g _21256_ (.A(cpuregs[13][31]), .B(_00008_[2]), .Y(_14651_));
NAND_g _21257_ (.A(cpuregs[9][31]), .B(_09032_), .Y(_14652_));
AND_g _21258_ (.A(_00008_[0]), .B(_14652_), .Y(_14653_));
NAND_g _21259_ (.A(_14651_), .B(_14653_), .Y(_14654_));
NAND_g _21260_ (.A(_14650_), .B(_14654_), .Y(_14655_));
NAND_g _21261_ (.A(_09031_), .B(_14655_), .Y(_14656_));
NAND_g _21262_ (.A(cpuregs[10][31]), .B(_09032_), .Y(_14657_));
NAND_g _21263_ (.A(cpuregs[14][31]), .B(_00008_[2]), .Y(_14658_));
AND_g _21264_ (.A(_09030_), .B(_14658_), .Y(_14659_));
NAND_g _21265_ (.A(_14657_), .B(_14659_), .Y(_14660_));
NAND_g _21266_ (.A(cpuregs[15][31]), .B(_00008_[2]), .Y(_14661_));
NAND_g _21267_ (.A(cpuregs[11][31]), .B(_09032_), .Y(_14662_));
AND_g _21268_ (.A(_00008_[0]), .B(_14662_), .Y(_14663_));
NAND_g _21269_ (.A(_14661_), .B(_14663_), .Y(_14664_));
NAND_g _21270_ (.A(_14660_), .B(_14664_), .Y(_14665_));
AND_g _21271_ (.A(_00008_[1]), .B(_14665_), .Y(_14666_));
NOR_g _21272_ (.A(_00008_[4]), .B(_14666_), .Y(_14667_));
NAND_g _21273_ (.A(_14656_), .B(_14667_), .Y(_14668_));
NAND_g _21274_ (.A(_14646_), .B(_14668_), .Y(_14669_));
NAND_g _21275_ (.A(_00008_[3]), .B(_14669_), .Y(_14670_));
NAND_g _21276_ (.A(cpuregs[23][31]), .B(_00008_[2]), .Y(_14671_));
NAND_g _21277_ (.A(cpuregs[19][31]), .B(_09032_), .Y(_14672_));
NAND_g _21278_ (.A(_14671_), .B(_14672_), .Y(_14673_));
NAND_g _21279_ (.A(_00008_[0]), .B(_14673_), .Y(_14674_));
NAND_g _21280_ (.A(cpuregs[22][31]), .B(_00008_[2]), .Y(_14675_));
NAND_g _21281_ (.A(cpuregs[18][31]), .B(_09032_), .Y(_14676_));
NAND_g _21282_ (.A(_14675_), .B(_14676_), .Y(_14677_));
NAND_g _21283_ (.A(_09030_), .B(_14677_), .Y(_14678_));
NAND_g _21284_ (.A(_14674_), .B(_14678_), .Y(_14679_));
NAND_g _21285_ (.A(_00008_[1]), .B(_14679_), .Y(_14680_));
NAND_g _21286_ (.A(cpuregs[17][31]), .B(_09032_), .Y(_14681_));
NAND_g _21287_ (.A(cpuregs[21][31]), .B(_00008_[2]), .Y(_14682_));
NAND_g _21288_ (.A(_14681_), .B(_14682_), .Y(_14683_));
NAND_g _21289_ (.A(_00008_[0]), .B(_14683_), .Y(_14684_));
NAND_g _21290_ (.A(cpuregs[20][31]), .B(_00008_[2]), .Y(_14685_));
NAND_g _21291_ (.A(cpuregs[16][31]), .B(_09032_), .Y(_14686_));
NAND_g _21292_ (.A(_14685_), .B(_14686_), .Y(_14687_));
NAND_g _21293_ (.A(_09030_), .B(_14687_), .Y(_14688_));
NAND_g _21294_ (.A(_14684_), .B(_14688_), .Y(_14689_));
NAND_g _21295_ (.A(_09031_), .B(_14689_), .Y(_14690_));
NAND_g _21296_ (.A(_14680_), .B(_14690_), .Y(_14691_));
NAND_g _21297_ (.A(_00008_[4]), .B(_14691_), .Y(_14692_));
NAND_g _21298_ (.A(cpuregs[6][31]), .B(_00008_[2]), .Y(_14693_));
NAND_g _21299_ (.A(cpuregs[2][31]), .B(_09032_), .Y(_14694_));
NAND_g _21300_ (.A(_14693_), .B(_14694_), .Y(_14695_));
NAND_g _21301_ (.A(_09030_), .B(_14695_), .Y(_14696_));
NAND_g _21302_ (.A(cpuregs[7][31]), .B(_00008_[2]), .Y(_14697_));
NAND_g _21303_ (.A(cpuregs[3][31]), .B(_09032_), .Y(_14698_));
NAND_g _21304_ (.A(_14697_), .B(_14698_), .Y(_14699_));
NAND_g _21305_ (.A(_00008_[0]), .B(_14699_), .Y(_14700_));
AND_g _21306_ (.A(_14696_), .B(_14700_), .Y(_14701_));
NAND_g _21307_ (.A(cpuregs[1][31]), .B(_09032_), .Y(_14702_));
NAND_g _21308_ (.A(cpuregs[5][31]), .B(_00008_[2]), .Y(_14703_));
NAND_g _21309_ (.A(_14702_), .B(_14703_), .Y(_14704_));
NAND_g _21310_ (.A(_00008_[0]), .B(_14704_), .Y(_14705_));
NAND_g _21311_ (.A(cpuregs[4][31]), .B(_00008_[2]), .Y(_14706_));
NAND_g _21312_ (.A(cpuregs[0][31]), .B(_09032_), .Y(_14707_));
NAND_g _21313_ (.A(_14706_), .B(_14707_), .Y(_14708_));
NAND_g _21314_ (.A(_09030_), .B(_14708_), .Y(_14709_));
AND_g _21315_ (.A(_14705_), .B(_14709_), .Y(_14710_));
NAND_g _21316_ (.A(_00008_[1]), .B(_14701_), .Y(_14711_));
AND_g _21317_ (.A(_09031_), .B(_14710_), .Y(_14712_));
NOR_g _21318_ (.A(_00008_[4]), .B(_14712_), .Y(_14713_));
NAND_g _21319_ (.A(_14711_), .B(_14713_), .Y(_14714_));
NAND_g _21320_ (.A(_14692_), .B(_14714_), .Y(_14715_));
NAND_g _21321_ (.A(_09033_), .B(_14715_), .Y(_14716_));
NAND_g _21322_ (.A(_14670_), .B(_14716_), .Y(_14717_));
NAND_g _21323_ (.A(_14624_), .B(_14717_), .Y(_14718_));
NAND_g _21324_ (.A(_14618_), .B(_14718_), .Y(_14719_));
NAND_g _21325_ (.A(_10595_), .B(_14719_), .Y(_14720_));
AND_g _21326_ (.A(pcpi_rs1[27]), .B(_14481_), .Y(_14721_));
NAND_g _21327_ (.A(_13880_), .B(_14721_), .Y(_14722_));
AND_g _21328_ (.A(pcpi_rs1[30]), .B(_14481_), .Y(_14723_));
NAND_g _21329_ (.A(_13879_), .B(_14723_), .Y(_14724_));
NAND_g _21330_ (.A(_14722_), .B(_14724_), .Y(_14725_));
NAND_g _21331_ (.A(_13883_), .B(_14725_), .Y(_14726_));
AND_g _21332_ (.A(_14489_), .B(_14720_), .Y(_14727_));
AND_g _21333_ (.A(_14726_), .B(_14727_), .Y(_14728_));
AND_g _21334_ (.A(_14616_), .B(_14728_), .Y(_14729_));
NOR_g _21335_ (.A(_14490_), .B(_14729_), .Y(_00373_));
NAND_g _21336_ (.A(instr_sh), .B(_13841_), .Y(_14730_));
NAND_g _21337_ (.A(_13845_), .B(_14438_), .Y(_14731_));
NAND_g _21338_ (.A(_14730_), .B(_14731_), .Y(_00374_));
NAND_g _21339_ (.A(instr_addi), .B(_14431_), .Y(_14732_));
AND_g _21340_ (.A(is_alu_reg_imm), .B(_13840_), .Y(_14733_));
AND_g _21341_ (.A(resetn), .B(_14733_), .Y(_14734_));
NAND_g _21342_ (.A(_14434_), .B(_14734_), .Y(_14735_));
NAND_g _21343_ (.A(_14732_), .B(_14735_), .Y(_00375_));
NAND_g _21344_ (.A(instr_slti), .B(_14431_), .Y(_14736_));
NAND_g _21345_ (.A(_13844_), .B(_14734_), .Y(_14737_));
NAND_g _21346_ (.A(_14736_), .B(_14737_), .Y(_00376_));
AND_g _21347_ (.A(_08867_), .B(_14450_), .Y(_14738_));
NAND_g _21348_ (.A(_14734_), .B(_14738_), .Y(_14739_));
NAND_g _21349_ (.A(instr_sltiu), .B(_14431_), .Y(_14740_));
NAND_g _21350_ (.A(_14739_), .B(_14740_), .Y(_00377_));
NAND_g _21351_ (.A(instr_xori), .B(_14431_), .Y(_14741_));
NAND_g _21352_ (.A(_14441_), .B(_14734_), .Y(_14742_));
NAND_g _21353_ (.A(_14741_), .B(_14742_), .Y(_00378_));
NAND_g _21354_ (.A(instr_ori), .B(_14431_), .Y(_14743_));
NAND_g _21355_ (.A(_14447_), .B(_14734_), .Y(_14744_));
NAND_g _21356_ (.A(_14743_), .B(_14744_), .Y(_00379_));
NAND_g _21357_ (.A(instr_andi), .B(_14431_), .Y(_14745_));
NAND_g _21358_ (.A(_14451_), .B(_14734_), .Y(_14746_));
NAND_g _21359_ (.A(_14745_), .B(_14746_), .Y(_00380_));
NAND_g _21360_ (.A(instr_sb), .B(_13841_), .Y(_14747_));
NAND_g _21361_ (.A(_13845_), .B(_14434_), .Y(_14748_));
NAND_g _21362_ (.A(_14747_), .B(_14748_), .Y(_00381_));
NAND_g _21363_ (.A(instr_slli), .B(_13841_), .Y(_14749_));
NOR_g _21364_ (.A(mem_rdata_q[25]), .B(mem_rdata_q[26]), .Y(_14750_));
NOR_g _21365_ (.A(mem_rdata_q[27]), .B(mem_rdata_q[28]), .Y(_14751_));
AND_g _21366_ (.A(_08872_), .B(_14751_), .Y(_14752_));
AND_g _21367_ (.A(_14750_), .B(_14752_), .Y(_14753_));
AND_g _21368_ (.A(_08870_), .B(_14753_), .Y(_14754_));
AND_g _21369_ (.A(_08871_), .B(_14754_), .Y(_14755_));
AND_g _21370_ (.A(_14438_), .B(_14755_), .Y(_14756_));
NOT_g _21371_ (.A(_14756_), .Y(_14757_));
NAND_g _21372_ (.A(_14733_), .B(_14756_), .Y(_14758_));
NAND_g _21373_ (.A(_14749_), .B(_14758_), .Y(_00382_));
NAND_g _21374_ (.A(instr_srli), .B(_13841_), .Y(_14759_));
AND_g _21375_ (.A(is_alu_reg_imm), .B(_14444_), .Y(_14760_));
AND_g _21376_ (.A(_13840_), .B(_14755_), .Y(_14761_));
NAND_g _21377_ (.A(_14760_), .B(_14761_), .Y(_14762_));
NAND_g _21378_ (.A(_14759_), .B(_14762_), .Y(_00383_));
NAND_g _21379_ (.A(instr_add), .B(_14431_), .Y(_14763_));
AND_g _21380_ (.A(resetn), .B(is_alu_reg_reg), .Y(_14764_));
AND_g _21381_ (.A(_14434_), .B(_14764_), .Y(_14765_));
NAND_g _21382_ (.A(_14761_), .B(_14765_), .Y(_14766_));
NAND_g _21383_ (.A(_14763_), .B(_14766_), .Y(_00384_));
NAND_g _21384_ (.A(instr_sub), .B(_14431_), .Y(_14767_));
AND_g _21385_ (.A(_08870_), .B(mem_rdata_q[30]), .Y(_14768_));
AND_g _21386_ (.A(_13840_), .B(_14753_), .Y(_14769_));
AND_g _21387_ (.A(_14768_), .B(_14769_), .Y(_14770_));
NAND_g _21388_ (.A(_14765_), .B(_14770_), .Y(_14771_));
NAND_g _21389_ (.A(_14767_), .B(_14771_), .Y(_00385_));
NAND_g _21390_ (.A(instr_sll), .B(_14431_), .Y(_14772_));
AND_g _21391_ (.A(is_alu_reg_reg), .B(_13840_), .Y(_14773_));
AND_g _21392_ (.A(_13840_), .B(_14764_), .Y(_14774_));
NAND_g _21393_ (.A(_14756_), .B(_14774_), .Y(_14775_));
NAND_g _21394_ (.A(_14772_), .B(_14775_), .Y(_00386_));
NAND_g _21395_ (.A(instr_slt), .B(_14431_), .Y(_14776_));
AND_g _21396_ (.A(_14761_), .B(_14764_), .Y(_14777_));
NAND_g _21397_ (.A(_13844_), .B(_14777_), .Y(_14778_));
NAND_g _21398_ (.A(_14776_), .B(_14778_), .Y(_00387_));
NAND_g _21399_ (.A(instr_sltu), .B(_14431_), .Y(_14779_));
NAND_g _21400_ (.A(_14738_), .B(_14777_), .Y(_14780_));
NAND_g _21401_ (.A(_14779_), .B(_14780_), .Y(_00388_));
NAND_g _21402_ (.A(instr_xor), .B(_14431_), .Y(_14781_));
NAND_g _21403_ (.A(_14441_), .B(_14777_), .Y(_14782_));
NAND_g _21404_ (.A(_14781_), .B(_14782_), .Y(_00389_));
NAND_g _21405_ (.A(instr_srl), .B(_14431_), .Y(_14783_));
AND_g _21406_ (.A(_14444_), .B(_14764_), .Y(_14784_));
NAND_g _21407_ (.A(_14761_), .B(_14784_), .Y(_14785_));
NAND_g _21408_ (.A(_14783_), .B(_14785_), .Y(_00390_));
NAND_g _21409_ (.A(instr_sra), .B(_14431_), .Y(_14786_));
NAND_g _21410_ (.A(_14770_), .B(_14784_), .Y(_14787_));
NAND_g _21411_ (.A(_14786_), .B(_14787_), .Y(_00391_));
NAND_g _21412_ (.A(instr_or), .B(_14431_), .Y(_14788_));
NAND_g _21413_ (.A(_14447_), .B(_14777_), .Y(_14789_));
NAND_g _21414_ (.A(_14788_), .B(_14789_), .Y(_00392_));
NAND_g _21415_ (.A(instr_and), .B(_14431_), .Y(_14790_));
NAND_g _21416_ (.A(_14451_), .B(_14777_), .Y(_14791_));
NAND_g _21417_ (.A(_14790_), .B(_14791_), .Y(_00393_));
NAND_g _21418_ (.A(instr_srai), .B(_13841_), .Y(_14792_));
NAND_g _21419_ (.A(_14760_), .B(_14770_), .Y(_14793_));
NAND_g _21420_ (.A(_14792_), .B(_14793_), .Y(_00394_));
NAND_g _21421_ (.A(instr_rdcycle), .B(_13841_), .Y(_14794_));
NOR_g _21422_ (.A(mem_rdata_q[24]), .B(_13841_), .Y(_14795_));
NAND_g _21423_ (.A(_14750_), .B(_14795_), .Y(_14796_));
NOR_g _21424_ (.A(mem_rdata_q[27]), .B(_14796_), .Y(_14797_));
NOR_g _21425_ (.A(mem_rdata_q[15]), .B(mem_rdata_q[16]), .Y(_14798_));
NOR_g _21426_ (.A(mem_rdata_q[17]), .B(mem_rdata_q[18]), .Y(_14799_));
AND_g _21427_ (.A(_14798_), .B(_14799_), .Y(_14800_));
AND_g _21428_ (.A(_14768_), .B(_14800_), .Y(_14801_));
AND_g _21429_ (.A(mem_rdata_q[31]), .B(mem_rdata_q[0]), .Y(_14802_));
AND_g _21430_ (.A(mem_rdata_q[1]), .B(_08874_), .Y(_14803_));
AND_g _21431_ (.A(_14802_), .B(_14803_), .Y(_14804_));
NOR_g _21432_ (.A(mem_rdata_q[19]), .B(mem_rdata_q[22]), .Y(_14805_));
NOR_g _21433_ (.A(mem_rdata_q[23]), .B(mem_rdata_q[28]), .Y(_14806_));
AND_g _21434_ (.A(_14805_), .B(_14806_), .Y(_14807_));
AND_g _21435_ (.A(_14804_), .B(_14807_), .Y(_14808_));
AND_g _21436_ (.A(_08875_), .B(mem_rdata_q[4]), .Y(_14809_));
AND_g _21437_ (.A(mem_rdata_q[5]), .B(mem_rdata_q[6]), .Y(_14810_));
AND_g _21438_ (.A(_14809_), .B(_14810_), .Y(_14811_));
AND_g _21439_ (.A(_13844_), .B(_14811_), .Y(_14812_));
AND_g _21440_ (.A(_14808_), .B(_14812_), .Y(_14813_));
NAND_g _21441_ (.A(_14801_), .B(_14813_), .Y(_14814_));
NOR_g _21442_ (.A(mem_rdata_q[21]), .B(_14814_), .Y(_14815_));
NAND_g _21443_ (.A(_14797_), .B(_14815_), .Y(_14816_));
NAND_g _21444_ (.A(_14794_), .B(_14816_), .Y(_00395_));
NAND_g _21445_ (.A(instr_rdcycleh), .B(_13841_), .Y(_14817_));
NOR_g _21446_ (.A(_08869_), .B(_14796_), .Y(_14818_));
NAND_g _21447_ (.A(_14815_), .B(_14818_), .Y(_14819_));
NAND_g _21448_ (.A(_14817_), .B(_14819_), .Y(_00396_));
NAND_g _21449_ (.A(instr_rdinstr), .B(_13841_), .Y(_14820_));
NAND_g _21450_ (.A(_08868_), .B(mem_rdata_q[21]), .Y(_14821_));
NOR_g _21451_ (.A(_14814_), .B(_14821_), .Y(_14822_));
NAND_g _21452_ (.A(_14797_), .B(_14822_), .Y(_14823_));
NAND_g _21453_ (.A(_14820_), .B(_14823_), .Y(_00397_));
NAND_g _21454_ (.A(instr_rdinstrh), .B(_13841_), .Y(_14824_));
NAND_g _21455_ (.A(_14818_), .B(_14822_), .Y(_14825_));
NAND_g _21456_ (.A(_14824_), .B(_14825_), .Y(_00398_));
NAND_g _21457_ (.A(mem_rdata[7]), .B(_09903_), .Y(_14826_));
NAND_g _21458_ (.A(mem_rdata_q[7]), .B(_09904_), .Y(_14827_));
NAND_g _21459_ (.A(_14826_), .B(_14827_), .Y(_00421_));
NAND_g _21460_ (.A(_14393_), .B(_00421_), .Y(_14828_));
NAND_g _21461_ (.A(decoded_rd[0]), .B(_14394_), .Y(_14829_));
NAND_g _21462_ (.A(_14828_), .B(_14829_), .Y(_00399_));
NAND_g _21463_ (.A(mem_rdata[8]), .B(_09903_), .Y(_14830_));
NAND_g _21464_ (.A(mem_rdata_q[8]), .B(_09904_), .Y(_14831_));
NAND_g _21465_ (.A(_14830_), .B(_14831_), .Y(_00422_));
NAND_g _21466_ (.A(_14393_), .B(_00422_), .Y(_14832_));
NAND_g _21467_ (.A(decoded_rd[1]), .B(_14394_), .Y(_14833_));
NAND_g _21468_ (.A(_14832_), .B(_14833_), .Y(_00400_));
NAND_g _21469_ (.A(mem_rdata[9]), .B(_09903_), .Y(_14834_));
NAND_g _21470_ (.A(mem_rdata_q[9]), .B(_09904_), .Y(_14835_));
NAND_g _21471_ (.A(_14834_), .B(_14835_), .Y(_00423_));
NAND_g _21472_ (.A(_14393_), .B(_00423_), .Y(_14836_));
NAND_g _21473_ (.A(decoded_rd[2]), .B(_14394_), .Y(_14837_));
NAND_g _21474_ (.A(_14836_), .B(_14837_), .Y(_00401_));
NAND_g _21475_ (.A(mem_rdata[10]), .B(_09903_), .Y(_14838_));
NAND_g _21476_ (.A(mem_rdata_q[10]), .B(_09904_), .Y(_14839_));
NAND_g _21477_ (.A(_14838_), .B(_14839_), .Y(_00424_));
NAND_g _21478_ (.A(_14393_), .B(_00424_), .Y(_14840_));
NAND_g _21479_ (.A(decoded_rd[3]), .B(_14394_), .Y(_14841_));
NAND_g _21480_ (.A(_14840_), .B(_14841_), .Y(_00402_));
NAND_g _21481_ (.A(mem_rdata[11]), .B(_09903_), .Y(_14842_));
NAND_g _21482_ (.A(mem_rdata_q[11]), .B(_09904_), .Y(_14843_));
NAND_g _21483_ (.A(_14842_), .B(_14843_), .Y(_00425_));
NAND_g _21484_ (.A(_14393_), .B(_00425_), .Y(_14844_));
NAND_g _21485_ (.A(decoded_rd[4]), .B(_14394_), .Y(_14845_));
NAND_g _21486_ (.A(_14844_), .B(_14845_), .Y(_00403_));
NAND_g _21487_ (.A(mem_rdata[20]), .B(_09903_), .Y(_14846_));
NAND_g _21488_ (.A(mem_rdata_q[20]), .B(_09904_), .Y(_14847_));
NAND_g _21489_ (.A(_14846_), .B(_14847_), .Y(_00434_));
NAND_g _21490_ (.A(_14393_), .B(_00434_), .Y(_14848_));
NAND_g _21491_ (.A(decoded_imm_j[11]), .B(_14394_), .Y(_14849_));
NAND_g _21492_ (.A(_14848_), .B(_14849_), .Y(_00404_));
NAND_g _21493_ (.A(mem_rdata[21]), .B(_09903_), .Y(_14850_));
NAND_g _21494_ (.A(mem_rdata_q[21]), .B(_09904_), .Y(_14851_));
NAND_g _21495_ (.A(_14850_), .B(_14851_), .Y(_00435_));
NAND_g _21496_ (.A(_14393_), .B(_00435_), .Y(_14852_));
NAND_g _21497_ (.A(decoded_imm_j[1]), .B(_14394_), .Y(_14853_));
NAND_g _21498_ (.A(_14852_), .B(_14853_), .Y(_00405_));
NAND_g _21499_ (.A(mem_rdata[22]), .B(_09903_), .Y(_14854_));
NAND_g _21500_ (.A(mem_rdata_q[22]), .B(_09904_), .Y(_14855_));
NAND_g _21501_ (.A(_14854_), .B(_14855_), .Y(_00436_));
NAND_g _21502_ (.A(_14393_), .B(_00436_), .Y(_14856_));
NAND_g _21503_ (.A(decoded_imm_j[2]), .B(_14394_), .Y(_14857_));
NAND_g _21504_ (.A(_14856_), .B(_14857_), .Y(_00406_));
NAND_g _21505_ (.A(mem_rdata[23]), .B(_09903_), .Y(_14858_));
NAND_g _21506_ (.A(mem_rdata_q[23]), .B(_09904_), .Y(_14859_));
NAND_g _21507_ (.A(_14858_), .B(_14859_), .Y(_00437_));
NAND_g _21508_ (.A(_14393_), .B(_00437_), .Y(_14860_));
NAND_g _21509_ (.A(decoded_imm_j[3]), .B(_14394_), .Y(_14861_));
NAND_g _21510_ (.A(_14860_), .B(_14861_), .Y(_00407_));
NAND_g _21511_ (.A(mem_rdata_q[7]), .B(_13845_), .Y(_14862_));
NOR_g _21512_ (.A(instr_jalr), .B(is_lb_lh_lw_lbu_lhu), .Y(_14863_));
NAND_g _21513_ (.A(_08863_), .B(_14863_), .Y(_14864_));
NOT_g _21514_ (.A(_14864_), .Y(_14865_));
AND_g _21515_ (.A(mem_rdata_q[20]), .B(_13840_), .Y(_14866_));
NAND_g _21516_ (.A(_14864_), .B(_14866_), .Y(_14867_));
NAND_g _21517_ (.A(decoded_imm[0]), .B(_13841_), .Y(_14868_));
AND_g _21518_ (.A(_14862_), .B(_14867_), .Y(_14869_));
NAND_g _21519_ (.A(_14868_), .B(_14869_), .Y(_00408_));
NAND_g _21520_ (.A(mem_rdata[30]), .B(_09903_), .Y(_14870_));
NAND_g _21521_ (.A(mem_rdata_q[30]), .B(_09904_), .Y(_14871_));
NAND_g _21522_ (.A(_14870_), .B(_14871_), .Y(_00444_));
NAND_g _21523_ (.A(_14393_), .B(_00444_), .Y(_14872_));
NAND_g _21524_ (.A(decoded_imm_j[10]), .B(_14394_), .Y(_14873_));
NAND_g _21525_ (.A(_14872_), .B(_14873_), .Y(_00409_));
NOR_g _21526_ (.A(_00516_), .B(_00517_), .Y(_14874_));
AND_g _21527_ (.A(_14399_), .B(_14874_), .Y(_14875_));
AND_g _21528_ (.A(_14409_), .B(_14412_), .Y(_14876_));
AND_g _21529_ (.A(_14875_), .B(_14876_), .Y(_14877_));
AND_g _21530_ (.A(_14416_), .B(_14877_), .Y(_14878_));
NAND_g _21531_ (.A(is_lb_lh_lw_lbu_lhu), .B(_14394_), .Y(_14879_));
NAND_g _21532_ (.A(_14393_), .B(_14878_), .Y(_14880_));
NAND_g _21533_ (.A(_14879_), .B(_14880_), .Y(_00410_));
NAND_g _21534_ (.A(is_slli_srli_srai), .B(_13841_), .Y(_14881_));
NAND_g _21535_ (.A(_14444_), .B(_14754_), .Y(_14882_));
NAND_g _21536_ (.A(_14757_), .B(_14882_), .Y(_14883_));
NAND_g _21537_ (.A(_14733_), .B(_14883_), .Y(_14884_));
NAND_g _21538_ (.A(_14881_), .B(_14884_), .Y(_00411_));
NAND_g _21539_ (.A(is_alu_reg_imm), .B(_14437_), .Y(_14885_));
NOR_g _21540_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi), .B(_13840_), .Y(_14886_));
NOR_g _21541_ (.A(instr_jalr), .B(_13841_), .Y(_14887_));
AND_g _21542_ (.A(_14885_), .B(_14887_), .Y(_14888_));
NOR_g _21543_ (.A(_14886_), .B(_14888_), .Y(_00412_));
NAND_g _21544_ (.A(is_sll_srl_sra), .B(_13841_), .Y(_14889_));
NAND_g _21545_ (.A(_14773_), .B(_14883_), .Y(_14890_));
NAND_g _21546_ (.A(_14889_), .B(_14890_), .Y(_00413_));
NAND_g _21547_ (.A(_13900_), .B(_14394_), .Y(_14891_));
AND_g _21548_ (.A(_14426_), .B(_14875_), .Y(_14892_));
NAND_g _21549_ (.A(_14393_), .B(_14892_), .Y(_14893_));
NAND_g _21550_ (.A(_14891_), .B(_14893_), .Y(_00414_));
AND_g _21551_ (.A(_08796_), .B(_10725_), .Y(_14894_));
NAND_g _21552_ (.A(_10739_), .B(_14894_), .Y(_14895_));
AND_g _21553_ (.A(_13841_), .B(_14895_), .Y(_00415_));
NAND_g _21554_ (.A(_14421_), .B(_14875_), .Y(_14896_));
NAND_g _21555_ (.A(_14393_), .B(_14896_), .Y(_14897_));
NAND_g _21556_ (.A(_08863_), .B(_14394_), .Y(_14898_));
AND_g _21557_ (.A(_14897_), .B(_14898_), .Y(_00416_));
NAND_g _21558_ (.A(_14417_), .B(_14875_), .Y(_14899_));
AND_g _21559_ (.A(_14393_), .B(_14899_), .Y(_14900_));
NOR_g _21560_ (.A(is_alu_reg_reg), .B(_14393_), .Y(_14901_));
NOR_g _21561_ (.A(_14900_), .B(_14901_), .Y(_00417_));
AND_g _21562_ (.A(_00519_), .B(_14877_), .Y(_14902_));
NAND_g _21563_ (.A(is_sb_sh_sw), .B(_14394_), .Y(_14903_));
NAND_g _21564_ (.A(_14393_), .B(_14902_), .Y(_14904_));
NAND_g _21565_ (.A(_14903_), .B(_14904_), .Y(_00418_));
NAND_g _21566_ (.A(_08790_), .B(_10719_), .Y(_14905_));
AND_g _21567_ (.A(_14431_), .B(_14905_), .Y(_00419_));
NAND_g _21568_ (.A(mem_instr), .B(_14271_), .Y(_14906_));
NAND_g _21569_ (.A(_14263_), .B(_14281_), .Y(_14907_));
NAND_g _21570_ (.A(_14906_), .B(_14907_), .Y(_00420_));
NAND_g _21571_ (.A(mem_rdata[15]), .B(_09903_), .Y(_14908_));
NAND_g _21572_ (.A(mem_rdata_q[15]), .B(_09904_), .Y(_14909_));
NAND_g _21573_ (.A(_14908_), .B(_14909_), .Y(_00429_));
NAND_g _21574_ (.A(mem_rdata[16]), .B(_09903_), .Y(_14910_));
NAND_g _21575_ (.A(mem_rdata_q[16]), .B(_09904_), .Y(_14911_));
NAND_g _21576_ (.A(_14910_), .B(_14911_), .Y(_00430_));
NAND_g _21577_ (.A(mem_rdata[17]), .B(_09903_), .Y(_14912_));
NAND_g _21578_ (.A(mem_rdata_q[17]), .B(_09904_), .Y(_14913_));
NAND_g _21579_ (.A(_14912_), .B(_14913_), .Y(_00431_));
NAND_g _21580_ (.A(mem_rdata[18]), .B(_09903_), .Y(_14914_));
NAND_g _21581_ (.A(mem_rdata_q[18]), .B(_09904_), .Y(_14915_));
NAND_g _21582_ (.A(_14914_), .B(_14915_), .Y(_00432_));
NAND_g _21583_ (.A(mem_rdata[19]), .B(_09903_), .Y(_14916_));
NAND_g _21584_ (.A(mem_rdata_q[19]), .B(_09904_), .Y(_14917_));
NAND_g _21585_ (.A(_14916_), .B(_14917_), .Y(_00433_));
NAND_g _21586_ (.A(mem_rdata[24]), .B(_09903_), .Y(_14918_));
NAND_g _21587_ (.A(mem_rdata_q[24]), .B(_09904_), .Y(_14919_));
NAND_g _21588_ (.A(_14918_), .B(_14919_), .Y(_00438_));
NAND_g _21589_ (.A(mem_rdata[25]), .B(_09903_), .Y(_14920_));
NAND_g _21590_ (.A(mem_rdata_q[25]), .B(_09904_), .Y(_14921_));
NAND_g _21591_ (.A(_14920_), .B(_14921_), .Y(_00439_));
NAND_g _21592_ (.A(mem_rdata[26]), .B(_09903_), .Y(_14922_));
NAND_g _21593_ (.A(mem_rdata_q[26]), .B(_09904_), .Y(_14923_));
NAND_g _21594_ (.A(_14922_), .B(_14923_), .Y(_00440_));
NAND_g _21595_ (.A(mem_rdata[27]), .B(_09903_), .Y(_14924_));
NAND_g _21596_ (.A(mem_rdata_q[27]), .B(_09904_), .Y(_14925_));
NAND_g _21597_ (.A(_14924_), .B(_14925_), .Y(_00441_));
NAND_g _21598_ (.A(mem_rdata[28]), .B(_09903_), .Y(_14926_));
NAND_g _21599_ (.A(mem_rdata_q[28]), .B(_09904_), .Y(_14927_));
NAND_g _21600_ (.A(_14926_), .B(_14927_), .Y(_00442_));
NAND_g _21601_ (.A(mem_rdata[29]), .B(_09903_), .Y(_14928_));
NAND_g _21602_ (.A(mem_rdata_q[29]), .B(_09904_), .Y(_14929_));
NAND_g _21603_ (.A(_14928_), .B(_14929_), .Y(_00443_));
NAND_g _21604_ (.A(mem_rdata[31]), .B(_09903_), .Y(_14930_));
NAND_g _21605_ (.A(mem_rdata_q[31]), .B(_09904_), .Y(_14931_));
NAND_g _21606_ (.A(_14930_), .B(_14931_), .Y(_00445_));
NAND_g _21607_ (.A(reg_out[2]), .B(_09913_), .Y(_14932_));
NAND_g _21608_ (.A(_09922_), .B(_14932_), .Y(_14933_));
NAND_g _21609_ (.A(_14263_), .B(_14933_), .Y(_14934_));
NAND_g _21610_ (.A(pcpi_rs1[2]), .B(_14262_), .Y(_14935_));
NAND_g _21611_ (.A(_14934_), .B(_14935_), .Y(mem_la_addr[2]));
NAND_g _21612_ (.A(_14270_), .B(mem_la_addr[2]), .Y(_14936_));
NAND_g _21613_ (.A(mem_addr[2]), .B(_14271_), .Y(_14937_));
NAND_g _21614_ (.A(_14936_), .B(_14937_), .Y(_00446_));
NAND_g _21615_ (.A(reg_out[3]), .B(_09913_), .Y(_14938_));
NAND_g _21616_ (.A(_09928_), .B(_14938_), .Y(_14939_));
NAND_g _21617_ (.A(_14263_), .B(_14939_), .Y(_14940_));
NAND_g _21618_ (.A(pcpi_rs1[3]), .B(_14262_), .Y(_14941_));
NAND_g _21619_ (.A(_14940_), .B(_14941_), .Y(mem_la_addr[3]));
NAND_g _21620_ (.A(_14270_), .B(mem_la_addr[3]), .Y(_14942_));
NAND_g _21621_ (.A(mem_addr[3]), .B(_14271_), .Y(_14943_));
NAND_g _21622_ (.A(_14942_), .B(_14943_), .Y(_00447_));
NAND_g _21623_ (.A(reg_out[4]), .B(_09913_), .Y(_14944_));
NAND_g _21624_ (.A(_09934_), .B(_14944_), .Y(_14945_));
NAND_g _21625_ (.A(_14263_), .B(_14945_), .Y(_14946_));
NAND_g _21626_ (.A(pcpi_rs1[4]), .B(_14262_), .Y(_14947_));
NAND_g _21627_ (.A(_14946_), .B(_14947_), .Y(mem_la_addr[4]));
NAND_g _21628_ (.A(_14270_), .B(mem_la_addr[4]), .Y(_14948_));
NAND_g _21629_ (.A(mem_addr[4]), .B(_14271_), .Y(_14949_));
NAND_g _21630_ (.A(_14948_), .B(_14949_), .Y(_00448_));
NAND_g _21631_ (.A(reg_out[5]), .B(_09913_), .Y(_14950_));
NAND_g _21632_ (.A(_09940_), .B(_14950_), .Y(_14951_));
NAND_g _21633_ (.A(_14263_), .B(_14951_), .Y(_14952_));
NAND_g _21634_ (.A(pcpi_rs1[5]), .B(_14262_), .Y(_14953_));
NAND_g _21635_ (.A(_14952_), .B(_14953_), .Y(mem_la_addr[5]));
NAND_g _21636_ (.A(_14270_), .B(mem_la_addr[5]), .Y(_14954_));
NAND_g _21637_ (.A(mem_addr[5]), .B(_14271_), .Y(_14955_));
NAND_g _21638_ (.A(_14954_), .B(_14955_), .Y(_00449_));
NAND_g _21639_ (.A(reg_out[6]), .B(_09913_), .Y(_14956_));
NAND_g _21640_ (.A(_09946_), .B(_14956_), .Y(_14957_));
NAND_g _21641_ (.A(_14263_), .B(_14957_), .Y(_14958_));
NAND_g _21642_ (.A(pcpi_rs1[6]), .B(_14262_), .Y(_14959_));
NAND_g _21643_ (.A(_14958_), .B(_14959_), .Y(mem_la_addr[6]));
NAND_g _21644_ (.A(_14270_), .B(mem_la_addr[6]), .Y(_14960_));
NAND_g _21645_ (.A(mem_addr[6]), .B(_14271_), .Y(_14961_));
NAND_g _21646_ (.A(_14960_), .B(_14961_), .Y(_00450_));
NAND_g _21647_ (.A(reg_out[7]), .B(_09913_), .Y(_14962_));
NAND_g _21648_ (.A(_09952_), .B(_14962_), .Y(_14963_));
NAND_g _21649_ (.A(_14263_), .B(_14963_), .Y(_14964_));
NAND_g _21650_ (.A(pcpi_rs1[7]), .B(_14262_), .Y(_14965_));
NAND_g _21651_ (.A(_14964_), .B(_14965_), .Y(mem_la_addr[7]));
NAND_g _21652_ (.A(mem_addr[7]), .B(_14271_), .Y(_14966_));
NAND_g _21653_ (.A(_14270_), .B(mem_la_addr[7]), .Y(_14967_));
NAND_g _21654_ (.A(_14966_), .B(_14967_), .Y(_00451_));
NAND_g _21655_ (.A(reg_out[8]), .B(_09913_), .Y(_14968_));
NAND_g _21656_ (.A(_09958_), .B(_14968_), .Y(_14969_));
NAND_g _21657_ (.A(_14263_), .B(_14969_), .Y(_14970_));
NAND_g _21658_ (.A(pcpi_rs1[8]), .B(_14262_), .Y(_14971_));
NAND_g _21659_ (.A(_14970_), .B(_14971_), .Y(mem_la_addr[8]));
NAND_g _21660_ (.A(_14270_), .B(mem_la_addr[8]), .Y(_14972_));
NAND_g _21661_ (.A(mem_addr[8]), .B(_14271_), .Y(_14973_));
NAND_g _21662_ (.A(_14972_), .B(_14973_), .Y(_00452_));
NAND_g _21663_ (.A(reg_out[9]), .B(_09913_), .Y(_14974_));
NAND_g _21664_ (.A(_09964_), .B(_14974_), .Y(_14975_));
NAND_g _21665_ (.A(_14263_), .B(_14975_), .Y(_14976_));
NAND_g _21666_ (.A(pcpi_rs1[9]), .B(_14262_), .Y(_14977_));
NAND_g _21667_ (.A(_14976_), .B(_14977_), .Y(mem_la_addr[9]));
NAND_g _21668_ (.A(_14270_), .B(mem_la_addr[9]), .Y(_14978_));
NAND_g _21669_ (.A(mem_addr[9]), .B(_14271_), .Y(_14979_));
NAND_g _21670_ (.A(_14978_), .B(_14979_), .Y(_00453_));
NAND_g _21671_ (.A(reg_out[10]), .B(_09913_), .Y(_14980_));
NAND_g _21672_ (.A(_09970_), .B(_14980_), .Y(_14981_));
NAND_g _21673_ (.A(_14263_), .B(_14981_), .Y(_14982_));
NAND_g _21674_ (.A(pcpi_rs1[10]), .B(_14262_), .Y(_14983_));
NAND_g _21675_ (.A(_14982_), .B(_14983_), .Y(mem_la_addr[10]));
NAND_g _21676_ (.A(_14270_), .B(mem_la_addr[10]), .Y(_14984_));
NAND_g _21677_ (.A(mem_addr[10]), .B(_14271_), .Y(_14985_));
NAND_g _21678_ (.A(_14984_), .B(_14985_), .Y(_00454_));
NAND_g _21679_ (.A(reg_out[11]), .B(_09913_), .Y(_14986_));
NAND_g _21680_ (.A(_09976_), .B(_14986_), .Y(_14987_));
NAND_g _21681_ (.A(_14263_), .B(_14987_), .Y(_14988_));
NAND_g _21682_ (.A(pcpi_rs1[11]), .B(_14262_), .Y(_14989_));
NAND_g _21683_ (.A(_14988_), .B(_14989_), .Y(mem_la_addr[11]));
NAND_g _21684_ (.A(_14270_), .B(mem_la_addr[11]), .Y(_14990_));
NAND_g _21685_ (.A(mem_addr[11]), .B(_14271_), .Y(_14991_));
NAND_g _21686_ (.A(_14990_), .B(_14991_), .Y(_00455_));
NAND_g _21687_ (.A(reg_out[12]), .B(_09913_), .Y(_14992_));
NAND_g _21688_ (.A(_09982_), .B(_14992_), .Y(_14993_));
NAND_g _21689_ (.A(_14263_), .B(_14993_), .Y(_14994_));
NAND_g _21690_ (.A(pcpi_rs1[12]), .B(_14262_), .Y(_14995_));
NAND_g _21691_ (.A(_14994_), .B(_14995_), .Y(mem_la_addr[12]));
NAND_g _21692_ (.A(_14270_), .B(mem_la_addr[12]), .Y(_14996_));
NAND_g _21693_ (.A(mem_addr[12]), .B(_14271_), .Y(_14997_));
NAND_g _21694_ (.A(_14996_), .B(_14997_), .Y(_00456_));
NAND_g _21695_ (.A(reg_out[13]), .B(_09913_), .Y(_14998_));
NAND_g _21696_ (.A(_09988_), .B(_14998_), .Y(_01535_));
NAND_g _21697_ (.A(_14263_), .B(_01535_), .Y(_01536_));
NAND_g _21698_ (.A(pcpi_rs1[13]), .B(_14262_), .Y(_01537_));
NAND_g _21699_ (.A(_01536_), .B(_01537_), .Y(mem_la_addr[13]));
NAND_g _21700_ (.A(_14270_), .B(mem_la_addr[13]), .Y(_01538_));
NAND_g _21701_ (.A(mem_addr[13]), .B(_14271_), .Y(_01539_));
NAND_g _21702_ (.A(_01538_), .B(_01539_), .Y(_00457_));
NAND_g _21703_ (.A(reg_out[14]), .B(_09913_), .Y(_01540_));
NAND_g _21704_ (.A(_09994_), .B(_01540_), .Y(_01541_));
NAND_g _21705_ (.A(_14263_), .B(_01541_), .Y(_01542_));
NAND_g _21706_ (.A(pcpi_rs1[14]), .B(_14262_), .Y(_01543_));
NAND_g _21707_ (.A(_01542_), .B(_01543_), .Y(mem_la_addr[14]));
NAND_g _21708_ (.A(_14270_), .B(mem_la_addr[14]), .Y(_01544_));
NAND_g _21709_ (.A(mem_addr[14]), .B(_14271_), .Y(_01545_));
NAND_g _21710_ (.A(_01544_), .B(_01545_), .Y(_00458_));
NAND_g _21711_ (.A(reg_out[15]), .B(_09913_), .Y(_01546_));
NAND_g _21712_ (.A(_10000_), .B(_01546_), .Y(_01547_));
NAND_g _21713_ (.A(_14263_), .B(_01547_), .Y(_01548_));
NAND_g _21714_ (.A(pcpi_rs1[15]), .B(_14262_), .Y(_01549_));
NAND_g _21715_ (.A(_01548_), .B(_01549_), .Y(mem_la_addr[15]));
NAND_g _21716_ (.A(_14270_), .B(mem_la_addr[15]), .Y(_01550_));
NAND_g _21717_ (.A(mem_addr[15]), .B(_14271_), .Y(_01551_));
NAND_g _21718_ (.A(_01550_), .B(_01551_), .Y(_00459_));
NAND_g _21719_ (.A(reg_out[16]), .B(_09913_), .Y(_01552_));
NAND_g _21720_ (.A(_10006_), .B(_01552_), .Y(_01553_));
NAND_g _21721_ (.A(_14263_), .B(_01553_), .Y(_01554_));
NAND_g _21722_ (.A(pcpi_rs1[16]), .B(_14262_), .Y(_01555_));
NAND_g _21723_ (.A(_01554_), .B(_01555_), .Y(mem_la_addr[16]));
NAND_g _21724_ (.A(_14270_), .B(mem_la_addr[16]), .Y(_01556_));
NAND_g _21725_ (.A(mem_addr[16]), .B(_14271_), .Y(_01557_));
NAND_g _21726_ (.A(_01556_), .B(_01557_), .Y(_00460_));
NAND_g _21727_ (.A(reg_out[17]), .B(_09913_), .Y(_01558_));
NAND_g _21728_ (.A(_10012_), .B(_01558_), .Y(_01559_));
NAND_g _21729_ (.A(_14263_), .B(_01559_), .Y(_01560_));
NAND_g _21730_ (.A(pcpi_rs1[17]), .B(_14262_), .Y(_01561_));
NAND_g _21731_ (.A(_01560_), .B(_01561_), .Y(mem_la_addr[17]));
NAND_g _21732_ (.A(_14270_), .B(mem_la_addr[17]), .Y(_01562_));
NAND_g _21733_ (.A(mem_addr[17]), .B(_14271_), .Y(_01563_));
NAND_g _21734_ (.A(_01562_), .B(_01563_), .Y(_00461_));
NAND_g _21735_ (.A(reg_out[18]), .B(_09913_), .Y(_01564_));
NAND_g _21736_ (.A(_10018_), .B(_01564_), .Y(_01565_));
NAND_g _21737_ (.A(_14263_), .B(_01565_), .Y(_01566_));
NAND_g _21738_ (.A(pcpi_rs1[18]), .B(_14262_), .Y(_01567_));
NAND_g _21739_ (.A(_01566_), .B(_01567_), .Y(mem_la_addr[18]));
NAND_g _21740_ (.A(_14270_), .B(mem_la_addr[18]), .Y(_01568_));
NAND_g _21741_ (.A(mem_addr[18]), .B(_14271_), .Y(_01569_));
NAND_g _21742_ (.A(_01568_), .B(_01569_), .Y(_00462_));
NAND_g _21743_ (.A(reg_out[19]), .B(_09913_), .Y(_01570_));
NAND_g _21744_ (.A(_10024_), .B(_01570_), .Y(_01571_));
NAND_g _21745_ (.A(_14263_), .B(_01571_), .Y(_01572_));
NAND_g _21746_ (.A(pcpi_rs1[19]), .B(_14262_), .Y(_01573_));
NAND_g _21747_ (.A(_01572_), .B(_01573_), .Y(mem_la_addr[19]));
NAND_g _21748_ (.A(mem_addr[19]), .B(_14271_), .Y(_01574_));
NAND_g _21749_ (.A(_14270_), .B(mem_la_addr[19]), .Y(_01575_));
NAND_g _21750_ (.A(_01574_), .B(_01575_), .Y(_00463_));
NAND_g _21751_ (.A(reg_out[20]), .B(_09913_), .Y(_01576_));
NAND_g _21752_ (.A(_10030_), .B(_01576_), .Y(_01577_));
NAND_g _21753_ (.A(_14263_), .B(_01577_), .Y(_01578_));
NAND_g _21754_ (.A(pcpi_rs1[20]), .B(_14262_), .Y(_01579_));
NAND_g _21755_ (.A(_01578_), .B(_01579_), .Y(mem_la_addr[20]));
NAND_g _21756_ (.A(_14270_), .B(mem_la_addr[20]), .Y(_01580_));
NAND_g _21757_ (.A(mem_addr[20]), .B(_14271_), .Y(_01581_));
NAND_g _21758_ (.A(_01580_), .B(_01581_), .Y(_00464_));
NAND_g _21759_ (.A(reg_out[21]), .B(_09913_), .Y(_01582_));
NAND_g _21760_ (.A(_10036_), .B(_01582_), .Y(_01583_));
NAND_g _21761_ (.A(_14263_), .B(_01583_), .Y(_01584_));
NAND_g _21762_ (.A(pcpi_rs1[21]), .B(_14262_), .Y(_01585_));
NAND_g _21763_ (.A(_01584_), .B(_01585_), .Y(mem_la_addr[21]));
NAND_g _21764_ (.A(_14270_), .B(mem_la_addr[21]), .Y(_01586_));
NAND_g _21765_ (.A(mem_addr[21]), .B(_14271_), .Y(_01587_));
NAND_g _21766_ (.A(_01586_), .B(_01587_), .Y(_00465_));
NAND_g _21767_ (.A(reg_out[22]), .B(_09913_), .Y(_01588_));
NAND_g _21768_ (.A(_10042_), .B(_01588_), .Y(_01589_));
NAND_g _21769_ (.A(_14263_), .B(_01589_), .Y(_01590_));
NAND_g _21770_ (.A(pcpi_rs1[22]), .B(_14262_), .Y(_01591_));
NAND_g _21771_ (.A(_01590_), .B(_01591_), .Y(mem_la_addr[22]));
NAND_g _21772_ (.A(_14270_), .B(mem_la_addr[22]), .Y(_01592_));
NAND_g _21773_ (.A(mem_addr[22]), .B(_14271_), .Y(_01593_));
NAND_g _21774_ (.A(_01592_), .B(_01593_), .Y(_00466_));
NAND_g _21775_ (.A(reg_out[23]), .B(_09913_), .Y(_01594_));
NAND_g _21776_ (.A(_10048_), .B(_01594_), .Y(_01595_));
NAND_g _21777_ (.A(_14263_), .B(_01595_), .Y(_01596_));
NAND_g _21778_ (.A(pcpi_rs1[23]), .B(_14262_), .Y(_01597_));
NAND_g _21779_ (.A(_01596_), .B(_01597_), .Y(mem_la_addr[23]));
NAND_g _21780_ (.A(_14270_), .B(mem_la_addr[23]), .Y(_01598_));
NAND_g _21781_ (.A(mem_addr[23]), .B(_14271_), .Y(_01599_));
NAND_g _21782_ (.A(_01598_), .B(_01599_), .Y(_00467_));
NAND_g _21783_ (.A(reg_out[24]), .B(_09913_), .Y(_01600_));
NAND_g _21784_ (.A(_10054_), .B(_01600_), .Y(_01601_));
NAND_g _21785_ (.A(_14263_), .B(_01601_), .Y(_01602_));
NAND_g _21786_ (.A(pcpi_rs1[24]), .B(_14262_), .Y(_01603_));
NAND_g _21787_ (.A(_01602_), .B(_01603_), .Y(mem_la_addr[24]));
NAND_g _21788_ (.A(mem_addr[24]), .B(_14271_), .Y(_01604_));
NAND_g _21789_ (.A(_14270_), .B(mem_la_addr[24]), .Y(_01605_));
NAND_g _21790_ (.A(_01604_), .B(_01605_), .Y(_00468_));
NAND_g _21791_ (.A(reg_out[25]), .B(_09913_), .Y(_01606_));
NAND_g _21792_ (.A(_10060_), .B(_01606_), .Y(_01607_));
NAND_g _21793_ (.A(_14263_), .B(_01607_), .Y(_01608_));
NAND_g _21794_ (.A(pcpi_rs1[25]), .B(_14262_), .Y(_01609_));
NAND_g _21795_ (.A(_01608_), .B(_01609_), .Y(mem_la_addr[25]));
NAND_g _21796_ (.A(_14270_), .B(mem_la_addr[25]), .Y(_01610_));
NAND_g _21797_ (.A(mem_addr[25]), .B(_14271_), .Y(_01611_));
NAND_g _21798_ (.A(_01610_), .B(_01611_), .Y(_00469_));
NAND_g _21799_ (.A(reg_out[26]), .B(_09913_), .Y(_01612_));
NAND_g _21800_ (.A(_10065_), .B(_01612_), .Y(_01613_));
NAND_g _21801_ (.A(_14263_), .B(_01613_), .Y(_01614_));
NAND_g _21802_ (.A(pcpi_rs1[26]), .B(_14262_), .Y(_01615_));
NAND_g _21803_ (.A(_01614_), .B(_01615_), .Y(mem_la_addr[26]));
NAND_g _21804_ (.A(_14270_), .B(mem_la_addr[26]), .Y(_01616_));
NAND_g _21805_ (.A(mem_addr[26]), .B(_14271_), .Y(_01617_));
NAND_g _21806_ (.A(_01616_), .B(_01617_), .Y(_00470_));
NAND_g _21807_ (.A(reg_out[27]), .B(_09913_), .Y(_01618_));
NAND_g _21808_ (.A(_10071_), .B(_01618_), .Y(_01619_));
NAND_g _21809_ (.A(_14263_), .B(_01619_), .Y(_01620_));
NAND_g _21810_ (.A(pcpi_rs1[27]), .B(_14262_), .Y(_01621_));
NAND_g _21811_ (.A(_01620_), .B(_01621_), .Y(mem_la_addr[27]));
NAND_g _21812_ (.A(_14270_), .B(mem_la_addr[27]), .Y(_01622_));
NAND_g _21813_ (.A(mem_addr[27]), .B(_14271_), .Y(_01623_));
NAND_g _21814_ (.A(_01622_), .B(_01623_), .Y(_00471_));
NAND_g _21815_ (.A(reg_out[28]), .B(_09913_), .Y(_01624_));
NAND_g _21816_ (.A(_10076_), .B(_01624_), .Y(_01625_));
NAND_g _21817_ (.A(_14263_), .B(_01625_), .Y(_01626_));
NAND_g _21818_ (.A(pcpi_rs1[28]), .B(_14262_), .Y(_01627_));
NAND_g _21819_ (.A(_01626_), .B(_01627_), .Y(mem_la_addr[28]));
NAND_g _21820_ (.A(_14270_), .B(mem_la_addr[28]), .Y(_01628_));
NAND_g _21821_ (.A(mem_addr[28]), .B(_14271_), .Y(_01629_));
NAND_g _21822_ (.A(_01628_), .B(_01629_), .Y(_00472_));
NAND_g _21823_ (.A(reg_out[29]), .B(_09913_), .Y(_01630_));
NAND_g _21824_ (.A(_10082_), .B(_01630_), .Y(_01631_));
NAND_g _21825_ (.A(_14263_), .B(_01631_), .Y(_01632_));
NAND_g _21826_ (.A(pcpi_rs1[29]), .B(_14262_), .Y(_01633_));
NAND_g _21827_ (.A(_01632_), .B(_01633_), .Y(mem_la_addr[29]));
NAND_g _21828_ (.A(_14270_), .B(mem_la_addr[29]), .Y(_01634_));
NAND_g _21829_ (.A(mem_addr[29]), .B(_14271_), .Y(_01635_));
NAND_g _21830_ (.A(_01634_), .B(_01635_), .Y(_00473_));
NAND_g _21831_ (.A(reg_out[30]), .B(_09913_), .Y(_01636_));
NAND_g _21832_ (.A(_10088_), .B(_01636_), .Y(_01637_));
NAND_g _21833_ (.A(_14263_), .B(_01637_), .Y(_01638_));
NAND_g _21834_ (.A(pcpi_rs1[30]), .B(_14262_), .Y(_01639_));
NAND_g _21835_ (.A(_01638_), .B(_01639_), .Y(mem_la_addr[30]));
NAND_g _21836_ (.A(_14270_), .B(mem_la_addr[30]), .Y(_01640_));
NAND_g _21837_ (.A(mem_addr[30]), .B(_14271_), .Y(_01641_));
NAND_g _21838_ (.A(_01640_), .B(_01641_), .Y(_00474_));
NAND_g _21839_ (.A(reg_out[31]), .B(_09913_), .Y(_01642_));
NAND_g _21840_ (.A(_10093_), .B(_01642_), .Y(_01643_));
NAND_g _21841_ (.A(_14263_), .B(_01643_), .Y(_01644_));
NAND_g _21842_ (.A(pcpi_rs1[31]), .B(_14262_), .Y(_01645_));
NAND_g _21843_ (.A(_01644_), .B(_01645_), .Y(mem_la_addr[31]));
NAND_g _21844_ (.A(_14270_), .B(mem_la_addr[31]), .Y(_01646_));
NAND_g _21845_ (.A(mem_addr[31]), .B(_14271_), .Y(_01647_));
NAND_g _21846_ (.A(_01646_), .B(_01647_), .Y(_00475_));
NAND_g _21847_ (.A(mem_wordsize[0]), .B(mem_wordsize[1]), .Y(_01648_));
AND_g _21848_ (.A(pcpi_rs2[0]), .B(_01648_), .Y(mem_la_wdata[0]));
AND_g _21849_ (.A(_14260_), .B(_14268_), .Y(_01649_));
NAND_g _21850_ (.A(_14260_), .B(_14268_), .Y(_01650_));
NAND_g _21851_ (.A(mem_la_wdata[0]), .B(_01649_), .Y(_01651_));
NAND_g _21852_ (.A(mem_wdata[0]), .B(_01650_), .Y(_01652_));
NAND_g _21853_ (.A(_01651_), .B(_01652_), .Y(_00476_));
AND_g _21854_ (.A(pcpi_rs2[1]), .B(_01648_), .Y(mem_la_wdata[1]));
NAND_g _21855_ (.A(_01649_), .B(mem_la_wdata[1]), .Y(_01653_));
NAND_g _21856_ (.A(mem_wdata[1]), .B(_01650_), .Y(_01654_));
NAND_g _21857_ (.A(_01653_), .B(_01654_), .Y(_00477_));
AND_g _21858_ (.A(pcpi_rs2[2]), .B(_01648_), .Y(mem_la_wdata[2]));
NAND_g _21859_ (.A(_01649_), .B(mem_la_wdata[2]), .Y(_01655_));
NAND_g _21860_ (.A(mem_wdata[2]), .B(_01650_), .Y(_01656_));
NAND_g _21861_ (.A(_01655_), .B(_01656_), .Y(_00478_));
AND_g _21862_ (.A(pcpi_rs2[3]), .B(_01648_), .Y(mem_la_wdata[3]));
NAND_g _21863_ (.A(_01649_), .B(mem_la_wdata[3]), .Y(_01657_));
NAND_g _21864_ (.A(mem_wdata[3]), .B(_01650_), .Y(_01658_));
NAND_g _21865_ (.A(_01657_), .B(_01658_), .Y(_00479_));
AND_g _21866_ (.A(pcpi_rs2[4]), .B(_01648_), .Y(mem_la_wdata[4]));
NAND_g _21867_ (.A(_01649_), .B(mem_la_wdata[4]), .Y(_01659_));
NAND_g _21868_ (.A(mem_wdata[4]), .B(_01650_), .Y(_01660_));
NAND_g _21869_ (.A(_01659_), .B(_01660_), .Y(_00480_));
AND_g _21870_ (.A(pcpi_rs2[5]), .B(_01648_), .Y(mem_la_wdata[5]));
NAND_g _21871_ (.A(_01649_), .B(mem_la_wdata[5]), .Y(_01661_));
NAND_g _21872_ (.A(mem_wdata[5]), .B(_01650_), .Y(_01662_));
NAND_g _21873_ (.A(_01661_), .B(_01662_), .Y(_00481_));
AND_g _21874_ (.A(pcpi_rs2[6]), .B(_01648_), .Y(mem_la_wdata[6]));
NAND_g _21875_ (.A(_01649_), .B(mem_la_wdata[6]), .Y(_01663_));
NAND_g _21876_ (.A(mem_wdata[6]), .B(_01650_), .Y(_01664_));
NAND_g _21877_ (.A(_01663_), .B(_01664_), .Y(_00482_));
AND_g _21878_ (.A(pcpi_rs2[7]), .B(_01648_), .Y(mem_la_wdata[7]));
NAND_g _21879_ (.A(_01649_), .B(mem_la_wdata[7]), .Y(_01665_));
NAND_g _21880_ (.A(mem_wdata[7]), .B(_01650_), .Y(_01666_));
NAND_g _21881_ (.A(_01665_), .B(_01666_), .Y(_00483_));
AND_g _21882_ (.A(_08842_), .B(mem_wordsize[1]), .Y(_01667_));
NAND_g _21883_ (.A(pcpi_rs2[0]), .B(_01667_), .Y(_01668_));
NAND_g _21884_ (.A(pcpi_rs2[8]), .B(_08843_), .Y(_01669_));
NAND_g _21885_ (.A(_01668_), .B(_01669_), .Y(mem_la_wdata[8]));
NAND_g _21886_ (.A(mem_wdata[8]), .B(_01650_), .Y(_01670_));
NAND_g _21887_ (.A(_01649_), .B(mem_la_wdata[8]), .Y(_01671_));
NAND_g _21888_ (.A(_01670_), .B(_01671_), .Y(_00484_));
NAND_g _21889_ (.A(pcpi_rs2[1]), .B(_01667_), .Y(_01672_));
NAND_g _21890_ (.A(pcpi_rs2[9]), .B(_08843_), .Y(_01673_));
NAND_g _21891_ (.A(_01672_), .B(_01673_), .Y(mem_la_wdata[9]));
NAND_g _21892_ (.A(mem_wdata[9]), .B(_01650_), .Y(_01674_));
NAND_g _21893_ (.A(_01649_), .B(mem_la_wdata[9]), .Y(_01675_));
NAND_g _21894_ (.A(_01674_), .B(_01675_), .Y(_00485_));
NAND_g _21895_ (.A(pcpi_rs2[2]), .B(_01667_), .Y(_01676_));
NAND_g _21896_ (.A(pcpi_rs2[10]), .B(_08843_), .Y(_01677_));
NAND_g _21897_ (.A(_01676_), .B(_01677_), .Y(mem_la_wdata[10]));
NAND_g _21898_ (.A(mem_wdata[10]), .B(_01650_), .Y(_01678_));
NAND_g _21899_ (.A(_01649_), .B(mem_la_wdata[10]), .Y(_01679_));
NAND_g _21900_ (.A(_01678_), .B(_01679_), .Y(_00486_));
NAND_g _21901_ (.A(pcpi_rs2[3]), .B(_01667_), .Y(_01680_));
NAND_g _21902_ (.A(pcpi_rs2[11]), .B(_08843_), .Y(_01681_));
NAND_g _21903_ (.A(_01680_), .B(_01681_), .Y(mem_la_wdata[11]));
NAND_g _21904_ (.A(mem_wdata[11]), .B(_01650_), .Y(_01682_));
NAND_g _21905_ (.A(_01649_), .B(mem_la_wdata[11]), .Y(_01683_));
NAND_g _21906_ (.A(_01682_), .B(_01683_), .Y(_00487_));
NAND_g _21907_ (.A(pcpi_rs2[4]), .B(_01667_), .Y(_01684_));
NAND_g _21908_ (.A(pcpi_rs2[12]), .B(_08843_), .Y(_01685_));
NAND_g _21909_ (.A(_01684_), .B(_01685_), .Y(mem_la_wdata[12]));
NAND_g _21910_ (.A(mem_wdata[12]), .B(_01650_), .Y(_01686_));
NAND_g _21911_ (.A(_01649_), .B(mem_la_wdata[12]), .Y(_01687_));
NAND_g _21912_ (.A(_01686_), .B(_01687_), .Y(_00488_));
NAND_g _21913_ (.A(pcpi_rs2[5]), .B(_01667_), .Y(_01688_));
NAND_g _21914_ (.A(pcpi_rs2[13]), .B(_08843_), .Y(_01689_));
NAND_g _21915_ (.A(_01688_), .B(_01689_), .Y(mem_la_wdata[13]));
NAND_g _21916_ (.A(mem_wdata[13]), .B(_01650_), .Y(_01690_));
NAND_g _21917_ (.A(_01649_), .B(mem_la_wdata[13]), .Y(_01691_));
NAND_g _21918_ (.A(_01690_), .B(_01691_), .Y(_00489_));
NAND_g _21919_ (.A(pcpi_rs2[6]), .B(_01667_), .Y(_01692_));
NAND_g _21920_ (.A(pcpi_rs2[14]), .B(_08843_), .Y(_01693_));
NAND_g _21921_ (.A(_01692_), .B(_01693_), .Y(mem_la_wdata[14]));
NAND_g _21922_ (.A(mem_wdata[14]), .B(_01650_), .Y(_01694_));
NAND_g _21923_ (.A(_01649_), .B(mem_la_wdata[14]), .Y(_01695_));
NAND_g _21924_ (.A(_01694_), .B(_01695_), .Y(_00490_));
NAND_g _21925_ (.A(pcpi_rs2[7]), .B(_01667_), .Y(_01696_));
NAND_g _21926_ (.A(pcpi_rs2[15]), .B(_08843_), .Y(_01697_));
NAND_g _21927_ (.A(_01696_), .B(_01697_), .Y(mem_la_wdata[15]));
NAND_g _21928_ (.A(mem_wdata[15]), .B(_01650_), .Y(_01698_));
NAND_g _21929_ (.A(_01649_), .B(mem_la_wdata[15]), .Y(_01699_));
NAND_g _21930_ (.A(_01698_), .B(_01699_), .Y(_00491_));
NOR_g _21931_ (.A(mem_wordsize[0]), .B(mem_wordsize[1]), .Y(_01700_));
NAND_g _21932_ (.A(_08842_), .B(_08843_), .Y(_01701_));
NAND_g _21933_ (.A(pcpi_rs2[16]), .B(_01700_), .Y(_01702_));
NAND_g _21934_ (.A(mem_la_wdata[0]), .B(_01701_), .Y(_01703_));
NAND_g _21935_ (.A(_01702_), .B(_01703_), .Y(mem_la_wdata[16]));
NAND_g _21936_ (.A(_01649_), .B(mem_la_wdata[16]), .Y(_01704_));
NAND_g _21937_ (.A(mem_wdata[16]), .B(_01650_), .Y(_01705_));
NAND_g _21938_ (.A(_01704_), .B(_01705_), .Y(_00492_));
NAND_g _21939_ (.A(pcpi_rs2[17]), .B(_01700_), .Y(_01706_));
NAND_g _21940_ (.A(mem_la_wdata[1]), .B(_01701_), .Y(_01707_));
NAND_g _21941_ (.A(_01706_), .B(_01707_), .Y(mem_la_wdata[17]));
NAND_g _21942_ (.A(_01649_), .B(mem_la_wdata[17]), .Y(_01708_));
NAND_g _21943_ (.A(mem_wdata[17]), .B(_01650_), .Y(_01709_));
NAND_g _21944_ (.A(_01708_), .B(_01709_), .Y(_00493_));
NAND_g _21945_ (.A(pcpi_rs2[18]), .B(_01700_), .Y(_01710_));
NAND_g _21946_ (.A(mem_la_wdata[2]), .B(_01701_), .Y(_01711_));
NAND_g _21947_ (.A(_01710_), .B(_01711_), .Y(mem_la_wdata[18]));
NAND_g _21948_ (.A(_01649_), .B(mem_la_wdata[18]), .Y(_01712_));
NAND_g _21949_ (.A(mem_wdata[18]), .B(_01650_), .Y(_01713_));
NAND_g _21950_ (.A(_01712_), .B(_01713_), .Y(_00494_));
NAND_g _21951_ (.A(pcpi_rs2[19]), .B(_01700_), .Y(_01714_));
NAND_g _21952_ (.A(mem_la_wdata[3]), .B(_01701_), .Y(_01715_));
NAND_g _21953_ (.A(_01714_), .B(_01715_), .Y(mem_la_wdata[19]));
NAND_g _21954_ (.A(_01649_), .B(mem_la_wdata[19]), .Y(_01716_));
NAND_g _21955_ (.A(mem_wdata[19]), .B(_01650_), .Y(_01717_));
NAND_g _21956_ (.A(_01716_), .B(_01717_), .Y(_00495_));
NAND_g _21957_ (.A(pcpi_rs2[20]), .B(_01700_), .Y(_01718_));
NAND_g _21958_ (.A(mem_la_wdata[4]), .B(_01701_), .Y(_01719_));
NAND_g _21959_ (.A(_01718_), .B(_01719_), .Y(mem_la_wdata[20]));
NAND_g _21960_ (.A(_01649_), .B(mem_la_wdata[20]), .Y(_01720_));
NAND_g _21961_ (.A(mem_wdata[20]), .B(_01650_), .Y(_01721_));
NAND_g _21962_ (.A(_01720_), .B(_01721_), .Y(_00496_));
NAND_g _21963_ (.A(pcpi_rs2[21]), .B(_01700_), .Y(_01722_));
NAND_g _21964_ (.A(mem_la_wdata[5]), .B(_01701_), .Y(_01723_));
NAND_g _21965_ (.A(_01722_), .B(_01723_), .Y(mem_la_wdata[21]));
NAND_g _21966_ (.A(_01649_), .B(mem_la_wdata[21]), .Y(_01724_));
NAND_g _21967_ (.A(mem_wdata[21]), .B(_01650_), .Y(_01725_));
NAND_g _21968_ (.A(_01724_), .B(_01725_), .Y(_00497_));
NAND_g _21969_ (.A(pcpi_rs2[22]), .B(_01700_), .Y(_01726_));
NAND_g _21970_ (.A(mem_la_wdata[6]), .B(_01701_), .Y(_01727_));
NAND_g _21971_ (.A(_01726_), .B(_01727_), .Y(mem_la_wdata[22]));
NAND_g _21972_ (.A(_01649_), .B(mem_la_wdata[22]), .Y(_01728_));
NAND_g _21973_ (.A(mem_wdata[22]), .B(_01650_), .Y(_01729_));
NAND_g _21974_ (.A(_01728_), .B(_01729_), .Y(_00498_));
NAND_g _21975_ (.A(pcpi_rs2[23]), .B(_01700_), .Y(_01730_));
NAND_g _21976_ (.A(mem_la_wdata[7]), .B(_01701_), .Y(_01731_));
NAND_g _21977_ (.A(_01730_), .B(_01731_), .Y(mem_la_wdata[23]));
NAND_g _21978_ (.A(_01649_), .B(mem_la_wdata[23]), .Y(_01732_));
NAND_g _21979_ (.A(mem_wdata[23]), .B(_01650_), .Y(_01733_));
NAND_g _21980_ (.A(_01732_), .B(_01733_), .Y(_00499_));
AND_g _21981_ (.A(mem_wordsize[0]), .B(_08843_), .Y(_01734_));
NAND_g _21982_ (.A(pcpi_rs2[8]), .B(_01734_), .Y(_01735_));
NAND_g _21983_ (.A(pcpi_rs2[24]), .B(_01700_), .Y(_01736_));
AND_g _21984_ (.A(_01668_), .B(_01735_), .Y(_01737_));
NAND_g _21985_ (.A(_01736_), .B(_01737_), .Y(mem_la_wdata[24]));
NAND_g _21986_ (.A(mem_wdata[24]), .B(_01650_), .Y(_01738_));
NAND_g _21987_ (.A(_01649_), .B(mem_la_wdata[24]), .Y(_01739_));
NAND_g _21988_ (.A(_01738_), .B(_01739_), .Y(_00500_));
NAND_g _21989_ (.A(pcpi_rs2[25]), .B(_01700_), .Y(_01740_));
NAND_g _21990_ (.A(pcpi_rs2[9]), .B(_01734_), .Y(_01741_));
AND_g _21991_ (.A(_01672_), .B(_01741_), .Y(_01742_));
NAND_g _21992_ (.A(_01740_), .B(_01742_), .Y(mem_la_wdata[25]));
NAND_g _21993_ (.A(mem_wdata[25]), .B(_01650_), .Y(_01743_));
NAND_g _21994_ (.A(_01649_), .B(mem_la_wdata[25]), .Y(_01744_));
NAND_g _21995_ (.A(_01743_), .B(_01744_), .Y(_00501_));
NAND_g _21996_ (.A(pcpi_rs2[26]), .B(_01700_), .Y(_01745_));
NAND_g _21997_ (.A(pcpi_rs2[10]), .B(_01734_), .Y(_01746_));
AND_g _21998_ (.A(_01676_), .B(_01746_), .Y(_01747_));
NAND_g _21999_ (.A(_01745_), .B(_01747_), .Y(mem_la_wdata[26]));
NAND_g _22000_ (.A(mem_wdata[26]), .B(_01650_), .Y(_01748_));
NAND_g _22001_ (.A(_01649_), .B(mem_la_wdata[26]), .Y(_01749_));
NAND_g _22002_ (.A(_01748_), .B(_01749_), .Y(_00502_));
NAND_g _22003_ (.A(pcpi_rs2[11]), .B(_01734_), .Y(_01750_));
NAND_g _22004_ (.A(pcpi_rs2[27]), .B(_01700_), .Y(_01751_));
AND_g _22005_ (.A(_01680_), .B(_01750_), .Y(_01752_));
NAND_g _22006_ (.A(_01751_), .B(_01752_), .Y(mem_la_wdata[27]));
NAND_g _22007_ (.A(mem_wdata[27]), .B(_01650_), .Y(_01753_));
NAND_g _22008_ (.A(_01649_), .B(mem_la_wdata[27]), .Y(_01754_));
NAND_g _22009_ (.A(_01753_), .B(_01754_), .Y(_00503_));
NAND_g _22010_ (.A(pcpi_rs2[12]), .B(_01734_), .Y(_01755_));
NAND_g _22011_ (.A(pcpi_rs2[28]), .B(_01700_), .Y(_01756_));
AND_g _22012_ (.A(_01684_), .B(_01755_), .Y(_01757_));
NAND_g _22013_ (.A(_01756_), .B(_01757_), .Y(mem_la_wdata[28]));
NAND_g _22014_ (.A(mem_wdata[28]), .B(_01650_), .Y(_01758_));
NAND_g _22015_ (.A(_01649_), .B(mem_la_wdata[28]), .Y(_01759_));
NAND_g _22016_ (.A(_01758_), .B(_01759_), .Y(_00504_));
NAND_g _22017_ (.A(pcpi_rs2[13]), .B(_01734_), .Y(_01760_));
NAND_g _22018_ (.A(pcpi_rs2[29]), .B(_01700_), .Y(_01761_));
AND_g _22019_ (.A(_01688_), .B(_01760_), .Y(_01762_));
NAND_g _22020_ (.A(_01761_), .B(_01762_), .Y(mem_la_wdata[29]));
NAND_g _22021_ (.A(mem_wdata[29]), .B(_01650_), .Y(_01763_));
NAND_g _22022_ (.A(_01649_), .B(mem_la_wdata[29]), .Y(_01764_));
NAND_g _22023_ (.A(_01763_), .B(_01764_), .Y(_00505_));
NAND_g _22024_ (.A(pcpi_rs2[14]), .B(_01734_), .Y(_01765_));
NAND_g _22025_ (.A(pcpi_rs2[30]), .B(_01700_), .Y(_01766_));
AND_g _22026_ (.A(_01692_), .B(_01765_), .Y(_01767_));
NAND_g _22027_ (.A(_01766_), .B(_01767_), .Y(mem_la_wdata[30]));
NAND_g _22028_ (.A(mem_wdata[30]), .B(_01650_), .Y(_01768_));
NAND_g _22029_ (.A(_01649_), .B(mem_la_wdata[30]), .Y(_01769_));
NAND_g _22030_ (.A(_01768_), .B(_01769_), .Y(_00506_));
NAND_g _22031_ (.A(pcpi_rs2[15]), .B(_01734_), .Y(_01770_));
NAND_g _22032_ (.A(pcpi_rs2[31]), .B(_01700_), .Y(_01771_));
AND_g _22033_ (.A(_01696_), .B(_01770_), .Y(_01772_));
NAND_g _22034_ (.A(_01771_), .B(_01772_), .Y(mem_la_wdata[31]));
NAND_g _22035_ (.A(mem_wdata[31]), .B(_01650_), .Y(_01773_));
NAND_g _22036_ (.A(_01649_), .B(mem_la_wdata[31]), .Y(_01774_));
NAND_g _22037_ (.A(_01773_), .B(_01774_), .Y(_00507_));
NAND_g _22038_ (.A(mem_wstrb[0]), .B(_14271_), .Y(_01775_));
NOR_g _22039_ (.A(mem_wordsize[0]), .B(pcpi_rs1[1]), .Y(_01776_));
NAND_g _22040_ (.A(_08961_), .B(_01776_), .Y(_01777_));
AND_g _22041_ (.A(mem_wordsize[0]), .B(pcpi_rs1[1]), .Y(_01778_));
NAND_g _22042_ (.A(mem_wordsize[0]), .B(pcpi_rs1[1]), .Y(_01779_));
AND_g _22043_ (.A(_08843_), .B(_01779_), .Y(_01780_));
NAND_g _22044_ (.A(_08843_), .B(_01779_), .Y(_01781_));
NAND_g _22045_ (.A(_01777_), .B(_01781_), .Y(mem_la_wstrb[0]));
NOR_g _22046_ (.A(_14269_), .B(_01650_), .Y(_01782_));
NAND_g _22047_ (.A(mem_la_wstrb[0]), .B(_01782_), .Y(_01783_));
NAND_g _22048_ (.A(_01775_), .B(_01783_), .Y(_00508_));
NAND_g _22049_ (.A(pcpi_rs1[0]), .B(_01776_), .Y(_01784_));
NAND_g _22050_ (.A(_01781_), .B(_01784_), .Y(mem_la_wstrb[1]));
NAND_g _22051_ (.A(_01782_), .B(mem_la_wstrb[1]), .Y(_01785_));
NAND_g _22052_ (.A(mem_wstrb[1]), .B(_14271_), .Y(_01786_));
NAND_g _22053_ (.A(_01785_), .B(_01786_), .Y(_00509_));
AND_g _22054_ (.A(pcpi_rs1[1]), .B(_01667_), .Y(_01787_));
NAND_g _22055_ (.A(_08961_), .B(_01787_), .Y(_01788_));
AND_g _22056_ (.A(_08843_), .B(_01778_), .Y(_01789_));
NAND_g _22057_ (.A(_08843_), .B(_01778_), .Y(_01790_));
NAND_g _22058_ (.A(_01788_), .B(_01790_), .Y(_01791_));
NOT_g _22059_ (.A(_01791_), .Y(_01792_));
NAND_g _22060_ (.A(_01701_), .B(_01792_), .Y(mem_la_wstrb[2]));
NAND_g _22061_ (.A(_01782_), .B(mem_la_wstrb[2]), .Y(_01793_));
NAND_g _22062_ (.A(mem_wstrb[2]), .B(_14271_), .Y(_01794_));
NAND_g _22063_ (.A(_01793_), .B(_01794_), .Y(_00510_));
NAND_g _22064_ (.A(mem_wstrb[3]), .B(_14271_), .Y(_01795_));
AND_g _22065_ (.A(pcpi_rs1[0]), .B(_01787_), .Y(_01796_));
NOR_g _22066_ (.A(_01700_), .B(_01796_), .Y(_01797_));
NAND_g _22067_ (.A(_01790_), .B(_01797_), .Y(mem_la_wstrb[3]));
NAND_g _22068_ (.A(_01782_), .B(mem_la_wstrb[3]), .Y(_01798_));
NAND_g _22069_ (.A(_01795_), .B(_01798_), .Y(_00511_));
AND_g _22070_ (.A(_14273_), .B(_14278_), .Y(_01799_));
NAND_g _22071_ (.A(_08804_), .B(_14272_), .Y(_01800_));
AND_g _22072_ (.A(_14279_), .B(_01800_), .Y(_01801_));
NAND_g _22073_ (.A(_01799_), .B(_01801_), .Y(_01802_));
NAND_g _22074_ (.A(mem_state[0]), .B(_01802_), .Y(_01803_));
AND_g _22075_ (.A(mem_state[0]), .B(_08873_), .Y(_01804_));
AND_g _22076_ (.A(_09903_), .B(_01804_), .Y(_01805_));
AND_g _22077_ (.A(_09899_), .B(_14260_), .Y(_01806_));
NAND_g _22078_ (.A(_01805_), .B(_01806_), .Y(_01807_));
NAND_g _22079_ (.A(_14265_), .B(_14281_), .Y(_01808_));
AND_g _22080_ (.A(_01807_), .B(_01808_), .Y(_01809_));
NAND_g _22081_ (.A(_01803_), .B(_01809_), .Y(_00512_));
NAND_g _22082_ (.A(mem_state[1]), .B(_01802_), .Y(_01810_));
AND_g _22083_ (.A(_01650_), .B(_01807_), .Y(_01811_));
NAND_g _22084_ (.A(_01810_), .B(_01811_), .Y(_00513_));
NOR_g _22085_ (.A(decoded_imm[31]), .B(_13840_), .Y(_01812_));
NAND_g _22086_ (.A(mem_rdata_q[31]), .B(_10738_), .Y(_01813_));
NAND_g _22087_ (.A(mem_rdata_q[31]), .B(_14864_), .Y(_01814_));
AND_g _22088_ (.A(_13840_), .B(_01814_), .Y(_01815_));
NAND_g _22089_ (.A(instr_jal), .B(decoded_imm_j[31]), .Y(_01816_));
NOR_g _22090_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(is_sb_sh_sw), .Y(_01817_));
NAND_g _22091_ (.A(_08790_), .B(_08864_), .Y(_01818_));
NAND_g _22092_ (.A(mem_rdata_q[31]), .B(_01818_), .Y(_01819_));
AND_g _22093_ (.A(_01816_), .B(_01819_), .Y(_01820_));
AND_g _22094_ (.A(_01815_), .B(_01820_), .Y(_01821_));
AND_g _22095_ (.A(_01813_), .B(_01821_), .Y(_01822_));
NOR_g _22096_ (.A(_01812_), .B(_01822_), .Y(_00521_));
NOR_g _22097_ (.A(decoded_imm[30]), .B(_13840_), .Y(_01823_));
NAND_g _22098_ (.A(mem_rdata_q[30]), .B(_10738_), .Y(_01824_));
AND_g _22099_ (.A(_01821_), .B(_01824_), .Y(_01825_));
NOR_g _22100_ (.A(_01823_), .B(_01825_), .Y(_00522_));
NOR_g _22101_ (.A(decoded_imm[29]), .B(_13840_), .Y(_01826_));
NAND_g _22102_ (.A(mem_rdata_q[29]), .B(_10738_), .Y(_01827_));
AND_g _22103_ (.A(_01821_), .B(_01827_), .Y(_01828_));
NOR_g _22104_ (.A(_01826_), .B(_01828_), .Y(_00523_));
NOR_g _22105_ (.A(decoded_imm[28]), .B(_13840_), .Y(_01829_));
NAND_g _22106_ (.A(mem_rdata_q[28]), .B(_10738_), .Y(_01830_));
AND_g _22107_ (.A(_01821_), .B(_01830_), .Y(_01831_));
NOR_g _22108_ (.A(_01829_), .B(_01831_), .Y(_00524_));
NOR_g _22109_ (.A(decoded_imm[27]), .B(_13840_), .Y(_01832_));
NAND_g _22110_ (.A(mem_rdata_q[27]), .B(_10738_), .Y(_01833_));
AND_g _22111_ (.A(_01821_), .B(_01833_), .Y(_01834_));
NOR_g _22112_ (.A(_01832_), .B(_01834_), .Y(_00525_));
NOR_g _22113_ (.A(decoded_imm[26]), .B(_13840_), .Y(_01835_));
NAND_g _22114_ (.A(mem_rdata_q[26]), .B(_10738_), .Y(_01836_));
AND_g _22115_ (.A(_01821_), .B(_01836_), .Y(_01837_));
NOR_g _22116_ (.A(_01835_), .B(_01837_), .Y(_00526_));
NOR_g _22117_ (.A(decoded_imm[25]), .B(_13840_), .Y(_01838_));
NAND_g _22118_ (.A(mem_rdata_q[25]), .B(_10738_), .Y(_01839_));
AND_g _22119_ (.A(_01821_), .B(_01839_), .Y(_01840_));
NOR_g _22120_ (.A(_01838_), .B(_01840_), .Y(_00527_));
NOR_g _22121_ (.A(decoded_imm[24]), .B(_13840_), .Y(_01841_));
NAND_g _22122_ (.A(mem_rdata_q[24]), .B(_10738_), .Y(_01842_));
AND_g _22123_ (.A(_01821_), .B(_01842_), .Y(_01843_));
NOR_g _22124_ (.A(_01841_), .B(_01843_), .Y(_00528_));
NOR_g _22125_ (.A(decoded_imm[23]), .B(_13840_), .Y(_01844_));
NAND_g _22126_ (.A(mem_rdata_q[23]), .B(_10738_), .Y(_01845_));
AND_g _22127_ (.A(_01821_), .B(_01845_), .Y(_01846_));
NOR_g _22128_ (.A(_01844_), .B(_01846_), .Y(_00529_));
NOR_g _22129_ (.A(decoded_imm[22]), .B(_13840_), .Y(_01847_));
NAND_g _22130_ (.A(mem_rdata_q[22]), .B(_10738_), .Y(_01848_));
AND_g _22131_ (.A(_01821_), .B(_01848_), .Y(_01849_));
NOR_g _22132_ (.A(_01847_), .B(_01849_), .Y(_00530_));
NOR_g _22133_ (.A(decoded_imm[21]), .B(_13840_), .Y(_01850_));
NAND_g _22134_ (.A(mem_rdata_q[21]), .B(_10738_), .Y(_01851_));
AND_g _22135_ (.A(_01821_), .B(_01851_), .Y(_01852_));
NOR_g _22136_ (.A(_01850_), .B(_01852_), .Y(_00531_));
NOR_g _22137_ (.A(decoded_imm[20]), .B(_13840_), .Y(_01853_));
NAND_g _22138_ (.A(mem_rdata_q[20]), .B(_10738_), .Y(_01854_));
AND_g _22139_ (.A(_01821_), .B(_01854_), .Y(_01855_));
NOR_g _22140_ (.A(_01853_), .B(_01855_), .Y(_00532_));
NOR_g _22141_ (.A(decoded_imm[19]), .B(_13840_), .Y(_01856_));
NAND_g _22142_ (.A(instr_jal), .B(decoded_imm_j[19]), .Y(_01857_));
NAND_g _22143_ (.A(mem_rdata_q[19]), .B(_10738_), .Y(_01858_));
AND_g _22144_ (.A(_01857_), .B(_01858_), .Y(_01859_));
AND_g _22145_ (.A(_01815_), .B(_01819_), .Y(_01860_));
AND_g _22146_ (.A(_01859_), .B(_01860_), .Y(_01861_));
NOR_g _22147_ (.A(_01856_), .B(_01861_), .Y(_00533_));
NOR_g _22148_ (.A(decoded_imm[18]), .B(_13840_), .Y(_01862_));
NAND_g _22149_ (.A(instr_jal), .B(decoded_imm_j[18]), .Y(_01863_));
NAND_g _22150_ (.A(mem_rdata_q[18]), .B(_10738_), .Y(_01864_));
AND_g _22151_ (.A(_01863_), .B(_01864_), .Y(_01865_));
AND_g _22152_ (.A(_01860_), .B(_01865_), .Y(_01866_));
NOR_g _22153_ (.A(_01862_), .B(_01866_), .Y(_00534_));
NOR_g _22154_ (.A(decoded_imm[17]), .B(_13840_), .Y(_01867_));
NAND_g _22155_ (.A(mem_rdata_q[17]), .B(_10738_), .Y(_01868_));
NAND_g _22156_ (.A(instr_jal), .B(decoded_imm_j[17]), .Y(_01869_));
AND_g _22157_ (.A(_01868_), .B(_01869_), .Y(_01870_));
AND_g _22158_ (.A(_01860_), .B(_01870_), .Y(_01871_));
NOR_g _22159_ (.A(_01867_), .B(_01871_), .Y(_00535_));
NOR_g _22160_ (.A(decoded_imm[16]), .B(_13840_), .Y(_01872_));
NAND_g _22161_ (.A(mem_rdata_q[16]), .B(_10738_), .Y(_01873_));
NAND_g _22162_ (.A(instr_jal), .B(decoded_imm_j[16]), .Y(_01874_));
AND_g _22163_ (.A(_01873_), .B(_01874_), .Y(_01875_));
AND_g _22164_ (.A(_01860_), .B(_01875_), .Y(_01876_));
NOR_g _22165_ (.A(_01872_), .B(_01876_), .Y(_00536_));
NOR_g _22166_ (.A(decoded_imm[15]), .B(_13840_), .Y(_01877_));
NAND_g _22167_ (.A(instr_jal), .B(decoded_imm_j[15]), .Y(_01878_));
NAND_g _22168_ (.A(mem_rdata_q[15]), .B(_10738_), .Y(_01879_));
AND_g _22169_ (.A(_01878_), .B(_01879_), .Y(_01880_));
AND_g _22170_ (.A(_01860_), .B(_01880_), .Y(_01881_));
NOR_g _22171_ (.A(_01877_), .B(_01881_), .Y(_00537_));
NOR_g _22172_ (.A(decoded_imm[14]), .B(_13840_), .Y(_01882_));
AND_g _22173_ (.A(instr_jal), .B(decoded_imm_j[14]), .Y(_01883_));
NOR_g _22174_ (.A(_08867_), .B(_10737_), .Y(_01884_));
NOR_g _22175_ (.A(_01883_), .B(_01884_), .Y(_01885_));
AND_g _22176_ (.A(_01860_), .B(_01885_), .Y(_01886_));
NOR_g _22177_ (.A(_01882_), .B(_01886_), .Y(_00538_));
NOR_g _22178_ (.A(decoded_imm[13]), .B(_13840_), .Y(_01887_));
AND_g _22179_ (.A(instr_jal), .B(decoded_imm_j[13]), .Y(_01888_));
NOR_g _22180_ (.A(_08866_), .B(_10737_), .Y(_01889_));
NOR_g _22181_ (.A(_01888_), .B(_01889_), .Y(_01890_));
AND_g _22182_ (.A(_01860_), .B(_01890_), .Y(_01891_));
NOR_g _22183_ (.A(_01887_), .B(_01891_), .Y(_00539_));
NOR_g _22184_ (.A(decoded_imm[12]), .B(_13840_), .Y(_01892_));
NOR_g _22185_ (.A(_08865_), .B(_10737_), .Y(_01893_));
AND_g _22186_ (.A(instr_jal), .B(decoded_imm_j[12]), .Y(_01894_));
NOR_g _22187_ (.A(_01893_), .B(_01894_), .Y(_01895_));
AND_g _22188_ (.A(_01860_), .B(_01895_), .Y(_01896_));
NOR_g _22189_ (.A(_01892_), .B(_01896_), .Y(_00540_));
NOR_g _22190_ (.A(decoded_imm[11]), .B(_13840_), .Y(_01897_));
NAND_g _22191_ (.A(is_sb_sh_sw), .B(mem_rdata_q[31]), .Y(_01898_));
NAND_g _22192_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(mem_rdata_q[7]), .Y(_01899_));
NAND_g _22193_ (.A(instr_jal), .B(decoded_imm_j[11]), .Y(_01900_));
AND_g _22194_ (.A(_01899_), .B(_01900_), .Y(_01901_));
AND_g _22195_ (.A(_01898_), .B(_01901_), .Y(_01902_));
AND_g _22196_ (.A(_01815_), .B(_01902_), .Y(_01903_));
NOR_g _22197_ (.A(_01897_), .B(_01903_), .Y(_00541_));
NAND_g _22198_ (.A(_14865_), .B(_01817_), .Y(_01904_));
NAND_g _22199_ (.A(mem_rdata_q[30]), .B(_01904_), .Y(_01905_));
NAND_g _22200_ (.A(instr_jal), .B(decoded_imm_j[10]), .Y(_01906_));
NOR_g _22201_ (.A(decoded_imm[10]), .B(_13840_), .Y(_01907_));
AND_g _22202_ (.A(_13840_), .B(_01906_), .Y(_01908_));
AND_g _22203_ (.A(_01905_), .B(_01908_), .Y(_01909_));
NOR_g _22204_ (.A(_01907_), .B(_01909_), .Y(_00542_));
NAND_g _22205_ (.A(mem_rdata_q[29]), .B(_01904_), .Y(_01910_));
NAND_g _22206_ (.A(instr_jal), .B(decoded_imm_j[9]), .Y(_01911_));
NOR_g _22207_ (.A(decoded_imm[9]), .B(_13840_), .Y(_01912_));
AND_g _22208_ (.A(_13840_), .B(_01911_), .Y(_01913_));
AND_g _22209_ (.A(_01910_), .B(_01913_), .Y(_01914_));
NOR_g _22210_ (.A(_01912_), .B(_01914_), .Y(_00543_));
NAND_g _22211_ (.A(mem_rdata_q[28]), .B(_01904_), .Y(_01915_));
NAND_g _22212_ (.A(instr_jal), .B(decoded_imm_j[8]), .Y(_01916_));
NOR_g _22213_ (.A(decoded_imm[8]), .B(_13840_), .Y(_01917_));
AND_g _22214_ (.A(_13840_), .B(_01916_), .Y(_01918_));
AND_g _22215_ (.A(_01915_), .B(_01918_), .Y(_01919_));
NOR_g _22216_ (.A(_01917_), .B(_01919_), .Y(_00544_));
NAND_g _22217_ (.A(mem_rdata_q[27]), .B(_01904_), .Y(_01920_));
NAND_g _22218_ (.A(instr_jal), .B(decoded_imm_j[7]), .Y(_01921_));
NOR_g _22219_ (.A(decoded_imm[7]), .B(_13840_), .Y(_01922_));
AND_g _22220_ (.A(_13840_), .B(_01921_), .Y(_01923_));
AND_g _22221_ (.A(_01920_), .B(_01923_), .Y(_01924_));
NOR_g _22222_ (.A(_01922_), .B(_01924_), .Y(_00545_));
NAND_g _22223_ (.A(mem_rdata_q[26]), .B(_01904_), .Y(_01925_));
NAND_g _22224_ (.A(instr_jal), .B(decoded_imm_j[6]), .Y(_01926_));
NOR_g _22225_ (.A(decoded_imm[6]), .B(_13840_), .Y(_01927_));
AND_g _22226_ (.A(_13840_), .B(_01926_), .Y(_01928_));
AND_g _22227_ (.A(_01925_), .B(_01928_), .Y(_01929_));
NOR_g _22228_ (.A(_01927_), .B(_01929_), .Y(_00546_));
NAND_g _22229_ (.A(mem_rdata_q[25]), .B(_01904_), .Y(_01930_));
NAND_g _22230_ (.A(instr_jal), .B(decoded_imm_j[5]), .Y(_01931_));
NOR_g _22231_ (.A(decoded_imm[5]), .B(_13840_), .Y(_01932_));
AND_g _22232_ (.A(_13840_), .B(_01931_), .Y(_01933_));
AND_g _22233_ (.A(_01930_), .B(_01933_), .Y(_01934_));
NOR_g _22234_ (.A(_01932_), .B(_01934_), .Y(_00547_));
NAND_g _22235_ (.A(mem_rdata_q[24]), .B(_14864_), .Y(_01935_));
NAND_g _22236_ (.A(instr_jal), .B(decoded_imm_j[4]), .Y(_01936_));
NAND_g _22237_ (.A(mem_rdata_q[11]), .B(_01818_), .Y(_01937_));
AND_g _22238_ (.A(_13840_), .B(_01936_), .Y(_01938_));
AND_g _22239_ (.A(_01937_), .B(_01938_), .Y(_01939_));
AND_g _22240_ (.A(_01935_), .B(_01939_), .Y(_01940_));
NOR_g _22241_ (.A(decoded_imm[4]), .B(_13840_), .Y(_01941_));
NOR_g _22242_ (.A(_01940_), .B(_01941_), .Y(_00548_));
NAND_g _22243_ (.A(mem_rdata_q[23]), .B(_14864_), .Y(_01942_));
NAND_g _22244_ (.A(instr_jal), .B(decoded_imm_j[3]), .Y(_01943_));
NAND_g _22245_ (.A(mem_rdata_q[10]), .B(_01818_), .Y(_01944_));
AND_g _22246_ (.A(_13840_), .B(_01943_), .Y(_01945_));
AND_g _22247_ (.A(_01944_), .B(_01945_), .Y(_01946_));
AND_g _22248_ (.A(_01942_), .B(_01946_), .Y(_01947_));
NOR_g _22249_ (.A(decoded_imm[3]), .B(_13840_), .Y(_01948_));
NOR_g _22250_ (.A(_01947_), .B(_01948_), .Y(_00549_));
NAND_g _22251_ (.A(mem_rdata_q[22]), .B(_14864_), .Y(_01949_));
NAND_g _22252_ (.A(mem_rdata_q[9]), .B(_01818_), .Y(_01950_));
NAND_g _22253_ (.A(instr_jal), .B(decoded_imm_j[2]), .Y(_01951_));
AND_g _22254_ (.A(_01950_), .B(_01951_), .Y(_01952_));
NAND_g _22255_ (.A(_01949_), .B(_01952_), .Y(_01953_));
NAND_g _22256_ (.A(_13840_), .B(_01953_), .Y(_01954_));
NAND_g _22257_ (.A(decoded_imm[2]), .B(_13841_), .Y(_01955_));
NAND_g _22258_ (.A(_01954_), .B(_01955_), .Y(_00550_));
NAND_g _22259_ (.A(mem_rdata_q[21]), .B(_14864_), .Y(_01956_));
AND_g _22260_ (.A(mem_rdata_q[8]), .B(_01818_), .Y(_01957_));
NOR_g _22261_ (.A(_10099_), .B(_01957_), .Y(_01958_));
NAND_g _22262_ (.A(_01956_), .B(_01958_), .Y(_01959_));
NAND_g _22263_ (.A(_13840_), .B(_01959_), .Y(_01960_));
NAND_g _22264_ (.A(decoded_imm[1]), .B(_13841_), .Y(_01961_));
NAND_g _22265_ (.A(_01960_), .B(_01961_), .Y(_00551_));
NAND_g _22266_ (.A(_09073_), .B(_09913_), .Y(_01962_));
AND_g _22267_ (.A(reg_next_pc[0]), .B(resetn), .Y(_01963_));
AND_g _22268_ (.A(_01962_), .B(_01963_), .Y(_00552_));
AND_g _22269_ (.A(_09499_), .B(_09825_), .Y(_01964_));
NAND_g _22270_ (.A(_09499_), .B(_09825_), .Y(_01965_));
NAND_g _22271_ (.A(_09098_), .B(_01964_), .Y(_01966_));
NAND_g _22272_ (.A(cpuregs[29][0]), .B(_01965_), .Y(_01967_));
NAND_g _22273_ (.A(_01966_), .B(_01967_), .Y(_00553_));
NAND_g _22274_ (.A(_09109_), .B(_01964_), .Y(_01968_));
NAND_g _22275_ (.A(cpuregs[29][1]), .B(_01965_), .Y(_01969_));
NAND_g _22276_ (.A(_01968_), .B(_01969_), .Y(_00554_));
NAND_g _22277_ (.A(_09118_), .B(_01964_), .Y(_01970_));
NAND_g _22278_ (.A(cpuregs[29][2]), .B(_01965_), .Y(_01971_));
NAND_g _22279_ (.A(_01970_), .B(_01971_), .Y(_00555_));
NAND_g _22280_ (.A(_09131_), .B(_01964_), .Y(_01972_));
NAND_g _22281_ (.A(cpuregs[29][3]), .B(_01965_), .Y(_01973_));
NAND_g _22282_ (.A(_01972_), .B(_01973_), .Y(_00556_));
NAND_g _22283_ (.A(_09144_), .B(_01964_), .Y(_01974_));
NAND_g _22284_ (.A(cpuregs[29][4]), .B(_01965_), .Y(_01975_));
NAND_g _22285_ (.A(_01974_), .B(_01975_), .Y(_00557_));
NAND_g _22286_ (.A(_09157_), .B(_01964_), .Y(_01976_));
NAND_g _22287_ (.A(cpuregs[29][5]), .B(_01965_), .Y(_01977_));
NAND_g _22288_ (.A(_01976_), .B(_01977_), .Y(_00558_));
NAND_g _22289_ (.A(_09170_), .B(_01964_), .Y(_01978_));
NAND_g _22290_ (.A(cpuregs[29][6]), .B(_01965_), .Y(_01979_));
NAND_g _22291_ (.A(_01978_), .B(_01979_), .Y(_00559_));
NAND_g _22292_ (.A(_09183_), .B(_01964_), .Y(_01980_));
NAND_g _22293_ (.A(cpuregs[29][7]), .B(_01965_), .Y(_01981_));
NAND_g _22294_ (.A(_01980_), .B(_01981_), .Y(_00560_));
NAND_g _22295_ (.A(_09196_), .B(_01964_), .Y(_01982_));
NAND_g _22296_ (.A(cpuregs[29][8]), .B(_01965_), .Y(_01983_));
NAND_g _22297_ (.A(_01982_), .B(_01983_), .Y(_00561_));
NAND_g _22298_ (.A(_09209_), .B(_01964_), .Y(_01984_));
NAND_g _22299_ (.A(cpuregs[29][9]), .B(_01965_), .Y(_01985_));
NAND_g _22300_ (.A(_01984_), .B(_01985_), .Y(_00562_));
NAND_g _22301_ (.A(_09222_), .B(_01964_), .Y(_01986_));
NAND_g _22302_ (.A(cpuregs[29][10]), .B(_01965_), .Y(_01987_));
NAND_g _22303_ (.A(_01986_), .B(_01987_), .Y(_00563_));
NAND_g _22304_ (.A(_09235_), .B(_01964_), .Y(_01988_));
NAND_g _22305_ (.A(cpuregs[29][11]), .B(_01965_), .Y(_01989_));
NAND_g _22306_ (.A(_01988_), .B(_01989_), .Y(_00564_));
NAND_g _22307_ (.A(_09248_), .B(_01964_), .Y(_01990_));
NAND_g _22308_ (.A(cpuregs[29][12]), .B(_01965_), .Y(_01991_));
NAND_g _22309_ (.A(_01990_), .B(_01991_), .Y(_00565_));
NAND_g _22310_ (.A(_09261_), .B(_01964_), .Y(_01992_));
NAND_g _22311_ (.A(cpuregs[29][13]), .B(_01965_), .Y(_01993_));
NAND_g _22312_ (.A(_01992_), .B(_01993_), .Y(_00566_));
NAND_g _22313_ (.A(_09274_), .B(_01964_), .Y(_01994_));
NAND_g _22314_ (.A(cpuregs[29][14]), .B(_01965_), .Y(_01995_));
NAND_g _22315_ (.A(_01994_), .B(_01995_), .Y(_00567_));
NAND_g _22316_ (.A(_09287_), .B(_01964_), .Y(_01996_));
NAND_g _22317_ (.A(cpuregs[29][15]), .B(_01965_), .Y(_01997_));
NAND_g _22318_ (.A(_01996_), .B(_01997_), .Y(_00568_));
NAND_g _22319_ (.A(_09300_), .B(_01964_), .Y(_01998_));
NAND_g _22320_ (.A(cpuregs[29][16]), .B(_01965_), .Y(_01999_));
NAND_g _22321_ (.A(_01998_), .B(_01999_), .Y(_00569_));
NOR_g _22322_ (.A(cpuregs[29][17]), .B(_01964_), .Y(_02000_));
NOR_g _22323_ (.A(_09313_), .B(_01965_), .Y(_02001_));
NOR_g _22324_ (.A(_02000_), .B(_02001_), .Y(_00570_));
NAND_g _22325_ (.A(_09325_), .B(_01964_), .Y(_02002_));
NAND_g _22326_ (.A(cpuregs[29][18]), .B(_01965_), .Y(_02003_));
NAND_g _22327_ (.A(_02002_), .B(_02003_), .Y(_00571_));
NAND_g _22328_ (.A(_09338_), .B(_01964_), .Y(_02004_));
NAND_g _22329_ (.A(cpuregs[29][19]), .B(_01965_), .Y(_02005_));
NAND_g _22330_ (.A(_02004_), .B(_02005_), .Y(_00572_));
NAND_g _22331_ (.A(_09351_), .B(_01964_), .Y(_02006_));
NAND_g _22332_ (.A(cpuregs[29][20]), .B(_01965_), .Y(_02007_));
NAND_g _22333_ (.A(_02006_), .B(_02007_), .Y(_00573_));
NAND_g _22334_ (.A(_09364_), .B(_01964_), .Y(_02008_));
NAND_g _22335_ (.A(cpuregs[29][21]), .B(_01965_), .Y(_02009_));
NAND_g _22336_ (.A(_02008_), .B(_02009_), .Y(_00574_));
NAND_g _22337_ (.A(_09377_), .B(_01964_), .Y(_02010_));
NAND_g _22338_ (.A(cpuregs[29][22]), .B(_01965_), .Y(_02011_));
NAND_g _22339_ (.A(_02010_), .B(_02011_), .Y(_00575_));
NAND_g _22340_ (.A(_09390_), .B(_01964_), .Y(_02012_));
NAND_g _22341_ (.A(cpuregs[29][23]), .B(_01965_), .Y(_02013_));
NAND_g _22342_ (.A(_02012_), .B(_02013_), .Y(_00576_));
NAND_g _22343_ (.A(_09403_), .B(_01964_), .Y(_02014_));
NAND_g _22344_ (.A(cpuregs[29][24]), .B(_01965_), .Y(_02015_));
NAND_g _22345_ (.A(_02014_), .B(_02015_), .Y(_00577_));
NAND_g _22346_ (.A(_09416_), .B(_01964_), .Y(_02016_));
NAND_g _22347_ (.A(cpuregs[29][25]), .B(_01965_), .Y(_02017_));
NAND_g _22348_ (.A(_02016_), .B(_02017_), .Y(_00578_));
NAND_g _22349_ (.A(_09429_), .B(_01964_), .Y(_02018_));
NAND_g _22350_ (.A(cpuregs[29][26]), .B(_01965_), .Y(_02019_));
NAND_g _22351_ (.A(_02018_), .B(_02019_), .Y(_00579_));
NAND_g _22352_ (.A(_09442_), .B(_01964_), .Y(_02020_));
NAND_g _22353_ (.A(cpuregs[29][27]), .B(_01965_), .Y(_02021_));
NAND_g _22354_ (.A(_02020_), .B(_02021_), .Y(_00580_));
NAND_g _22355_ (.A(_09455_), .B(_01964_), .Y(_02022_));
NAND_g _22356_ (.A(cpuregs[29][28]), .B(_01965_), .Y(_02023_));
NAND_g _22357_ (.A(_02022_), .B(_02023_), .Y(_00581_));
NAND_g _22358_ (.A(_09468_), .B(_01964_), .Y(_02024_));
NAND_g _22359_ (.A(cpuregs[29][29]), .B(_01965_), .Y(_02025_));
NAND_g _22360_ (.A(_02024_), .B(_02025_), .Y(_00582_));
NAND_g _22361_ (.A(_09481_), .B(_01964_), .Y(_02026_));
NAND_g _22362_ (.A(cpuregs[29][30]), .B(_01965_), .Y(_02027_));
NAND_g _22363_ (.A(_02026_), .B(_02027_), .Y(_00583_));
NAND_g _22364_ (.A(_09493_), .B(_01964_), .Y(_02028_));
NAND_g _22365_ (.A(cpuregs[29][31]), .B(_01965_), .Y(_02029_));
NAND_g _22366_ (.A(_02028_), .B(_02029_), .Y(_00584_));
NAND_g _22367_ (.A(_14393_), .B(_00438_), .Y(_02030_));
NAND_g _22368_ (.A(decoded_imm_j[4]), .B(_14394_), .Y(_02031_));
NAND_g _22369_ (.A(_02030_), .B(_02031_), .Y(_00585_));
NAND_g _22370_ (.A(count_instr[0]), .B(_09893_), .Y(_02032_));
NOR_g _22371_ (.A(count_instr[0]), .B(_09893_), .Y(_02033_));
NOR_g _22372_ (.A(_08811_), .B(_02033_), .Y(_02034_));
AND_g _22373_ (.A(_02032_), .B(_02034_), .Y(_00586_));
AND_g _22374_ (.A(count_instr[1]), .B(count_instr[0]), .Y(_02035_));
AND_g _22375_ (.A(_09893_), .B(_02035_), .Y(_02036_));
NAND_g _22376_ (.A(_08788_), .B(_02032_), .Y(_02037_));
NAND_g _22377_ (.A(resetn), .B(_02037_), .Y(_02038_));
NOR_g _22378_ (.A(_02036_), .B(_02038_), .Y(_00587_));
NAND_g _22379_ (.A(count_instr[2]), .B(_02036_), .Y(_02039_));
NOR_g _22380_ (.A(count_instr[2]), .B(_02036_), .Y(_02040_));
NOR_g _22381_ (.A(_08811_), .B(_02040_), .Y(_02041_));
AND_g _22382_ (.A(_02039_), .B(_02041_), .Y(_00588_));
NAND_g _22383_ (.A(_08787_), .B(_02039_), .Y(_02042_));
AND_g _22384_ (.A(count_instr[3]), .B(count_instr[2]), .Y(_02043_));
AND_g _22385_ (.A(_02035_), .B(_02043_), .Y(_02044_));
AND_g _22386_ (.A(_09893_), .B(_02044_), .Y(_02045_));
NOR_g _22387_ (.A(_08811_), .B(_02045_), .Y(_02046_));
NOR_g _22388_ (.A(_08787_), .B(_02039_), .Y(_02047_));
AND_g _22389_ (.A(_02042_), .B(_02046_), .Y(_00589_));
NOR_g _22390_ (.A(count_instr[4]), .B(_02045_), .Y(_02048_));
NOR_g _22391_ (.A(_08811_), .B(_02048_), .Y(_02049_));
NAND_g _22392_ (.A(count_instr[4]), .B(_02045_), .Y(_02050_));
AND_g _22393_ (.A(_02049_), .B(_02050_), .Y(_00590_));
NAND_g _22394_ (.A(_08786_), .B(_02050_), .Y(_02051_));
AND_g _22395_ (.A(count_instr[5]), .B(count_instr[4]), .Y(_02052_));
AND_g _22396_ (.A(_02045_), .B(_02052_), .Y(_02053_));
NOR_g _22397_ (.A(_08811_), .B(_02053_), .Y(_02054_));
AND_g _22398_ (.A(_02047_), .B(_02052_), .Y(_02055_));
AND_g _22399_ (.A(_02051_), .B(_02054_), .Y(_00591_));
NOR_g _22400_ (.A(count_instr[6]), .B(_02053_), .Y(_02056_));
NOR_g _22401_ (.A(_08811_), .B(_02056_), .Y(_02057_));
AND_g _22402_ (.A(count_instr[6]), .B(_02053_), .Y(_02058_));
NAND_g _22403_ (.A(count_instr[6]), .B(_02053_), .Y(_02059_));
AND_g _22404_ (.A(_02057_), .B(_02059_), .Y(_00592_));
NOR_g _22405_ (.A(count_instr[7]), .B(_02058_), .Y(_02060_));
NOR_g _22406_ (.A(_08811_), .B(_02060_), .Y(_02061_));
NAND_g _22407_ (.A(count_instr[7]), .B(_02058_), .Y(_02062_));
NOT_g _22408_ (.A(_02062_), .Y(_02063_));
AND_g _22409_ (.A(count_instr[7]), .B(count_instr[6]), .Y(_02064_));
AND_g _22410_ (.A(_02052_), .B(_02064_), .Y(_02065_));
AND_g _22411_ (.A(_02045_), .B(_02065_), .Y(_02066_));
AND_g _22412_ (.A(_02055_), .B(_02064_), .Y(_02067_));
AND_g _22413_ (.A(_02061_), .B(_02062_), .Y(_00593_));
NAND_g _22414_ (.A(_08785_), .B(_02062_), .Y(_02068_));
NAND_g _22415_ (.A(resetn), .B(_02068_), .Y(_02069_));
AND_g _22416_ (.A(count_instr[8]), .B(_02066_), .Y(_02070_));
NOR_g _22417_ (.A(_02069_), .B(_02070_), .Y(_00594_));
NOR_g _22418_ (.A(count_instr[9]), .B(_02070_), .Y(_02071_));
AND_g _22419_ (.A(count_instr[9]), .B(count_instr[8]), .Y(_02072_));
NOR_g _22420_ (.A(_08811_), .B(_02071_), .Y(_02073_));
AND_g _22421_ (.A(count_instr[9]), .B(_02070_), .Y(_02074_));
NAND_g _22422_ (.A(count_instr[9]), .B(_02070_), .Y(_02075_));
AND_g _22423_ (.A(_02073_), .B(_02075_), .Y(_00595_));
NOR_g _22424_ (.A(count_instr[10]), .B(_02074_), .Y(_02076_));
NOR_g _22425_ (.A(_08811_), .B(_02076_), .Y(_02077_));
NAND_g _22426_ (.A(count_instr[10]), .B(_02074_), .Y(_02078_));
AND_g _22427_ (.A(_02077_), .B(_02078_), .Y(_00596_));
NAND_g _22428_ (.A(_08784_), .B(_02078_), .Y(_02079_));
AND_g _22429_ (.A(count_instr[11]), .B(count_instr[10]), .Y(_02080_));
AND_g _22430_ (.A(_02072_), .B(_02080_), .Y(_02081_));
AND_g _22431_ (.A(_02063_), .B(_02081_), .Y(_02082_));
AND_g _22432_ (.A(resetn), .B(_02079_), .Y(_02083_));
NAND_g _22433_ (.A(_02074_), .B(_02080_), .Y(_02084_));
AND_g _22434_ (.A(_02067_), .B(_02081_), .Y(_02085_));
AND_g _22435_ (.A(_02083_), .B(_02084_), .Y(_00597_));
NAND_g _22436_ (.A(_08783_), .B(_02084_), .Y(_02086_));
AND_g _22437_ (.A(resetn), .B(_02086_), .Y(_02087_));
NAND_g _22438_ (.A(count_instr[12]), .B(_02082_), .Y(_02088_));
NOT_g _22439_ (.A(_02088_), .Y(_02089_));
AND_g _22440_ (.A(count_instr[12]), .B(_02085_), .Y(_02090_));
AND_g _22441_ (.A(_02087_), .B(_02088_), .Y(_00598_));
NAND_g _22442_ (.A(_08782_), .B(_02088_), .Y(_02091_));
AND_g _22443_ (.A(resetn), .B(_02091_), .Y(_02092_));
NAND_g _22444_ (.A(count_instr[13]), .B(_02089_), .Y(_02093_));
AND_g _22445_ (.A(count_instr[13]), .B(count_instr[12]), .Y(_02094_));
AND_g _22446_ (.A(count_instr[13]), .B(_02090_), .Y(_02095_));
AND_g _22447_ (.A(_02092_), .B(_02093_), .Y(_00599_));
NAND_g _22448_ (.A(_08781_), .B(_02093_), .Y(_02096_));
AND_g _22449_ (.A(resetn), .B(_02096_), .Y(_02097_));
NAND_g _22450_ (.A(count_instr[14]), .B(_02095_), .Y(_02098_));
AND_g _22451_ (.A(_02097_), .B(_02098_), .Y(_00600_));
NAND_g _22452_ (.A(_08780_), .B(_02098_), .Y(_02099_));
AND_g _22453_ (.A(count_instr[15]), .B(count_instr[14]), .Y(_02100_));
AND_g _22454_ (.A(_02094_), .B(_02100_), .Y(_02101_));
NAND_g _22455_ (.A(_02082_), .B(_02101_), .Y(_02102_));
AND_g _22456_ (.A(resetn), .B(_02102_), .Y(_02103_));
AND_g _22457_ (.A(_02099_), .B(_02103_), .Y(_00601_));
AND_g _22458_ (.A(_02065_), .B(_02081_), .Y(_02104_));
AND_g _22459_ (.A(_02101_), .B(_02104_), .Y(_02105_));
AND_g _22460_ (.A(_02045_), .B(_02105_), .Y(_02106_));
AND_g _22461_ (.A(_02044_), .B(_02101_), .Y(_02107_));
AND_g _22462_ (.A(_02104_), .B(_02107_), .Y(_02108_));
AND_g _22463_ (.A(_09893_), .B(_02108_), .Y(_02109_));
AND_g _22464_ (.A(count_instr[14]), .B(_02044_), .Y(_02110_));
AND_g _22465_ (.A(count_instr[13]), .B(_02052_), .Y(_02111_));
AND_g _22466_ (.A(count_instr[15]), .B(count_instr[12]), .Y(_02112_));
AND_g _22467_ (.A(_02064_), .B(_02112_), .Y(_02113_));
AND_g _22468_ (.A(_02111_), .B(_02113_), .Y(_02114_));
AND_g _22469_ (.A(_02081_), .B(_02114_), .Y(_02115_));
AND_g _22470_ (.A(_02110_), .B(_02115_), .Y(_02116_));
AND_g _22471_ (.A(_09893_), .B(_02116_), .Y(_02117_));
NOR_g _22472_ (.A(count_instr[16]), .B(_02117_), .Y(_02118_));
NOR_g _22473_ (.A(_08811_), .B(_02118_), .Y(_02119_));
NAND_g _22474_ (.A(count_instr[16]), .B(_02109_), .Y(_02120_));
AND_g _22475_ (.A(_02119_), .B(_02120_), .Y(_00602_));
NAND_g _22476_ (.A(_08779_), .B(_02120_), .Y(_02121_));
AND_g _22477_ (.A(count_instr[17]), .B(count_instr[16]), .Y(_02122_));
AND_g _22478_ (.A(_02106_), .B(_02122_), .Y(_02123_));
NAND_g _22479_ (.A(resetn), .B(_02121_), .Y(_02124_));
AND_g _22480_ (.A(_02117_), .B(_02122_), .Y(_02125_));
NOR_g _22481_ (.A(_02124_), .B(_02125_), .Y(_00603_));
NOR_g _22482_ (.A(count_instr[18]), .B(_02125_), .Y(_02126_));
NOR_g _22483_ (.A(_08811_), .B(_02126_), .Y(_02127_));
NAND_g _22484_ (.A(count_instr[18]), .B(_02123_), .Y(_02128_));
AND_g _22485_ (.A(count_instr[18]), .B(_02125_), .Y(_02129_));
AND_g _22486_ (.A(_02127_), .B(_02128_), .Y(_00604_));
NAND_g _22487_ (.A(_08778_), .B(_02128_), .Y(_02130_));
NAND_g _22488_ (.A(resetn), .B(_02130_), .Y(_02131_));
AND_g _22489_ (.A(count_instr[19]), .B(_02129_), .Y(_02132_));
NOR_g _22490_ (.A(_02131_), .B(_02132_), .Y(_00605_));
NOR_g _22491_ (.A(count_instr[20]), .B(_02132_), .Y(_02133_));
NOR_g _22492_ (.A(_08811_), .B(_02133_), .Y(_02134_));
NAND_g _22493_ (.A(count_instr[20]), .B(_02132_), .Y(_02135_));
NOT_g _22494_ (.A(_02135_), .Y(_02136_));
AND_g _22495_ (.A(_02134_), .B(_02135_), .Y(_00606_));
NOR_g _22496_ (.A(count_instr[21]), .B(_02136_), .Y(_02137_));
NOR_g _22497_ (.A(_08811_), .B(_02137_), .Y(_02138_));
NAND_g _22498_ (.A(count_instr[21]), .B(_02136_), .Y(_02139_));
AND_g _22499_ (.A(_02138_), .B(_02139_), .Y(_00607_));
NAND_g _22500_ (.A(_08777_), .B(_02139_), .Y(_02140_));
NAND_g _22501_ (.A(resetn), .B(_02140_), .Y(_02141_));
NOR_g _22502_ (.A(_08777_), .B(_02139_), .Y(_02142_));
NOR_g _22503_ (.A(_02141_), .B(_02142_), .Y(_00608_));
AND_g _22504_ (.A(count_instr[23]), .B(_02142_), .Y(_02143_));
NOR_g _22505_ (.A(count_instr[23]), .B(_02142_), .Y(_02144_));
NOT_g _22506_ (.A(_02144_), .Y(_02145_));
NAND_g _22507_ (.A(resetn), .B(_02145_), .Y(_02146_));
NOR_g _22508_ (.A(_02143_), .B(_02146_), .Y(_00609_));
NAND_g _22509_ (.A(count_instr[24]), .B(_02143_), .Y(_02147_));
NOR_g _22510_ (.A(count_instr[24]), .B(_02143_), .Y(_02148_));
NOR_g _22511_ (.A(_08811_), .B(_02148_), .Y(_02149_));
AND_g _22512_ (.A(_02147_), .B(_02149_), .Y(_00610_));
NAND_g _22513_ (.A(_08776_), .B(_02147_), .Y(_02150_));
AND_g _22514_ (.A(count_instr[25]), .B(count_instr[24]), .Y(_02151_));
AND_g _22515_ (.A(_02143_), .B(_02151_), .Y(_02152_));
NOR_g _22516_ (.A(_08811_), .B(_02152_), .Y(_02153_));
AND_g _22517_ (.A(_02150_), .B(_02153_), .Y(_00611_));
NOR_g _22518_ (.A(count_instr[26]), .B(_02152_), .Y(_02154_));
NOR_g _22519_ (.A(_08811_), .B(_02154_), .Y(_02155_));
AND_g _22520_ (.A(count_instr[26]), .B(_02152_), .Y(_02156_));
NAND_g _22521_ (.A(count_instr[26]), .B(_02152_), .Y(_02157_));
AND_g _22522_ (.A(_02155_), .B(_02157_), .Y(_00612_));
NOR_g _22523_ (.A(count_instr[27]), .B(_02156_), .Y(_02158_));
NOR_g _22524_ (.A(_08811_), .B(_02158_), .Y(_02159_));
NAND_g _22525_ (.A(count_instr[27]), .B(_02156_), .Y(_02160_));
AND_g _22526_ (.A(_02159_), .B(_02160_), .Y(_00613_));
NAND_g _22527_ (.A(_08775_), .B(_02160_), .Y(_02161_));
NAND_g _22528_ (.A(resetn), .B(_02161_), .Y(_02162_));
NOR_g _22529_ (.A(_08775_), .B(_02160_), .Y(_02163_));
NOR_g _22530_ (.A(_02162_), .B(_02163_), .Y(_00614_));
NOR_g _22531_ (.A(count_instr[29]), .B(_02163_), .Y(_02164_));
NOR_g _22532_ (.A(_08811_), .B(_02164_), .Y(_02165_));
NAND_g _22533_ (.A(count_instr[29]), .B(_02163_), .Y(_02166_));
AND_g _22534_ (.A(_02165_), .B(_02166_), .Y(_00615_));
NAND_g _22535_ (.A(_08774_), .B(_02166_), .Y(_02167_));
NAND_g _22536_ (.A(resetn), .B(_02167_), .Y(_02168_));
NOR_g _22537_ (.A(_08774_), .B(_02166_), .Y(_02169_));
NOR_g _22538_ (.A(_02168_), .B(_02169_), .Y(_00616_));
AND_g _22539_ (.A(count_instr[31]), .B(_02169_), .Y(_02170_));
NOR_g _22540_ (.A(count_instr[31]), .B(_02169_), .Y(_02171_));
NOT_g _22541_ (.A(_02171_), .Y(_02172_));
NAND_g _22542_ (.A(resetn), .B(_02172_), .Y(_02173_));
NOR_g _22543_ (.A(_02170_), .B(_02173_), .Y(_00617_));
AND_g _22544_ (.A(count_instr[32]), .B(_02170_), .Y(_02174_));
NOR_g _22545_ (.A(count_instr[32]), .B(_02170_), .Y(_02175_));
NOT_g _22546_ (.A(_02175_), .Y(_02176_));
NAND_g _22547_ (.A(resetn), .B(_02176_), .Y(_02177_));
NOR_g _22548_ (.A(_02174_), .B(_02177_), .Y(_00618_));
NOR_g _22549_ (.A(count_instr[33]), .B(_02174_), .Y(_02178_));
NOT_g _22550_ (.A(_02178_), .Y(_02179_));
AND_g _22551_ (.A(count_instr[33]), .B(_02174_), .Y(_02180_));
NOR_g _22552_ (.A(_08811_), .B(_02180_), .Y(_02181_));
AND_g _22553_ (.A(_02179_), .B(_02181_), .Y(_00619_));
NAND_g _22554_ (.A(count_instr[34]), .B(_02180_), .Y(_02182_));
NOR_g _22555_ (.A(count_instr[34]), .B(_02180_), .Y(_02183_));
NOR_g _22556_ (.A(_08811_), .B(_02183_), .Y(_02184_));
AND_g _22557_ (.A(_02182_), .B(_02184_), .Y(_00620_));
NAND_g _22558_ (.A(_08773_), .B(_02182_), .Y(_02185_));
NAND_g _22559_ (.A(resetn), .B(_02185_), .Y(_02186_));
NOR_g _22560_ (.A(_08773_), .B(_02182_), .Y(_02187_));
AND_g _22561_ (.A(count_instr[35]), .B(count_instr[34]), .Y(_02188_));
NOR_g _22562_ (.A(_02186_), .B(_02187_), .Y(_00621_));
NOR_g _22563_ (.A(count_instr[36]), .B(_02187_), .Y(_02189_));
NOR_g _22564_ (.A(_08811_), .B(_02189_), .Y(_02190_));
NAND_g _22565_ (.A(count_instr[36]), .B(_02187_), .Y(_02191_));
AND_g _22566_ (.A(_02190_), .B(_02191_), .Y(_00622_));
NAND_g _22567_ (.A(_08772_), .B(_02191_), .Y(_02192_));
AND_g _22568_ (.A(count_instr[37]), .B(count_instr[36]), .Y(_02193_));
AND_g _22569_ (.A(_02188_), .B(_02193_), .Y(_02194_));
AND_g _22570_ (.A(_02180_), .B(_02194_), .Y(_02195_));
NOR_g _22571_ (.A(_08811_), .B(_02195_), .Y(_02196_));
AND_g _22572_ (.A(_02192_), .B(_02196_), .Y(_00623_));
NOR_g _22573_ (.A(count_instr[38]), .B(_02195_), .Y(_02197_));
NOR_g _22574_ (.A(_08811_), .B(_02197_), .Y(_02198_));
NAND_g _22575_ (.A(count_instr[38]), .B(_02195_), .Y(_02199_));
AND_g _22576_ (.A(_02198_), .B(_02199_), .Y(_00624_));
XNOR_g _22577_ (.A(count_instr[39]), .B(_02199_), .Y(_02200_));
NOR_g _22578_ (.A(_08771_), .B(_02199_), .Y(_02201_));
AND_g _22579_ (.A(resetn), .B(_02200_), .Y(_00625_));
NAND_g _22580_ (.A(count_instr[40]), .B(_02201_), .Y(_02202_));
NOR_g _22581_ (.A(count_instr[40]), .B(_02201_), .Y(_02203_));
NOR_g _22582_ (.A(_08811_), .B(_02203_), .Y(_02204_));
AND_g _22583_ (.A(_02202_), .B(_02204_), .Y(_00626_));
AND_g _22584_ (.A(count_instr[41]), .B(count_instr[40]), .Y(_02205_));
AND_g _22585_ (.A(_02201_), .B(_02205_), .Y(_02206_));
NAND_g _22586_ (.A(_08770_), .B(_02202_), .Y(_02207_));
NAND_g _22587_ (.A(resetn), .B(_02207_), .Y(_02208_));
NOR_g _22588_ (.A(_02206_), .B(_02208_), .Y(_00627_));
AND_g _22589_ (.A(count_instr[42]), .B(_02206_), .Y(_02209_));
NOR_g _22590_ (.A(count_instr[42]), .B(_02206_), .Y(_02210_));
NOT_g _22591_ (.A(_02210_), .Y(_02211_));
NAND_g _22592_ (.A(resetn), .B(_02211_), .Y(_02212_));
NOR_g _22593_ (.A(_02209_), .B(_02212_), .Y(_00628_));
NOR_g _22594_ (.A(count_instr[43]), .B(_02209_), .Y(_02213_));
AND_g _22595_ (.A(count_instr[43]), .B(count_instr[42]), .Y(_02214_));
AND_g _22596_ (.A(_02206_), .B(_02214_), .Y(_02215_));
NAND_g _22597_ (.A(_02206_), .B(_02214_), .Y(_02216_));
NAND_g _22598_ (.A(resetn), .B(_02216_), .Y(_02217_));
AND_g _22599_ (.A(count_instr[43]), .B(_02209_), .Y(_02218_));
NOR_g _22600_ (.A(_02213_), .B(_02217_), .Y(_00629_));
AND_g _22601_ (.A(_02205_), .B(_02214_), .Y(_02219_));
AND_g _22602_ (.A(_02201_), .B(_02219_), .Y(_02220_));
NOR_g _22603_ (.A(count_instr[44]), .B(_02220_), .Y(_02221_));
NOR_g _22604_ (.A(_08811_), .B(_02221_), .Y(_02222_));
NAND_g _22605_ (.A(count_instr[44]), .B(_02215_), .Y(_02223_));
AND_g _22606_ (.A(count_instr[44]), .B(_02220_), .Y(_02224_));
AND_g _22607_ (.A(_02222_), .B(_02223_), .Y(_00630_));
NAND_g _22608_ (.A(_08769_), .B(_02223_), .Y(_02225_));
AND_g _22609_ (.A(resetn), .B(_02225_), .Y(_02226_));
AND_g _22610_ (.A(count_instr[45]), .B(count_instr[44]), .Y(_02227_));
NAND_g _22611_ (.A(_02218_), .B(_02227_), .Y(_02228_));
AND_g _22612_ (.A(count_instr[45]), .B(_02224_), .Y(_02229_));
AND_g _22613_ (.A(_02226_), .B(_02228_), .Y(_00631_));
NAND_g _22614_ (.A(_08768_), .B(_02228_), .Y(_02230_));
AND_g _22615_ (.A(resetn), .B(_02230_), .Y(_02231_));
NAND_g _22616_ (.A(count_instr[46]), .B(_02229_), .Y(_02232_));
AND_g _22617_ (.A(_02231_), .B(_02232_), .Y(_00632_));
NAND_g _22618_ (.A(_08767_), .B(_02232_), .Y(_02233_));
AND_g _22619_ (.A(count_instr[47]), .B(count_instr[46]), .Y(_02234_));
AND_g _22620_ (.A(_02227_), .B(_02234_), .Y(_02235_));
NAND_g _22621_ (.A(_02215_), .B(_02235_), .Y(_02236_));
AND_g _22622_ (.A(resetn), .B(_02236_), .Y(_02237_));
AND_g _22623_ (.A(_02233_), .B(_02237_), .Y(_00633_));
AND_g _22624_ (.A(_02219_), .B(_02235_), .Y(_02238_));
AND_g _22625_ (.A(_02201_), .B(_02238_), .Y(_02239_));
NAND_g _22626_ (.A(count_instr[48]), .B(_02239_), .Y(_02240_));
NOR_g _22627_ (.A(count_instr[48]), .B(_02239_), .Y(_02241_));
NOR_g _22628_ (.A(_08811_), .B(_02241_), .Y(_02242_));
AND_g _22629_ (.A(_02240_), .B(_02242_), .Y(_00634_));
NAND_g _22630_ (.A(_08766_), .B(_02240_), .Y(_02243_));
AND_g _22631_ (.A(count_instr[49]), .B(count_instr[48]), .Y(_02244_));
AND_g _22632_ (.A(_02239_), .B(_02244_), .Y(_02245_));
NOR_g _22633_ (.A(_08811_), .B(_02245_), .Y(_02246_));
AND_g _22634_ (.A(_02243_), .B(_02246_), .Y(_00635_));
NOR_g _22635_ (.A(count_instr[50]), .B(_02245_), .Y(_02247_));
NOR_g _22636_ (.A(_08811_), .B(_02247_), .Y(_02248_));
AND_g _22637_ (.A(count_instr[50]), .B(_02245_), .Y(_02249_));
NAND_g _22638_ (.A(count_instr[50]), .B(_02245_), .Y(_02250_));
AND_g _22639_ (.A(_02248_), .B(_02250_), .Y(_00636_));
NOR_g _22640_ (.A(count_instr[51]), .B(_02249_), .Y(_02251_));
NOR_g _22641_ (.A(_08811_), .B(_02251_), .Y(_02252_));
NAND_g _22642_ (.A(count_instr[51]), .B(_02249_), .Y(_02253_));
AND_g _22643_ (.A(count_instr[51]), .B(count_instr[50]), .Y(_02254_));
AND_g _22644_ (.A(_02252_), .B(_02253_), .Y(_00637_));
NAND_g _22645_ (.A(_08765_), .B(_02253_), .Y(_02255_));
NAND_g _22646_ (.A(resetn), .B(_02255_), .Y(_02256_));
NOR_g _22647_ (.A(_08765_), .B(_02253_), .Y(_02257_));
NOR_g _22648_ (.A(_02256_), .B(_02257_), .Y(_00638_));
NOR_g _22649_ (.A(count_instr[53]), .B(_02257_), .Y(_02258_));
AND_g _22650_ (.A(count_instr[53]), .B(count_instr[52]), .Y(_02259_));
AND_g _22651_ (.A(_02254_), .B(_02259_), .Y(_02260_));
AND_g _22652_ (.A(_02245_), .B(_02260_), .Y(_02261_));
NOR_g _22653_ (.A(_08811_), .B(_02258_), .Y(_02262_));
NAND_g _22654_ (.A(count_instr[53]), .B(_02257_), .Y(_02263_));
AND_g _22655_ (.A(_02262_), .B(_02263_), .Y(_00639_));
NAND_g _22656_ (.A(_08764_), .B(_02263_), .Y(_02264_));
AND_g _22657_ (.A(resetn), .B(_02264_), .Y(_02265_));
NAND_g _22658_ (.A(count_instr[54]), .B(_02261_), .Y(_02266_));
AND_g _22659_ (.A(_02265_), .B(_02266_), .Y(_00640_));
XNOR_g _22660_ (.A(count_instr[55]), .B(_02266_), .Y(_02267_));
AND_g _22661_ (.A(resetn), .B(_02267_), .Y(_00641_));
AND_g _22662_ (.A(count_instr[55]), .B(count_instr[54]), .Y(_02268_));
AND_g _22663_ (.A(_02244_), .B(_02268_), .Y(_02269_));
AND_g _22664_ (.A(_02260_), .B(_02269_), .Y(_02270_));
AND_g _22665_ (.A(_02239_), .B(_02270_), .Y(_02271_));
NOR_g _22666_ (.A(count_instr[56]), .B(_02271_), .Y(_02272_));
NOR_g _22667_ (.A(_08811_), .B(_02272_), .Y(_02273_));
AND_g _22668_ (.A(count_instr[56]), .B(_02271_), .Y(_02274_));
NAND_g _22669_ (.A(count_instr[56]), .B(_02271_), .Y(_02275_));
AND_g _22670_ (.A(_02273_), .B(_02275_), .Y(_00642_));
NOR_g _22671_ (.A(count_instr[57]), .B(_02274_), .Y(_02276_));
NOR_g _22672_ (.A(_08811_), .B(_02276_), .Y(_02277_));
NAND_g _22673_ (.A(count_instr[57]), .B(_02274_), .Y(_02278_));
AND_g _22674_ (.A(_02277_), .B(_02278_), .Y(_00643_));
NAND_g _22675_ (.A(_08763_), .B(_02278_), .Y(_02279_));
NAND_g _22676_ (.A(resetn), .B(_02279_), .Y(_02280_));
NOR_g _22677_ (.A(_08763_), .B(_02278_), .Y(_02281_));
NOR_g _22678_ (.A(_02280_), .B(_02281_), .Y(_00644_));
NOR_g _22679_ (.A(count_instr[59]), .B(_02281_), .Y(_02282_));
NOR_g _22680_ (.A(_08811_), .B(_02282_), .Y(_02283_));
NAND_g _22681_ (.A(count_instr[59]), .B(_02281_), .Y(_02284_));
AND_g _22682_ (.A(_02283_), .B(_02284_), .Y(_00645_));
NAND_g _22683_ (.A(_08762_), .B(_02284_), .Y(_02285_));
NAND_g _22684_ (.A(resetn), .B(_02285_), .Y(_02286_));
NOR_g _22685_ (.A(_08762_), .B(_02284_), .Y(_02287_));
NOR_g _22686_ (.A(_02286_), .B(_02287_), .Y(_00646_));
NOR_g _22687_ (.A(count_instr[61]), .B(_02287_), .Y(_02288_));
NOR_g _22688_ (.A(_08811_), .B(_02288_), .Y(_02289_));
NAND_g _22689_ (.A(count_instr[61]), .B(_02287_), .Y(_02290_));
NOT_g _22690_ (.A(_02290_), .Y(_02291_));
AND_g _22691_ (.A(_02289_), .B(_02290_), .Y(_00647_));
NAND_g _22692_ (.A(_08761_), .B(_02290_), .Y(_02292_));
AND_g _22693_ (.A(resetn), .B(_02292_), .Y(_02293_));
NAND_g _22694_ (.A(count_instr[62]), .B(_02291_), .Y(_02294_));
AND_g _22695_ (.A(_02293_), .B(_02294_), .Y(_00648_));
XNOR_g _22696_ (.A(count_instr[63]), .B(_02294_), .Y(_02295_));
AND_g _22697_ (.A(resetn), .B(_02295_), .Y(_00649_));
AND_g _22698_ (.A(_09087_), .B(_14286_), .Y(_02296_));
NAND_g _22699_ (.A(_09087_), .B(_14286_), .Y(_02297_));
NAND_g _22700_ (.A(_09098_), .B(_02296_), .Y(_02298_));
NAND_g _22701_ (.A(cpuregs[12][0]), .B(_02297_), .Y(_02299_));
NAND_g _22702_ (.A(_02298_), .B(_02299_), .Y(_00650_));
NAND_g _22703_ (.A(_09109_), .B(_02296_), .Y(_02300_));
NAND_g _22704_ (.A(cpuregs[12][1]), .B(_02297_), .Y(_02301_));
NAND_g _22705_ (.A(_02300_), .B(_02301_), .Y(_00651_));
NAND_g _22706_ (.A(cpuregs[12][2]), .B(_02297_), .Y(_02302_));
NAND_g _22707_ (.A(_09118_), .B(_02296_), .Y(_02303_));
NAND_g _22708_ (.A(_02302_), .B(_02303_), .Y(_00652_));
NAND_g _22709_ (.A(cpuregs[12][3]), .B(_02297_), .Y(_02304_));
NAND_g _22710_ (.A(_09131_), .B(_02296_), .Y(_02305_));
NAND_g _22711_ (.A(_02304_), .B(_02305_), .Y(_00653_));
NAND_g _22712_ (.A(cpuregs[12][4]), .B(_02297_), .Y(_02306_));
NAND_g _22713_ (.A(_09144_), .B(_02296_), .Y(_02307_));
NAND_g _22714_ (.A(_02306_), .B(_02307_), .Y(_00654_));
NAND_g _22715_ (.A(cpuregs[12][5]), .B(_02297_), .Y(_02308_));
NAND_g _22716_ (.A(_09157_), .B(_02296_), .Y(_02309_));
NAND_g _22717_ (.A(_02308_), .B(_02309_), .Y(_00655_));
NAND_g _22718_ (.A(cpuregs[12][6]), .B(_02297_), .Y(_02310_));
NAND_g _22719_ (.A(_09170_), .B(_02296_), .Y(_02311_));
NAND_g _22720_ (.A(_02310_), .B(_02311_), .Y(_00656_));
NAND_g _22721_ (.A(cpuregs[12][7]), .B(_02297_), .Y(_02312_));
NAND_g _22722_ (.A(_09183_), .B(_02296_), .Y(_02313_));
NAND_g _22723_ (.A(_02312_), .B(_02313_), .Y(_00657_));
NAND_g _22724_ (.A(cpuregs[12][8]), .B(_02297_), .Y(_02314_));
NAND_g _22725_ (.A(_09196_), .B(_02296_), .Y(_02315_));
NAND_g _22726_ (.A(_02314_), .B(_02315_), .Y(_00658_));
NAND_g _22727_ (.A(cpuregs[12][9]), .B(_02297_), .Y(_02316_));
NAND_g _22728_ (.A(_09209_), .B(_02296_), .Y(_02317_));
NAND_g _22729_ (.A(_02316_), .B(_02317_), .Y(_00659_));
NAND_g _22730_ (.A(cpuregs[12][10]), .B(_02297_), .Y(_02318_));
NAND_g _22731_ (.A(_09222_), .B(_02296_), .Y(_02319_));
NAND_g _22732_ (.A(_02318_), .B(_02319_), .Y(_00660_));
NAND_g _22733_ (.A(cpuregs[12][11]), .B(_02297_), .Y(_02320_));
NAND_g _22734_ (.A(_09235_), .B(_02296_), .Y(_02321_));
NAND_g _22735_ (.A(_02320_), .B(_02321_), .Y(_00661_));
NAND_g _22736_ (.A(_09248_), .B(_02296_), .Y(_02322_));
NAND_g _22737_ (.A(cpuregs[12][12]), .B(_02297_), .Y(_02323_));
NAND_g _22738_ (.A(_02322_), .B(_02323_), .Y(_00662_));
NAND_g _22739_ (.A(cpuregs[12][13]), .B(_02297_), .Y(_02324_));
NAND_g _22740_ (.A(_09261_), .B(_02296_), .Y(_02325_));
NAND_g _22741_ (.A(_02324_), .B(_02325_), .Y(_00663_));
NAND_g _22742_ (.A(cpuregs[12][14]), .B(_02297_), .Y(_02326_));
NAND_g _22743_ (.A(_09274_), .B(_02296_), .Y(_02327_));
NAND_g _22744_ (.A(_02326_), .B(_02327_), .Y(_00664_));
NAND_g _22745_ (.A(cpuregs[12][15]), .B(_02297_), .Y(_02328_));
NAND_g _22746_ (.A(_09287_), .B(_02296_), .Y(_02329_));
NAND_g _22747_ (.A(_02328_), .B(_02329_), .Y(_00665_));
NOR_g _22748_ (.A(cpuregs[12][16]), .B(_02296_), .Y(_02330_));
NOR_g _22749_ (.A(_09300_), .B(_02297_), .Y(_02331_));
NOR_g _22750_ (.A(_02330_), .B(_02331_), .Y(_00666_));
NOR_g _22751_ (.A(cpuregs[12][17]), .B(_02296_), .Y(_02332_));
NOR_g _22752_ (.A(_09313_), .B(_02297_), .Y(_02333_));
NOR_g _22753_ (.A(_02332_), .B(_02333_), .Y(_00667_));
NAND_g _22754_ (.A(cpuregs[12][18]), .B(_02297_), .Y(_02334_));
NAND_g _22755_ (.A(_09325_), .B(_02296_), .Y(_02335_));
NAND_g _22756_ (.A(_02334_), .B(_02335_), .Y(_00668_));
NAND_g _22757_ (.A(cpuregs[12][19]), .B(_02297_), .Y(_02336_));
NAND_g _22758_ (.A(_09338_), .B(_02296_), .Y(_02337_));
NAND_g _22759_ (.A(_02336_), .B(_02337_), .Y(_00669_));
NAND_g _22760_ (.A(cpuregs[12][20]), .B(_02297_), .Y(_02338_));
NAND_g _22761_ (.A(_09351_), .B(_02296_), .Y(_02339_));
NAND_g _22762_ (.A(_02338_), .B(_02339_), .Y(_00670_));
NAND_g _22763_ (.A(_09364_), .B(_02296_), .Y(_02340_));
NAND_g _22764_ (.A(cpuregs[12][21]), .B(_02297_), .Y(_02341_));
NAND_g _22765_ (.A(_02340_), .B(_02341_), .Y(_00671_));
NAND_g _22766_ (.A(_09377_), .B(_02296_), .Y(_02342_));
NAND_g _22767_ (.A(cpuregs[12][22]), .B(_02297_), .Y(_02343_));
NAND_g _22768_ (.A(_02342_), .B(_02343_), .Y(_00672_));
NAND_g _22769_ (.A(cpuregs[12][23]), .B(_02297_), .Y(_02344_));
NAND_g _22770_ (.A(_09390_), .B(_02296_), .Y(_02345_));
NAND_g _22771_ (.A(_02344_), .B(_02345_), .Y(_00673_));
NAND_g _22772_ (.A(_09403_), .B(_02296_), .Y(_02346_));
NAND_g _22773_ (.A(cpuregs[12][24]), .B(_02297_), .Y(_02347_));
NAND_g _22774_ (.A(_02346_), .B(_02347_), .Y(_00674_));
NAND_g _22775_ (.A(cpuregs[12][25]), .B(_02297_), .Y(_02348_));
NAND_g _22776_ (.A(_09416_), .B(_02296_), .Y(_02349_));
NAND_g _22777_ (.A(_02348_), .B(_02349_), .Y(_00675_));
NAND_g _22778_ (.A(cpuregs[12][26]), .B(_02297_), .Y(_02350_));
NAND_g _22779_ (.A(_09429_), .B(_02296_), .Y(_02351_));
NAND_g _22780_ (.A(_02350_), .B(_02351_), .Y(_00676_));
NAND_g _22781_ (.A(cpuregs[12][27]), .B(_02297_), .Y(_02352_));
NAND_g _22782_ (.A(_09442_), .B(_02296_), .Y(_02353_));
NAND_g _22783_ (.A(_02352_), .B(_02353_), .Y(_00677_));
NAND_g _22784_ (.A(cpuregs[12][28]), .B(_02297_), .Y(_02354_));
NAND_g _22785_ (.A(_09455_), .B(_02296_), .Y(_02355_));
NAND_g _22786_ (.A(_02354_), .B(_02355_), .Y(_00678_));
NAND_g _22787_ (.A(cpuregs[12][29]), .B(_02297_), .Y(_02356_));
NAND_g _22788_ (.A(_09468_), .B(_02296_), .Y(_02357_));
NAND_g _22789_ (.A(_02356_), .B(_02357_), .Y(_00679_));
NAND_g _22790_ (.A(cpuregs[12][30]), .B(_02297_), .Y(_02358_));
NAND_g _22791_ (.A(_09481_), .B(_02296_), .Y(_02359_));
NAND_g _22792_ (.A(_02358_), .B(_02359_), .Y(_00680_));
NAND_g _22793_ (.A(_09493_), .B(_02296_), .Y(_02360_));
NAND_g _22794_ (.A(cpuregs[12][31]), .B(_02297_), .Y(_02361_));
NAND_g _22795_ (.A(_02360_), .B(_02361_), .Y(_00681_));
AND_g _22796_ (.A(_09085_), .B(_09567_), .Y(_02362_));
NAND_g _22797_ (.A(_09085_), .B(_09567_), .Y(_02363_));
NAND_g _22798_ (.A(_09098_), .B(_02362_), .Y(_02364_));
NAND_g _22799_ (.A(cpuregs[3][0]), .B(_02363_), .Y(_02365_));
NAND_g _22800_ (.A(_02364_), .B(_02365_), .Y(_00682_));
NAND_g _22801_ (.A(_09109_), .B(_02362_), .Y(_02366_));
NAND_g _22802_ (.A(cpuregs[3][1]), .B(_02363_), .Y(_02367_));
NAND_g _22803_ (.A(_02366_), .B(_02367_), .Y(_00683_));
NAND_g _22804_ (.A(_09118_), .B(_02362_), .Y(_02368_));
NAND_g _22805_ (.A(cpuregs[3][2]), .B(_02363_), .Y(_02369_));
NAND_g _22806_ (.A(_02368_), .B(_02369_), .Y(_00684_));
NAND_g _22807_ (.A(_09131_), .B(_02362_), .Y(_02370_));
NAND_g _22808_ (.A(cpuregs[3][3]), .B(_02363_), .Y(_02371_));
NAND_g _22809_ (.A(_02370_), .B(_02371_), .Y(_00685_));
NAND_g _22810_ (.A(_09144_), .B(_02362_), .Y(_02372_));
NAND_g _22811_ (.A(cpuregs[3][4]), .B(_02363_), .Y(_02373_));
NAND_g _22812_ (.A(_02372_), .B(_02373_), .Y(_00686_));
NAND_g _22813_ (.A(_09157_), .B(_02362_), .Y(_02374_));
NAND_g _22814_ (.A(cpuregs[3][5]), .B(_02363_), .Y(_02375_));
NAND_g _22815_ (.A(_02374_), .B(_02375_), .Y(_00687_));
NAND_g _22816_ (.A(_09170_), .B(_02362_), .Y(_02376_));
NAND_g _22817_ (.A(cpuregs[3][6]), .B(_02363_), .Y(_02377_));
NAND_g _22818_ (.A(_02376_), .B(_02377_), .Y(_00688_));
NAND_g _22819_ (.A(_09183_), .B(_02362_), .Y(_02378_));
NAND_g _22820_ (.A(cpuregs[3][7]), .B(_02363_), .Y(_02379_));
NAND_g _22821_ (.A(_02378_), .B(_02379_), .Y(_00689_));
NAND_g _22822_ (.A(_09196_), .B(_02362_), .Y(_02380_));
NAND_g _22823_ (.A(cpuregs[3][8]), .B(_02363_), .Y(_02381_));
NAND_g _22824_ (.A(_02380_), .B(_02381_), .Y(_00690_));
NAND_g _22825_ (.A(_09209_), .B(_02362_), .Y(_02382_));
NAND_g _22826_ (.A(cpuregs[3][9]), .B(_02363_), .Y(_02383_));
NAND_g _22827_ (.A(_02382_), .B(_02383_), .Y(_00691_));
NAND_g _22828_ (.A(_09222_), .B(_02362_), .Y(_02384_));
NAND_g _22829_ (.A(cpuregs[3][10]), .B(_02363_), .Y(_02385_));
NAND_g _22830_ (.A(_02384_), .B(_02385_), .Y(_00692_));
NAND_g _22831_ (.A(_09235_), .B(_02362_), .Y(_02386_));
NAND_g _22832_ (.A(cpuregs[3][11]), .B(_02363_), .Y(_02387_));
NAND_g _22833_ (.A(_02386_), .B(_02387_), .Y(_00693_));
NAND_g _22834_ (.A(_09248_), .B(_02362_), .Y(_02388_));
NAND_g _22835_ (.A(cpuregs[3][12]), .B(_02363_), .Y(_02389_));
NAND_g _22836_ (.A(_02388_), .B(_02389_), .Y(_00694_));
NAND_g _22837_ (.A(_09261_), .B(_02362_), .Y(_02390_));
NAND_g _22838_ (.A(cpuregs[3][13]), .B(_02363_), .Y(_02391_));
NAND_g _22839_ (.A(_02390_), .B(_02391_), .Y(_00695_));
NAND_g _22840_ (.A(_09274_), .B(_02362_), .Y(_02392_));
NAND_g _22841_ (.A(cpuregs[3][14]), .B(_02363_), .Y(_02393_));
NAND_g _22842_ (.A(_02392_), .B(_02393_), .Y(_00696_));
NAND_g _22843_ (.A(_09287_), .B(_02362_), .Y(_02394_));
NAND_g _22844_ (.A(cpuregs[3][15]), .B(_02363_), .Y(_02395_));
NAND_g _22845_ (.A(_02394_), .B(_02395_), .Y(_00697_));
NAND_g _22846_ (.A(_09300_), .B(_02362_), .Y(_02396_));
NAND_g _22847_ (.A(cpuregs[3][16]), .B(_02363_), .Y(_02397_));
NAND_g _22848_ (.A(_02396_), .B(_02397_), .Y(_00698_));
NOR_g _22849_ (.A(cpuregs[3][17]), .B(_02362_), .Y(_02398_));
NOR_g _22850_ (.A(_09313_), .B(_02363_), .Y(_02399_));
NOR_g _22851_ (.A(_02398_), .B(_02399_), .Y(_00699_));
NOR_g _22852_ (.A(cpuregs[3][18]), .B(_02362_), .Y(_02400_));
NOR_g _22853_ (.A(_09325_), .B(_02363_), .Y(_02401_));
NOR_g _22854_ (.A(_02400_), .B(_02401_), .Y(_00700_));
NAND_g _22855_ (.A(_09338_), .B(_02362_), .Y(_02402_));
NAND_g _22856_ (.A(cpuregs[3][19]), .B(_02363_), .Y(_02403_));
NAND_g _22857_ (.A(_02402_), .B(_02403_), .Y(_00701_));
NAND_g _22858_ (.A(_09351_), .B(_02362_), .Y(_02404_));
NAND_g _22859_ (.A(cpuregs[3][20]), .B(_02363_), .Y(_02405_));
NAND_g _22860_ (.A(_02404_), .B(_02405_), .Y(_00702_));
NAND_g _22861_ (.A(_09364_), .B(_02362_), .Y(_02406_));
NAND_g _22862_ (.A(cpuregs[3][21]), .B(_02363_), .Y(_02407_));
NAND_g _22863_ (.A(_02406_), .B(_02407_), .Y(_00703_));
NAND_g _22864_ (.A(_09377_), .B(_02362_), .Y(_02408_));
NAND_g _22865_ (.A(cpuregs[3][22]), .B(_02363_), .Y(_02409_));
NAND_g _22866_ (.A(_02408_), .B(_02409_), .Y(_00704_));
NAND_g _22867_ (.A(_09390_), .B(_02362_), .Y(_02410_));
NAND_g _22868_ (.A(cpuregs[3][23]), .B(_02363_), .Y(_02411_));
NAND_g _22869_ (.A(_02410_), .B(_02411_), .Y(_00705_));
NAND_g _22870_ (.A(_09403_), .B(_02362_), .Y(_02412_));
NAND_g _22871_ (.A(cpuregs[3][24]), .B(_02363_), .Y(_02413_));
NAND_g _22872_ (.A(_02412_), .B(_02413_), .Y(_00706_));
NAND_g _22873_ (.A(_09416_), .B(_02362_), .Y(_02414_));
NAND_g _22874_ (.A(cpuregs[3][25]), .B(_02363_), .Y(_02415_));
NAND_g _22875_ (.A(_02414_), .B(_02415_), .Y(_00707_));
NAND_g _22876_ (.A(_09429_), .B(_02362_), .Y(_02416_));
NAND_g _22877_ (.A(cpuregs[3][26]), .B(_02363_), .Y(_02417_));
NAND_g _22878_ (.A(_02416_), .B(_02417_), .Y(_00708_));
NAND_g _22879_ (.A(_09442_), .B(_02362_), .Y(_02418_));
NAND_g _22880_ (.A(cpuregs[3][27]), .B(_02363_), .Y(_02419_));
NAND_g _22881_ (.A(_02418_), .B(_02419_), .Y(_00709_));
NAND_g _22882_ (.A(_09455_), .B(_02362_), .Y(_02420_));
NAND_g _22883_ (.A(cpuregs[3][28]), .B(_02363_), .Y(_02421_));
NAND_g _22884_ (.A(_02420_), .B(_02421_), .Y(_00710_));
NAND_g _22885_ (.A(_09468_), .B(_02362_), .Y(_02422_));
NAND_g _22886_ (.A(cpuregs[3][29]), .B(_02363_), .Y(_02423_));
NAND_g _22887_ (.A(_02422_), .B(_02423_), .Y(_00711_));
NAND_g _22888_ (.A(_09481_), .B(_02362_), .Y(_02424_));
NAND_g _22889_ (.A(cpuregs[3][30]), .B(_02363_), .Y(_02425_));
NAND_g _22890_ (.A(_02424_), .B(_02425_), .Y(_00712_));
NAND_g _22891_ (.A(_09493_), .B(_02362_), .Y(_02426_));
NAND_g _22892_ (.A(cpuregs[3][31]), .B(_02363_), .Y(_02427_));
NAND_g _22893_ (.A(_02426_), .B(_02427_), .Y(_00713_));
AND_g _22894_ (.A(_09085_), .B(_14285_), .Y(_02428_));
NAND_g _22895_ (.A(_09085_), .B(_14285_), .Y(_02429_));
NAND_g _22896_ (.A(_09098_), .B(_02428_), .Y(_02430_));
NAND_g _22897_ (.A(cpuregs[23][0]), .B(_02429_), .Y(_02431_));
NAND_g _22898_ (.A(_02430_), .B(_02431_), .Y(_00714_));
NAND_g _22899_ (.A(_09109_), .B(_02428_), .Y(_02432_));
NAND_g _22900_ (.A(cpuregs[23][1]), .B(_02429_), .Y(_02433_));
NAND_g _22901_ (.A(_02432_), .B(_02433_), .Y(_00715_));
NAND_g _22902_ (.A(_09118_), .B(_02428_), .Y(_02434_));
NAND_g _22903_ (.A(cpuregs[23][2]), .B(_02429_), .Y(_02435_));
NAND_g _22904_ (.A(_02434_), .B(_02435_), .Y(_00716_));
NAND_g _22905_ (.A(_09131_), .B(_02428_), .Y(_02436_));
NAND_g _22906_ (.A(cpuregs[23][3]), .B(_02429_), .Y(_02437_));
NAND_g _22907_ (.A(_02436_), .B(_02437_), .Y(_00717_));
NAND_g _22908_ (.A(_09144_), .B(_02428_), .Y(_02438_));
NAND_g _22909_ (.A(cpuregs[23][4]), .B(_02429_), .Y(_02439_));
NAND_g _22910_ (.A(_02438_), .B(_02439_), .Y(_00718_));
NAND_g _22911_ (.A(_09157_), .B(_02428_), .Y(_02440_));
NAND_g _22912_ (.A(cpuregs[23][5]), .B(_02429_), .Y(_02441_));
NAND_g _22913_ (.A(_02440_), .B(_02441_), .Y(_00719_));
NAND_g _22914_ (.A(_09170_), .B(_02428_), .Y(_02442_));
NAND_g _22915_ (.A(cpuregs[23][6]), .B(_02429_), .Y(_02443_));
NAND_g _22916_ (.A(_02442_), .B(_02443_), .Y(_00720_));
NAND_g _22917_ (.A(_09183_), .B(_02428_), .Y(_02444_));
NAND_g _22918_ (.A(cpuregs[23][7]), .B(_02429_), .Y(_02445_));
NAND_g _22919_ (.A(_02444_), .B(_02445_), .Y(_00721_));
NAND_g _22920_ (.A(_09196_), .B(_02428_), .Y(_02446_));
NAND_g _22921_ (.A(cpuregs[23][8]), .B(_02429_), .Y(_02447_));
NAND_g _22922_ (.A(_02446_), .B(_02447_), .Y(_00722_));
NAND_g _22923_ (.A(_09209_), .B(_02428_), .Y(_02448_));
NAND_g _22924_ (.A(cpuregs[23][9]), .B(_02429_), .Y(_02449_));
NAND_g _22925_ (.A(_02448_), .B(_02449_), .Y(_00723_));
NAND_g _22926_ (.A(_09222_), .B(_02428_), .Y(_02450_));
NAND_g _22927_ (.A(cpuregs[23][10]), .B(_02429_), .Y(_02451_));
NAND_g _22928_ (.A(_02450_), .B(_02451_), .Y(_00724_));
NAND_g _22929_ (.A(_09235_), .B(_02428_), .Y(_02452_));
NAND_g _22930_ (.A(cpuregs[23][11]), .B(_02429_), .Y(_02453_));
NAND_g _22931_ (.A(_02452_), .B(_02453_), .Y(_00725_));
NAND_g _22932_ (.A(_09248_), .B(_02428_), .Y(_02454_));
NAND_g _22933_ (.A(cpuregs[23][12]), .B(_02429_), .Y(_02455_));
NAND_g _22934_ (.A(_02454_), .B(_02455_), .Y(_00726_));
NAND_g _22935_ (.A(_09261_), .B(_02428_), .Y(_02456_));
NAND_g _22936_ (.A(cpuregs[23][13]), .B(_02429_), .Y(_02457_));
NAND_g _22937_ (.A(_02456_), .B(_02457_), .Y(_00727_));
NAND_g _22938_ (.A(_09274_), .B(_02428_), .Y(_02458_));
NAND_g _22939_ (.A(cpuregs[23][14]), .B(_02429_), .Y(_02459_));
NAND_g _22940_ (.A(_02458_), .B(_02459_), .Y(_00728_));
NAND_g _22941_ (.A(_09287_), .B(_02428_), .Y(_02460_));
NAND_g _22942_ (.A(cpuregs[23][15]), .B(_02429_), .Y(_02461_));
NAND_g _22943_ (.A(_02460_), .B(_02461_), .Y(_00729_));
NAND_g _22944_ (.A(_09300_), .B(_02428_), .Y(_02462_));
NAND_g _22945_ (.A(cpuregs[23][16]), .B(_02429_), .Y(_02463_));
NAND_g _22946_ (.A(_02462_), .B(_02463_), .Y(_00730_));
NOR_g _22947_ (.A(cpuregs[23][17]), .B(_02428_), .Y(_02464_));
NOR_g _22948_ (.A(_09313_), .B(_02429_), .Y(_02465_));
NOR_g _22949_ (.A(_02464_), .B(_02465_), .Y(_00731_));
NOR_g _22950_ (.A(cpuregs[23][18]), .B(_02428_), .Y(_02466_));
NOR_g _22951_ (.A(_09325_), .B(_02429_), .Y(_02467_));
NOR_g _22952_ (.A(_02466_), .B(_02467_), .Y(_00732_));
NAND_g _22953_ (.A(_09338_), .B(_02428_), .Y(_02468_));
NAND_g _22954_ (.A(cpuregs[23][19]), .B(_02429_), .Y(_02469_));
NAND_g _22955_ (.A(_02468_), .B(_02469_), .Y(_00733_));
NAND_g _22956_ (.A(_09351_), .B(_02428_), .Y(_02470_));
NAND_g _22957_ (.A(cpuregs[23][20]), .B(_02429_), .Y(_02471_));
NAND_g _22958_ (.A(_02470_), .B(_02471_), .Y(_00734_));
NAND_g _22959_ (.A(_09364_), .B(_02428_), .Y(_02472_));
NAND_g _22960_ (.A(cpuregs[23][21]), .B(_02429_), .Y(_02473_));
NAND_g _22961_ (.A(_02472_), .B(_02473_), .Y(_00735_));
NAND_g _22962_ (.A(_09377_), .B(_02428_), .Y(_02474_));
NAND_g _22963_ (.A(cpuregs[23][22]), .B(_02429_), .Y(_02475_));
NAND_g _22964_ (.A(_02474_), .B(_02475_), .Y(_00736_));
NAND_g _22965_ (.A(_09390_), .B(_02428_), .Y(_02476_));
NAND_g _22966_ (.A(cpuregs[23][23]), .B(_02429_), .Y(_02477_));
NAND_g _22967_ (.A(_02476_), .B(_02477_), .Y(_00737_));
NAND_g _22968_ (.A(_09403_), .B(_02428_), .Y(_02478_));
NAND_g _22969_ (.A(cpuregs[23][24]), .B(_02429_), .Y(_02479_));
NAND_g _22970_ (.A(_02478_), .B(_02479_), .Y(_00738_));
NAND_g _22971_ (.A(_09416_), .B(_02428_), .Y(_02480_));
NAND_g _22972_ (.A(cpuregs[23][25]), .B(_02429_), .Y(_02481_));
NAND_g _22973_ (.A(_02480_), .B(_02481_), .Y(_00739_));
NAND_g _22974_ (.A(_09429_), .B(_02428_), .Y(_02482_));
NAND_g _22975_ (.A(cpuregs[23][26]), .B(_02429_), .Y(_02483_));
NAND_g _22976_ (.A(_02482_), .B(_02483_), .Y(_00740_));
NAND_g _22977_ (.A(_09442_), .B(_02428_), .Y(_02484_));
NAND_g _22978_ (.A(cpuregs[23][27]), .B(_02429_), .Y(_02485_));
NAND_g _22979_ (.A(_02484_), .B(_02485_), .Y(_00741_));
NAND_g _22980_ (.A(_09455_), .B(_02428_), .Y(_02486_));
NAND_g _22981_ (.A(cpuregs[23][28]), .B(_02429_), .Y(_02487_));
NAND_g _22982_ (.A(_02486_), .B(_02487_), .Y(_00742_));
NAND_g _22983_ (.A(_09468_), .B(_02428_), .Y(_02488_));
NAND_g _22984_ (.A(cpuregs[23][29]), .B(_02429_), .Y(_02489_));
NAND_g _22985_ (.A(_02488_), .B(_02489_), .Y(_00743_));
NAND_g _22986_ (.A(_09481_), .B(_02428_), .Y(_02490_));
NAND_g _22987_ (.A(cpuregs[23][30]), .B(_02429_), .Y(_02491_));
NAND_g _22988_ (.A(_02490_), .B(_02491_), .Y(_00744_));
NAND_g _22989_ (.A(_09493_), .B(_02428_), .Y(_02492_));
NAND_g _22990_ (.A(cpuregs[23][31]), .B(_02429_), .Y(_02493_));
NAND_g _22991_ (.A(_02492_), .B(_02493_), .Y(_00745_));
AND_g _22992_ (.A(_09100_), .B(_09566_), .Y(_02494_));
AND_g _22993_ (.A(_14286_), .B(_02494_), .Y(_02495_));
NAND_g _22994_ (.A(_14286_), .B(_02494_), .Y(_02496_));
NAND_g _22995_ (.A(_09098_), .B(_02495_), .Y(_02497_));
NAND_g _22996_ (.A(cpuregs[4][0]), .B(_02496_), .Y(_02498_));
NAND_g _22997_ (.A(_02497_), .B(_02498_), .Y(_00746_));
NAND_g _22998_ (.A(_09109_), .B(_02495_), .Y(_02499_));
NAND_g _22999_ (.A(cpuregs[4][1]), .B(_02496_), .Y(_02500_));
NAND_g _23000_ (.A(_02499_), .B(_02500_), .Y(_00747_));
NAND_g _23001_ (.A(_09118_), .B(_02495_), .Y(_02501_));
NAND_g _23002_ (.A(cpuregs[4][2]), .B(_02496_), .Y(_02502_));
NAND_g _23003_ (.A(_02501_), .B(_02502_), .Y(_00748_));
NAND_g _23004_ (.A(_09131_), .B(_02495_), .Y(_02503_));
NAND_g _23005_ (.A(cpuregs[4][3]), .B(_02496_), .Y(_02504_));
NAND_g _23006_ (.A(_02503_), .B(_02504_), .Y(_00749_));
NAND_g _23007_ (.A(_09144_), .B(_02495_), .Y(_02505_));
NAND_g _23008_ (.A(cpuregs[4][4]), .B(_02496_), .Y(_02506_));
NAND_g _23009_ (.A(_02505_), .B(_02506_), .Y(_00750_));
NAND_g _23010_ (.A(_09157_), .B(_02495_), .Y(_02507_));
NAND_g _23011_ (.A(cpuregs[4][5]), .B(_02496_), .Y(_02508_));
NAND_g _23012_ (.A(_02507_), .B(_02508_), .Y(_00751_));
NAND_g _23013_ (.A(_09170_), .B(_02495_), .Y(_02509_));
NAND_g _23014_ (.A(cpuregs[4][6]), .B(_02496_), .Y(_02510_));
NAND_g _23015_ (.A(_02509_), .B(_02510_), .Y(_00752_));
NAND_g _23016_ (.A(_09183_), .B(_02495_), .Y(_02511_));
NAND_g _23017_ (.A(cpuregs[4][7]), .B(_02496_), .Y(_02512_));
NAND_g _23018_ (.A(_02511_), .B(_02512_), .Y(_00753_));
NAND_g _23019_ (.A(_09196_), .B(_02495_), .Y(_02513_));
NAND_g _23020_ (.A(cpuregs[4][8]), .B(_02496_), .Y(_02514_));
NAND_g _23021_ (.A(_02513_), .B(_02514_), .Y(_00754_));
NAND_g _23022_ (.A(_09209_), .B(_02495_), .Y(_02515_));
NAND_g _23023_ (.A(cpuregs[4][9]), .B(_02496_), .Y(_02516_));
NAND_g _23024_ (.A(_02515_), .B(_02516_), .Y(_00755_));
NAND_g _23025_ (.A(_09222_), .B(_02495_), .Y(_02517_));
NAND_g _23026_ (.A(cpuregs[4][10]), .B(_02496_), .Y(_02518_));
NAND_g _23027_ (.A(_02517_), .B(_02518_), .Y(_00756_));
NAND_g _23028_ (.A(_09235_), .B(_02495_), .Y(_02519_));
NAND_g _23029_ (.A(cpuregs[4][11]), .B(_02496_), .Y(_02520_));
NAND_g _23030_ (.A(_02519_), .B(_02520_), .Y(_00757_));
NAND_g _23031_ (.A(_09248_), .B(_02495_), .Y(_02521_));
NAND_g _23032_ (.A(cpuregs[4][12]), .B(_02496_), .Y(_02522_));
NAND_g _23033_ (.A(_02521_), .B(_02522_), .Y(_00758_));
NAND_g _23034_ (.A(_09261_), .B(_02495_), .Y(_02523_));
NAND_g _23035_ (.A(cpuregs[4][13]), .B(_02496_), .Y(_02524_));
NAND_g _23036_ (.A(_02523_), .B(_02524_), .Y(_00759_));
NAND_g _23037_ (.A(_09274_), .B(_02495_), .Y(_02525_));
NAND_g _23038_ (.A(cpuregs[4][14]), .B(_02496_), .Y(_02526_));
NAND_g _23039_ (.A(_02525_), .B(_02526_), .Y(_00760_));
NAND_g _23040_ (.A(_09287_), .B(_02495_), .Y(_02527_));
NAND_g _23041_ (.A(cpuregs[4][15]), .B(_02496_), .Y(_02528_));
NAND_g _23042_ (.A(_02527_), .B(_02528_), .Y(_00761_));
NAND_g _23043_ (.A(_09300_), .B(_02495_), .Y(_02529_));
NAND_g _23044_ (.A(cpuregs[4][16]), .B(_02496_), .Y(_02530_));
NAND_g _23045_ (.A(_02529_), .B(_02530_), .Y(_00762_));
NOR_g _23046_ (.A(cpuregs[4][17]), .B(_02495_), .Y(_02531_));
NOR_g _23047_ (.A(_09313_), .B(_02496_), .Y(_02532_));
NOR_g _23048_ (.A(_02531_), .B(_02532_), .Y(_00763_));
AND_g _23049_ (.A(_08913_), .B(_02496_), .Y(_02533_));
NOR_g _23050_ (.A(_09325_), .B(_02496_), .Y(_02534_));
NOR_g _23051_ (.A(_02533_), .B(_02534_), .Y(_00764_));
NAND_g _23052_ (.A(_09338_), .B(_02495_), .Y(_02535_));
NAND_g _23053_ (.A(cpuregs[4][19]), .B(_02496_), .Y(_02536_));
NAND_g _23054_ (.A(_02535_), .B(_02536_), .Y(_00765_));
NAND_g _23055_ (.A(_09351_), .B(_02495_), .Y(_02537_));
NAND_g _23056_ (.A(cpuregs[4][20]), .B(_02496_), .Y(_02538_));
NAND_g _23057_ (.A(_02537_), .B(_02538_), .Y(_00766_));
NAND_g _23058_ (.A(_09364_), .B(_02495_), .Y(_02539_));
NAND_g _23059_ (.A(cpuregs[4][21]), .B(_02496_), .Y(_02540_));
NAND_g _23060_ (.A(_02539_), .B(_02540_), .Y(_00767_));
NAND_g _23061_ (.A(_09377_), .B(_02495_), .Y(_02541_));
NAND_g _23062_ (.A(cpuregs[4][22]), .B(_02496_), .Y(_02542_));
NAND_g _23063_ (.A(_02541_), .B(_02542_), .Y(_00768_));
NAND_g _23064_ (.A(_09390_), .B(_02495_), .Y(_02543_));
NAND_g _23065_ (.A(cpuregs[4][23]), .B(_02496_), .Y(_02544_));
NAND_g _23066_ (.A(_02543_), .B(_02544_), .Y(_00769_));
NAND_g _23067_ (.A(_09403_), .B(_02495_), .Y(_02545_));
NAND_g _23068_ (.A(cpuregs[4][24]), .B(_02496_), .Y(_02546_));
NAND_g _23069_ (.A(_02545_), .B(_02546_), .Y(_00770_));
NAND_g _23070_ (.A(_09416_), .B(_02495_), .Y(_02547_));
NAND_g _23071_ (.A(cpuregs[4][25]), .B(_02496_), .Y(_02548_));
NAND_g _23072_ (.A(_02547_), .B(_02548_), .Y(_00771_));
NAND_g _23073_ (.A(_09429_), .B(_02495_), .Y(_02549_));
NAND_g _23074_ (.A(cpuregs[4][26]), .B(_02496_), .Y(_02550_));
NAND_g _23075_ (.A(_02549_), .B(_02550_), .Y(_00772_));
NAND_g _23076_ (.A(_09442_), .B(_02495_), .Y(_02551_));
NAND_g _23077_ (.A(cpuregs[4][27]), .B(_02496_), .Y(_02552_));
NAND_g _23078_ (.A(_02551_), .B(_02552_), .Y(_00773_));
NAND_g _23079_ (.A(_09455_), .B(_02495_), .Y(_02553_));
NAND_g _23080_ (.A(cpuregs[4][28]), .B(_02496_), .Y(_02554_));
NAND_g _23081_ (.A(_02553_), .B(_02554_), .Y(_00774_));
NAND_g _23082_ (.A(_09468_), .B(_02495_), .Y(_02555_));
NAND_g _23083_ (.A(cpuregs[4][29]), .B(_02496_), .Y(_02556_));
NAND_g _23084_ (.A(_02555_), .B(_02556_), .Y(_00775_));
NAND_g _23085_ (.A(_09481_), .B(_02495_), .Y(_02557_));
NAND_g _23086_ (.A(cpuregs[4][30]), .B(_02496_), .Y(_02558_));
NAND_g _23087_ (.A(_02557_), .B(_02558_), .Y(_00776_));
NAND_g _23088_ (.A(_09493_), .B(_02495_), .Y(_02559_));
NAND_g _23089_ (.A(cpuregs[4][31]), .B(_02496_), .Y(_02560_));
NAND_g _23090_ (.A(_02559_), .B(_02560_), .Y(_00777_));
AND_g _23091_ (.A(_09496_), .B(_14285_), .Y(_02561_));
NAND_g _23092_ (.A(_09496_), .B(_14285_), .Y(_02562_));
NAND_g _23093_ (.A(_09098_), .B(_02561_), .Y(_02563_));
NAND_g _23094_ (.A(cpuregs[22][0]), .B(_02562_), .Y(_02564_));
NAND_g _23095_ (.A(_02563_), .B(_02564_), .Y(_00778_));
NAND_g _23096_ (.A(_09109_), .B(_02561_), .Y(_02565_));
NAND_g _23097_ (.A(cpuregs[22][1]), .B(_02562_), .Y(_02566_));
NAND_g _23098_ (.A(_02565_), .B(_02566_), .Y(_00779_));
NAND_g _23099_ (.A(_09118_), .B(_02561_), .Y(_02567_));
NAND_g _23100_ (.A(cpuregs[22][2]), .B(_02562_), .Y(_02568_));
NAND_g _23101_ (.A(_02567_), .B(_02568_), .Y(_00780_));
NAND_g _23102_ (.A(_09131_), .B(_02561_), .Y(_02569_));
NAND_g _23103_ (.A(cpuregs[22][3]), .B(_02562_), .Y(_02570_));
NAND_g _23104_ (.A(_02569_), .B(_02570_), .Y(_00781_));
NAND_g _23105_ (.A(_09144_), .B(_02561_), .Y(_02571_));
NAND_g _23106_ (.A(cpuregs[22][4]), .B(_02562_), .Y(_02572_));
NAND_g _23107_ (.A(_02571_), .B(_02572_), .Y(_00782_));
NAND_g _23108_ (.A(_09157_), .B(_02561_), .Y(_02573_));
NAND_g _23109_ (.A(cpuregs[22][5]), .B(_02562_), .Y(_02574_));
NAND_g _23110_ (.A(_02573_), .B(_02574_), .Y(_00783_));
NAND_g _23111_ (.A(_09170_), .B(_02561_), .Y(_02575_));
NAND_g _23112_ (.A(cpuregs[22][6]), .B(_02562_), .Y(_02576_));
NAND_g _23113_ (.A(_02575_), .B(_02576_), .Y(_00784_));
NAND_g _23114_ (.A(_09183_), .B(_02561_), .Y(_02577_));
NAND_g _23115_ (.A(cpuregs[22][7]), .B(_02562_), .Y(_02578_));
NAND_g _23116_ (.A(_02577_), .B(_02578_), .Y(_00785_));
NAND_g _23117_ (.A(_09196_), .B(_02561_), .Y(_02579_));
NAND_g _23118_ (.A(cpuregs[22][8]), .B(_02562_), .Y(_02580_));
NAND_g _23119_ (.A(_02579_), .B(_02580_), .Y(_00786_));
NAND_g _23120_ (.A(_09209_), .B(_02561_), .Y(_02581_));
NAND_g _23121_ (.A(cpuregs[22][9]), .B(_02562_), .Y(_02582_));
NAND_g _23122_ (.A(_02581_), .B(_02582_), .Y(_00787_));
NAND_g _23123_ (.A(_09222_), .B(_02561_), .Y(_02583_));
NAND_g _23124_ (.A(cpuregs[22][10]), .B(_02562_), .Y(_02584_));
NAND_g _23125_ (.A(_02583_), .B(_02584_), .Y(_00788_));
NAND_g _23126_ (.A(_09235_), .B(_02561_), .Y(_02585_));
NAND_g _23127_ (.A(cpuregs[22][11]), .B(_02562_), .Y(_02586_));
NAND_g _23128_ (.A(_02585_), .B(_02586_), .Y(_00789_));
NAND_g _23129_ (.A(_09248_), .B(_02561_), .Y(_02587_));
NAND_g _23130_ (.A(cpuregs[22][12]), .B(_02562_), .Y(_02588_));
NAND_g _23131_ (.A(_02587_), .B(_02588_), .Y(_00790_));
NAND_g _23132_ (.A(_09261_), .B(_02561_), .Y(_02589_));
NAND_g _23133_ (.A(cpuregs[22][13]), .B(_02562_), .Y(_02590_));
NAND_g _23134_ (.A(_02589_), .B(_02590_), .Y(_00791_));
NAND_g _23135_ (.A(_09274_), .B(_02561_), .Y(_02591_));
NAND_g _23136_ (.A(cpuregs[22][14]), .B(_02562_), .Y(_02592_));
NAND_g _23137_ (.A(_02591_), .B(_02592_), .Y(_00792_));
NAND_g _23138_ (.A(_09287_), .B(_02561_), .Y(_02593_));
NAND_g _23139_ (.A(cpuregs[22][15]), .B(_02562_), .Y(_02594_));
NAND_g _23140_ (.A(_02593_), .B(_02594_), .Y(_00793_));
NAND_g _23141_ (.A(_09300_), .B(_02561_), .Y(_02595_));
NAND_g _23142_ (.A(cpuregs[22][16]), .B(_02562_), .Y(_02596_));
NAND_g _23143_ (.A(_02595_), .B(_02596_), .Y(_00794_));
NOR_g _23144_ (.A(cpuregs[22][17]), .B(_02561_), .Y(_02597_));
NOR_g _23145_ (.A(_09313_), .B(_02562_), .Y(_02598_));
NOR_g _23146_ (.A(_02597_), .B(_02598_), .Y(_00795_));
NOR_g _23147_ (.A(cpuregs[22][18]), .B(_02561_), .Y(_02599_));
NOR_g _23148_ (.A(_09325_), .B(_02562_), .Y(_02600_));
NOR_g _23149_ (.A(_02599_), .B(_02600_), .Y(_00796_));
NAND_g _23150_ (.A(_09338_), .B(_02561_), .Y(_02601_));
NAND_g _23151_ (.A(cpuregs[22][19]), .B(_02562_), .Y(_02602_));
NAND_g _23152_ (.A(_02601_), .B(_02602_), .Y(_00797_));
NAND_g _23153_ (.A(_09351_), .B(_02561_), .Y(_02603_));
NAND_g _23154_ (.A(cpuregs[22][20]), .B(_02562_), .Y(_02604_));
NAND_g _23155_ (.A(_02603_), .B(_02604_), .Y(_00798_));
NAND_g _23156_ (.A(_09364_), .B(_02561_), .Y(_02605_));
NAND_g _23157_ (.A(cpuregs[22][21]), .B(_02562_), .Y(_02606_));
NAND_g _23158_ (.A(_02605_), .B(_02606_), .Y(_00799_));
NAND_g _23159_ (.A(_09377_), .B(_02561_), .Y(_02607_));
NAND_g _23160_ (.A(cpuregs[22][22]), .B(_02562_), .Y(_02608_));
NAND_g _23161_ (.A(_02607_), .B(_02608_), .Y(_00800_));
NAND_g _23162_ (.A(_09390_), .B(_02561_), .Y(_02609_));
NAND_g _23163_ (.A(cpuregs[22][23]), .B(_02562_), .Y(_02610_));
NAND_g _23164_ (.A(_02609_), .B(_02610_), .Y(_00801_));
NAND_g _23165_ (.A(_09403_), .B(_02561_), .Y(_02611_));
NAND_g _23166_ (.A(cpuregs[22][24]), .B(_02562_), .Y(_02612_));
NAND_g _23167_ (.A(_02611_), .B(_02612_), .Y(_00802_));
NAND_g _23168_ (.A(_09416_), .B(_02561_), .Y(_02613_));
NAND_g _23169_ (.A(cpuregs[22][25]), .B(_02562_), .Y(_02614_));
NAND_g _23170_ (.A(_02613_), .B(_02614_), .Y(_00803_));
NAND_g _23171_ (.A(_09429_), .B(_02561_), .Y(_02615_));
NAND_g _23172_ (.A(cpuregs[22][26]), .B(_02562_), .Y(_02616_));
NAND_g _23173_ (.A(_02615_), .B(_02616_), .Y(_00804_));
NAND_g _23174_ (.A(_09442_), .B(_02561_), .Y(_02617_));
NAND_g _23175_ (.A(cpuregs[22][27]), .B(_02562_), .Y(_02618_));
NAND_g _23176_ (.A(_02617_), .B(_02618_), .Y(_00805_));
NAND_g _23177_ (.A(_09455_), .B(_02561_), .Y(_02619_));
NAND_g _23178_ (.A(cpuregs[22][28]), .B(_02562_), .Y(_02620_));
NAND_g _23179_ (.A(_02619_), .B(_02620_), .Y(_00806_));
NAND_g _23180_ (.A(_09468_), .B(_02561_), .Y(_02621_));
NAND_g _23181_ (.A(cpuregs[22][29]), .B(_02562_), .Y(_02622_));
NAND_g _23182_ (.A(_02621_), .B(_02622_), .Y(_00807_));
NAND_g _23183_ (.A(_09481_), .B(_02561_), .Y(_02623_));
NAND_g _23184_ (.A(cpuregs[22][30]), .B(_02562_), .Y(_02624_));
NAND_g _23185_ (.A(_02623_), .B(_02624_), .Y(_00808_));
NAND_g _23186_ (.A(_09493_), .B(_02561_), .Y(_02625_));
NAND_g _23187_ (.A(cpuregs[22][31]), .B(_02562_), .Y(_02626_));
NAND_g _23188_ (.A(_02625_), .B(_02626_), .Y(_00809_));
AND_g _23189_ (.A(_09087_), .B(_09825_), .Y(_02627_));
NAND_g _23190_ (.A(_09087_), .B(_09825_), .Y(_02628_));
NAND_g _23191_ (.A(_09098_), .B(_02627_), .Y(_02629_));
NAND_g _23192_ (.A(cpuregs[13][0]), .B(_02628_), .Y(_02630_));
NAND_g _23193_ (.A(_02629_), .B(_02630_), .Y(_00810_));
NAND_g _23194_ (.A(_09109_), .B(_02627_), .Y(_02631_));
NAND_g _23195_ (.A(cpuregs[13][1]), .B(_02628_), .Y(_02632_));
NAND_g _23196_ (.A(_02631_), .B(_02632_), .Y(_00811_));
NAND_g _23197_ (.A(_09118_), .B(_02627_), .Y(_02633_));
NAND_g _23198_ (.A(cpuregs[13][2]), .B(_02628_), .Y(_02634_));
NAND_g _23199_ (.A(_02633_), .B(_02634_), .Y(_00812_));
NAND_g _23200_ (.A(_09131_), .B(_02627_), .Y(_02635_));
NAND_g _23201_ (.A(cpuregs[13][3]), .B(_02628_), .Y(_02636_));
NAND_g _23202_ (.A(_02635_), .B(_02636_), .Y(_00813_));
NAND_g _23203_ (.A(_09144_), .B(_02627_), .Y(_02637_));
NAND_g _23204_ (.A(cpuregs[13][4]), .B(_02628_), .Y(_02638_));
NAND_g _23205_ (.A(_02637_), .B(_02638_), .Y(_00814_));
NAND_g _23206_ (.A(_09157_), .B(_02627_), .Y(_02639_));
NAND_g _23207_ (.A(cpuregs[13][5]), .B(_02628_), .Y(_02640_));
NAND_g _23208_ (.A(_02639_), .B(_02640_), .Y(_00815_));
NAND_g _23209_ (.A(_09170_), .B(_02627_), .Y(_02641_));
NAND_g _23210_ (.A(cpuregs[13][6]), .B(_02628_), .Y(_02642_));
NAND_g _23211_ (.A(_02641_), .B(_02642_), .Y(_00816_));
NAND_g _23212_ (.A(_09183_), .B(_02627_), .Y(_02643_));
NAND_g _23213_ (.A(cpuregs[13][7]), .B(_02628_), .Y(_02644_));
NAND_g _23214_ (.A(_02643_), .B(_02644_), .Y(_00817_));
NAND_g _23215_ (.A(_09196_), .B(_02627_), .Y(_02645_));
NAND_g _23216_ (.A(cpuregs[13][8]), .B(_02628_), .Y(_02646_));
NAND_g _23217_ (.A(_02645_), .B(_02646_), .Y(_00818_));
NAND_g _23218_ (.A(_09209_), .B(_02627_), .Y(_02647_));
NAND_g _23219_ (.A(cpuregs[13][9]), .B(_02628_), .Y(_02648_));
NAND_g _23220_ (.A(_02647_), .B(_02648_), .Y(_00819_));
NAND_g _23221_ (.A(_09222_), .B(_02627_), .Y(_02649_));
NAND_g _23222_ (.A(cpuregs[13][10]), .B(_02628_), .Y(_02650_));
NAND_g _23223_ (.A(_02649_), .B(_02650_), .Y(_00820_));
NAND_g _23224_ (.A(_09235_), .B(_02627_), .Y(_02651_));
NAND_g _23225_ (.A(cpuregs[13][11]), .B(_02628_), .Y(_02652_));
NAND_g _23226_ (.A(_02651_), .B(_02652_), .Y(_00821_));
NAND_g _23227_ (.A(_09248_), .B(_02627_), .Y(_02653_));
NAND_g _23228_ (.A(cpuregs[13][12]), .B(_02628_), .Y(_02654_));
NAND_g _23229_ (.A(_02653_), .B(_02654_), .Y(_00822_));
NAND_g _23230_ (.A(_09261_), .B(_02627_), .Y(_02655_));
NAND_g _23231_ (.A(cpuregs[13][13]), .B(_02628_), .Y(_02656_));
NAND_g _23232_ (.A(_02655_), .B(_02656_), .Y(_00823_));
NAND_g _23233_ (.A(_09274_), .B(_02627_), .Y(_02657_));
NAND_g _23234_ (.A(cpuregs[13][14]), .B(_02628_), .Y(_02658_));
NAND_g _23235_ (.A(_02657_), .B(_02658_), .Y(_00824_));
NAND_g _23236_ (.A(_09287_), .B(_02627_), .Y(_02659_));
NAND_g _23237_ (.A(cpuregs[13][15]), .B(_02628_), .Y(_02660_));
NAND_g _23238_ (.A(_02659_), .B(_02660_), .Y(_00825_));
NOR_g _23239_ (.A(cpuregs[13][16]), .B(_02627_), .Y(_02661_));
NOR_g _23240_ (.A(_09300_), .B(_02628_), .Y(_02662_));
NOR_g _23241_ (.A(_02661_), .B(_02662_), .Y(_00826_));
NOR_g _23242_ (.A(cpuregs[13][17]), .B(_02627_), .Y(_02663_));
NOR_g _23243_ (.A(_09313_), .B(_02628_), .Y(_02664_));
NOR_g _23244_ (.A(_02663_), .B(_02664_), .Y(_00827_));
NAND_g _23245_ (.A(_09325_), .B(_02627_), .Y(_02665_));
NAND_g _23246_ (.A(cpuregs[13][18]), .B(_02628_), .Y(_02666_));
NAND_g _23247_ (.A(_02665_), .B(_02666_), .Y(_00828_));
NAND_g _23248_ (.A(_09338_), .B(_02627_), .Y(_02667_));
NAND_g _23249_ (.A(cpuregs[13][19]), .B(_02628_), .Y(_02668_));
NAND_g _23250_ (.A(_02667_), .B(_02668_), .Y(_00829_));
NAND_g _23251_ (.A(_09351_), .B(_02627_), .Y(_02669_));
NAND_g _23252_ (.A(cpuregs[13][20]), .B(_02628_), .Y(_02670_));
NAND_g _23253_ (.A(_02669_), .B(_02670_), .Y(_00830_));
NAND_g _23254_ (.A(_09364_), .B(_02627_), .Y(_02671_));
NAND_g _23255_ (.A(cpuregs[13][21]), .B(_02628_), .Y(_02672_));
NAND_g _23256_ (.A(_02671_), .B(_02672_), .Y(_00831_));
NAND_g _23257_ (.A(_09377_), .B(_02627_), .Y(_02673_));
NAND_g _23258_ (.A(cpuregs[13][22]), .B(_02628_), .Y(_02674_));
NAND_g _23259_ (.A(_02673_), .B(_02674_), .Y(_00832_));
NAND_g _23260_ (.A(_09390_), .B(_02627_), .Y(_02675_));
NAND_g _23261_ (.A(cpuregs[13][23]), .B(_02628_), .Y(_02676_));
NAND_g _23262_ (.A(_02675_), .B(_02676_), .Y(_00833_));
NAND_g _23263_ (.A(_09403_), .B(_02627_), .Y(_02677_));
NAND_g _23264_ (.A(cpuregs[13][24]), .B(_02628_), .Y(_02678_));
NAND_g _23265_ (.A(_02677_), .B(_02678_), .Y(_00834_));
NAND_g _23266_ (.A(_09416_), .B(_02627_), .Y(_02679_));
NAND_g _23267_ (.A(cpuregs[13][25]), .B(_02628_), .Y(_02680_));
NAND_g _23268_ (.A(_02679_), .B(_02680_), .Y(_00835_));
NAND_g _23269_ (.A(_09429_), .B(_02627_), .Y(_02681_));
NAND_g _23270_ (.A(cpuregs[13][26]), .B(_02628_), .Y(_02682_));
NAND_g _23271_ (.A(_02681_), .B(_02682_), .Y(_00836_));
NAND_g _23272_ (.A(_09442_), .B(_02627_), .Y(_02683_));
NAND_g _23273_ (.A(cpuregs[13][27]), .B(_02628_), .Y(_02684_));
NAND_g _23274_ (.A(_02683_), .B(_02684_), .Y(_00837_));
NAND_g _23275_ (.A(_09455_), .B(_02627_), .Y(_02685_));
NAND_g _23276_ (.A(cpuregs[13][28]), .B(_02628_), .Y(_02686_));
NAND_g _23277_ (.A(_02685_), .B(_02686_), .Y(_00838_));
NAND_g _23278_ (.A(_09468_), .B(_02627_), .Y(_02687_));
NAND_g _23279_ (.A(cpuregs[13][29]), .B(_02628_), .Y(_02688_));
NAND_g _23280_ (.A(_02687_), .B(_02688_), .Y(_00839_));
NAND_g _23281_ (.A(_09481_), .B(_02627_), .Y(_02689_));
NAND_g _23282_ (.A(cpuregs[13][30]), .B(_02628_), .Y(_02690_));
NAND_g _23283_ (.A(_02689_), .B(_02690_), .Y(_00840_));
NAND_g _23284_ (.A(_09493_), .B(_02627_), .Y(_02691_));
NAND_g _23285_ (.A(cpuregs[13][31]), .B(_02628_), .Y(_02692_));
NAND_g _23286_ (.A(_02691_), .B(_02692_), .Y(_00841_));
AND_g _23287_ (.A(_09077_), .B(_09078_), .Y(_02693_));
AND_g _23288_ (.A(_09085_), .B(_02693_), .Y(_02694_));
NAND_g _23289_ (.A(_09085_), .B(_02693_), .Y(_02695_));
NAND_g _23290_ (.A(_09098_), .B(_02694_), .Y(_02696_));
NAND_g _23291_ (.A(cpuregs[11][0]), .B(_02695_), .Y(_02697_));
NAND_g _23292_ (.A(_02696_), .B(_02697_), .Y(_00842_));
NAND_g _23293_ (.A(_09109_), .B(_02694_), .Y(_02698_));
NAND_g _23294_ (.A(cpuregs[11][1]), .B(_02695_), .Y(_02699_));
NAND_g _23295_ (.A(_02698_), .B(_02699_), .Y(_00843_));
NAND_g _23296_ (.A(_09118_), .B(_02694_), .Y(_02700_));
NAND_g _23297_ (.A(cpuregs[11][2]), .B(_02695_), .Y(_02701_));
NAND_g _23298_ (.A(_02700_), .B(_02701_), .Y(_00844_));
NAND_g _23299_ (.A(_09131_), .B(_02694_), .Y(_02702_));
NAND_g _23300_ (.A(cpuregs[11][3]), .B(_02695_), .Y(_02703_));
NAND_g _23301_ (.A(_02702_), .B(_02703_), .Y(_00845_));
NAND_g _23302_ (.A(_09144_), .B(_02694_), .Y(_02704_));
NAND_g _23303_ (.A(cpuregs[11][4]), .B(_02695_), .Y(_02705_));
NAND_g _23304_ (.A(_02704_), .B(_02705_), .Y(_00846_));
NAND_g _23305_ (.A(_09157_), .B(_02694_), .Y(_02706_));
NAND_g _23306_ (.A(cpuregs[11][5]), .B(_02695_), .Y(_02707_));
NAND_g _23307_ (.A(_02706_), .B(_02707_), .Y(_00847_));
NAND_g _23308_ (.A(_09170_), .B(_02694_), .Y(_02708_));
NAND_g _23309_ (.A(cpuregs[11][6]), .B(_02695_), .Y(_02709_));
NAND_g _23310_ (.A(_02708_), .B(_02709_), .Y(_00848_));
NAND_g _23311_ (.A(_09183_), .B(_02694_), .Y(_02710_));
NAND_g _23312_ (.A(cpuregs[11][7]), .B(_02695_), .Y(_02711_));
NAND_g _23313_ (.A(_02710_), .B(_02711_), .Y(_00849_));
NAND_g _23314_ (.A(_09196_), .B(_02694_), .Y(_02712_));
NAND_g _23315_ (.A(cpuregs[11][8]), .B(_02695_), .Y(_02713_));
NAND_g _23316_ (.A(_02712_), .B(_02713_), .Y(_00850_));
NAND_g _23317_ (.A(_09209_), .B(_02694_), .Y(_02714_));
NAND_g _23318_ (.A(cpuregs[11][9]), .B(_02695_), .Y(_02715_));
NAND_g _23319_ (.A(_02714_), .B(_02715_), .Y(_00851_));
NAND_g _23320_ (.A(_09222_), .B(_02694_), .Y(_02716_));
NAND_g _23321_ (.A(cpuregs[11][10]), .B(_02695_), .Y(_02717_));
NAND_g _23322_ (.A(_02716_), .B(_02717_), .Y(_00852_));
NAND_g _23323_ (.A(_09235_), .B(_02694_), .Y(_02718_));
NAND_g _23324_ (.A(cpuregs[11][11]), .B(_02695_), .Y(_02719_));
NAND_g _23325_ (.A(_02718_), .B(_02719_), .Y(_00853_));
NAND_g _23326_ (.A(_09248_), .B(_02694_), .Y(_02720_));
NAND_g _23327_ (.A(cpuregs[11][12]), .B(_02695_), .Y(_02721_));
NAND_g _23328_ (.A(_02720_), .B(_02721_), .Y(_00854_));
NAND_g _23329_ (.A(_09261_), .B(_02694_), .Y(_02722_));
NAND_g _23330_ (.A(cpuregs[11][13]), .B(_02695_), .Y(_02723_));
NAND_g _23331_ (.A(_02722_), .B(_02723_), .Y(_00855_));
NAND_g _23332_ (.A(_09274_), .B(_02694_), .Y(_02724_));
NAND_g _23333_ (.A(cpuregs[11][14]), .B(_02695_), .Y(_02725_));
NAND_g _23334_ (.A(_02724_), .B(_02725_), .Y(_00856_));
NAND_g _23335_ (.A(_09287_), .B(_02694_), .Y(_02726_));
NAND_g _23336_ (.A(cpuregs[11][15]), .B(_02695_), .Y(_02727_));
NAND_g _23337_ (.A(_02726_), .B(_02727_), .Y(_00857_));
NOR_g _23338_ (.A(cpuregs[11][16]), .B(_02694_), .Y(_02728_));
NOR_g _23339_ (.A(_09300_), .B(_02695_), .Y(_02729_));
NOR_g _23340_ (.A(_02728_), .B(_02729_), .Y(_00858_));
NOR_g _23341_ (.A(cpuregs[11][17]), .B(_02694_), .Y(_02730_));
NOR_g _23342_ (.A(_09313_), .B(_02695_), .Y(_02731_));
NOR_g _23343_ (.A(_02730_), .B(_02731_), .Y(_00859_));
NAND_g _23344_ (.A(_09325_), .B(_02694_), .Y(_02732_));
NAND_g _23345_ (.A(cpuregs[11][18]), .B(_02695_), .Y(_02733_));
NAND_g _23346_ (.A(_02732_), .B(_02733_), .Y(_00860_));
NAND_g _23347_ (.A(_09338_), .B(_02694_), .Y(_02734_));
NAND_g _23348_ (.A(cpuregs[11][19]), .B(_02695_), .Y(_02735_));
NAND_g _23349_ (.A(_02734_), .B(_02735_), .Y(_00861_));
NAND_g _23350_ (.A(_09351_), .B(_02694_), .Y(_02736_));
NAND_g _23351_ (.A(cpuregs[11][20]), .B(_02695_), .Y(_02737_));
NAND_g _23352_ (.A(_02736_), .B(_02737_), .Y(_00862_));
NAND_g _23353_ (.A(_09364_), .B(_02694_), .Y(_02738_));
NAND_g _23354_ (.A(cpuregs[11][21]), .B(_02695_), .Y(_02739_));
NAND_g _23355_ (.A(_02738_), .B(_02739_), .Y(_00863_));
NAND_g _23356_ (.A(_09377_), .B(_02694_), .Y(_02740_));
NAND_g _23357_ (.A(cpuregs[11][22]), .B(_02695_), .Y(_02741_));
NAND_g _23358_ (.A(_02740_), .B(_02741_), .Y(_00864_));
NAND_g _23359_ (.A(_09390_), .B(_02694_), .Y(_02742_));
NAND_g _23360_ (.A(cpuregs[11][23]), .B(_02695_), .Y(_02743_));
NAND_g _23361_ (.A(_02742_), .B(_02743_), .Y(_00865_));
NAND_g _23362_ (.A(_09403_), .B(_02694_), .Y(_02744_));
NAND_g _23363_ (.A(cpuregs[11][24]), .B(_02695_), .Y(_02745_));
NAND_g _23364_ (.A(_02744_), .B(_02745_), .Y(_00866_));
NAND_g _23365_ (.A(_09416_), .B(_02694_), .Y(_02746_));
NAND_g _23366_ (.A(cpuregs[11][25]), .B(_02695_), .Y(_02747_));
NAND_g _23367_ (.A(_02746_), .B(_02747_), .Y(_00867_));
NAND_g _23368_ (.A(_09429_), .B(_02694_), .Y(_02748_));
NAND_g _23369_ (.A(cpuregs[11][26]), .B(_02695_), .Y(_02749_));
NAND_g _23370_ (.A(_02748_), .B(_02749_), .Y(_00868_));
NAND_g _23371_ (.A(_09442_), .B(_02694_), .Y(_02750_));
NAND_g _23372_ (.A(cpuregs[11][27]), .B(_02695_), .Y(_02751_));
NAND_g _23373_ (.A(_02750_), .B(_02751_), .Y(_00869_));
NAND_g _23374_ (.A(_09455_), .B(_02694_), .Y(_02752_));
NAND_g _23375_ (.A(cpuregs[11][28]), .B(_02695_), .Y(_02753_));
NAND_g _23376_ (.A(_02752_), .B(_02753_), .Y(_00870_));
NAND_g _23377_ (.A(_09468_), .B(_02694_), .Y(_02754_));
NAND_g _23378_ (.A(cpuregs[11][29]), .B(_02695_), .Y(_02755_));
NAND_g _23379_ (.A(_02754_), .B(_02755_), .Y(_00871_));
NAND_g _23380_ (.A(_09481_), .B(_02694_), .Y(_02756_));
NAND_g _23381_ (.A(cpuregs[11][30]), .B(_02695_), .Y(_02757_));
NAND_g _23382_ (.A(_02756_), .B(_02757_), .Y(_00872_));
NAND_g _23383_ (.A(_09493_), .B(_02694_), .Y(_02758_));
NAND_g _23384_ (.A(cpuregs[11][31]), .B(_02695_), .Y(_02759_));
NAND_g _23385_ (.A(_02758_), .B(_02759_), .Y(_00873_));
AND_g _23386_ (.A(_08853_), .B(_14284_), .Y(_02760_));
AND_g _23387_ (.A(_09496_), .B(_02760_), .Y(_02761_));
NAND_g _23388_ (.A(_09496_), .B(_02760_), .Y(_02762_));
NAND_g _23389_ (.A(_09098_), .B(_02761_), .Y(_02763_));
NAND_g _23390_ (.A(cpuregs[18][0]), .B(_02762_), .Y(_02764_));
NAND_g _23391_ (.A(_02763_), .B(_02764_), .Y(_00874_));
NAND_g _23392_ (.A(_09109_), .B(_02761_), .Y(_02765_));
NAND_g _23393_ (.A(cpuregs[18][1]), .B(_02762_), .Y(_02766_));
NAND_g _23394_ (.A(_02765_), .B(_02766_), .Y(_00875_));
NAND_g _23395_ (.A(_09118_), .B(_02761_), .Y(_02767_));
NAND_g _23396_ (.A(cpuregs[18][2]), .B(_02762_), .Y(_02768_));
NAND_g _23397_ (.A(_02767_), .B(_02768_), .Y(_00876_));
NAND_g _23398_ (.A(_09131_), .B(_02761_), .Y(_02769_));
NAND_g _23399_ (.A(cpuregs[18][3]), .B(_02762_), .Y(_02770_));
NAND_g _23400_ (.A(_02769_), .B(_02770_), .Y(_00877_));
NAND_g _23401_ (.A(_09144_), .B(_02761_), .Y(_02771_));
NAND_g _23402_ (.A(cpuregs[18][4]), .B(_02762_), .Y(_02772_));
NAND_g _23403_ (.A(_02771_), .B(_02772_), .Y(_00878_));
NAND_g _23404_ (.A(_09157_), .B(_02761_), .Y(_02773_));
NAND_g _23405_ (.A(cpuregs[18][5]), .B(_02762_), .Y(_02774_));
NAND_g _23406_ (.A(_02773_), .B(_02774_), .Y(_00879_));
NAND_g _23407_ (.A(_09170_), .B(_02761_), .Y(_02775_));
NAND_g _23408_ (.A(cpuregs[18][6]), .B(_02762_), .Y(_02776_));
NAND_g _23409_ (.A(_02775_), .B(_02776_), .Y(_00880_));
NAND_g _23410_ (.A(_09183_), .B(_02761_), .Y(_02777_));
NAND_g _23411_ (.A(cpuregs[18][7]), .B(_02762_), .Y(_02778_));
NAND_g _23412_ (.A(_02777_), .B(_02778_), .Y(_00881_));
NAND_g _23413_ (.A(_09196_), .B(_02761_), .Y(_02779_));
NAND_g _23414_ (.A(cpuregs[18][8]), .B(_02762_), .Y(_02780_));
NAND_g _23415_ (.A(_02779_), .B(_02780_), .Y(_00882_));
NAND_g _23416_ (.A(_09209_), .B(_02761_), .Y(_02781_));
NAND_g _23417_ (.A(cpuregs[18][9]), .B(_02762_), .Y(_02782_));
NAND_g _23418_ (.A(_02781_), .B(_02782_), .Y(_00883_));
NAND_g _23419_ (.A(_09222_), .B(_02761_), .Y(_02783_));
NAND_g _23420_ (.A(cpuregs[18][10]), .B(_02762_), .Y(_02784_));
NAND_g _23421_ (.A(_02783_), .B(_02784_), .Y(_00884_));
NAND_g _23422_ (.A(_09235_), .B(_02761_), .Y(_02785_));
NAND_g _23423_ (.A(cpuregs[18][11]), .B(_02762_), .Y(_02786_));
NAND_g _23424_ (.A(_02785_), .B(_02786_), .Y(_00885_));
NAND_g _23425_ (.A(_09248_), .B(_02761_), .Y(_02787_));
NAND_g _23426_ (.A(cpuregs[18][12]), .B(_02762_), .Y(_02788_));
NAND_g _23427_ (.A(_02787_), .B(_02788_), .Y(_00886_));
NAND_g _23428_ (.A(_09261_), .B(_02761_), .Y(_02789_));
NAND_g _23429_ (.A(cpuregs[18][13]), .B(_02762_), .Y(_02790_));
NAND_g _23430_ (.A(_02789_), .B(_02790_), .Y(_00887_));
NAND_g _23431_ (.A(_09274_), .B(_02761_), .Y(_02791_));
NAND_g _23432_ (.A(cpuregs[18][14]), .B(_02762_), .Y(_02792_));
NAND_g _23433_ (.A(_02791_), .B(_02792_), .Y(_00888_));
NAND_g _23434_ (.A(_09287_), .B(_02761_), .Y(_02793_));
NAND_g _23435_ (.A(cpuregs[18][15]), .B(_02762_), .Y(_02794_));
NAND_g _23436_ (.A(_02793_), .B(_02794_), .Y(_00889_));
NAND_g _23437_ (.A(_09300_), .B(_02761_), .Y(_02795_));
NAND_g _23438_ (.A(cpuregs[18][16]), .B(_02762_), .Y(_02796_));
NAND_g _23439_ (.A(_02795_), .B(_02796_), .Y(_00890_));
NOR_g _23440_ (.A(cpuregs[18][17]), .B(_02761_), .Y(_02797_));
NOR_g _23441_ (.A(_09313_), .B(_02762_), .Y(_02798_));
NOR_g _23442_ (.A(_02797_), .B(_02798_), .Y(_00891_));
NOR_g _23443_ (.A(cpuregs[18][18]), .B(_02761_), .Y(_02799_));
NOR_g _23444_ (.A(_09325_), .B(_02762_), .Y(_02800_));
NOR_g _23445_ (.A(_02799_), .B(_02800_), .Y(_00892_));
NAND_g _23446_ (.A(_09338_), .B(_02761_), .Y(_02801_));
NAND_g _23447_ (.A(cpuregs[18][19]), .B(_02762_), .Y(_02802_));
NAND_g _23448_ (.A(_02801_), .B(_02802_), .Y(_00893_));
NAND_g _23449_ (.A(_09351_), .B(_02761_), .Y(_02803_));
NAND_g _23450_ (.A(cpuregs[18][20]), .B(_02762_), .Y(_02804_));
NAND_g _23451_ (.A(_02803_), .B(_02804_), .Y(_00894_));
NAND_g _23452_ (.A(_09364_), .B(_02761_), .Y(_02805_));
NAND_g _23453_ (.A(cpuregs[18][21]), .B(_02762_), .Y(_02806_));
NAND_g _23454_ (.A(_02805_), .B(_02806_), .Y(_00895_));
NAND_g _23455_ (.A(_09377_), .B(_02761_), .Y(_02807_));
NAND_g _23456_ (.A(cpuregs[18][22]), .B(_02762_), .Y(_02808_));
NAND_g _23457_ (.A(_02807_), .B(_02808_), .Y(_00896_));
NAND_g _23458_ (.A(_09390_), .B(_02761_), .Y(_02809_));
NAND_g _23459_ (.A(cpuregs[18][23]), .B(_02762_), .Y(_02810_));
NAND_g _23460_ (.A(_02809_), .B(_02810_), .Y(_00897_));
NAND_g _23461_ (.A(_09403_), .B(_02761_), .Y(_02811_));
NAND_g _23462_ (.A(cpuregs[18][24]), .B(_02762_), .Y(_02812_));
NAND_g _23463_ (.A(_02811_), .B(_02812_), .Y(_00898_));
NAND_g _23464_ (.A(_09416_), .B(_02761_), .Y(_02813_));
NAND_g _23465_ (.A(cpuregs[18][25]), .B(_02762_), .Y(_02814_));
NAND_g _23466_ (.A(_02813_), .B(_02814_), .Y(_00899_));
NAND_g _23467_ (.A(_09429_), .B(_02761_), .Y(_02815_));
NAND_g _23468_ (.A(cpuregs[18][26]), .B(_02762_), .Y(_02816_));
NAND_g _23469_ (.A(_02815_), .B(_02816_), .Y(_00900_));
NAND_g _23470_ (.A(_09442_), .B(_02761_), .Y(_02817_));
NAND_g _23471_ (.A(cpuregs[18][27]), .B(_02762_), .Y(_02818_));
NAND_g _23472_ (.A(_02817_), .B(_02818_), .Y(_00901_));
NAND_g _23473_ (.A(_09455_), .B(_02761_), .Y(_02819_));
NAND_g _23474_ (.A(cpuregs[18][28]), .B(_02762_), .Y(_02820_));
NAND_g _23475_ (.A(_02819_), .B(_02820_), .Y(_00902_));
NAND_g _23476_ (.A(_09468_), .B(_02761_), .Y(_02821_));
NAND_g _23477_ (.A(cpuregs[18][29]), .B(_02762_), .Y(_02822_));
NAND_g _23478_ (.A(_02821_), .B(_02822_), .Y(_00903_));
NAND_g _23479_ (.A(_09481_), .B(_02761_), .Y(_02823_));
NAND_g _23480_ (.A(cpuregs[18][30]), .B(_02762_), .Y(_02824_));
NAND_g _23481_ (.A(_02823_), .B(_02824_), .Y(_00904_));
NAND_g _23482_ (.A(_09493_), .B(_02761_), .Y(_02825_));
NAND_g _23483_ (.A(cpuregs[18][31]), .B(_02762_), .Y(_02826_));
NAND_g _23484_ (.A(_02825_), .B(_02826_), .Y(_00905_));
AND_g _23485_ (.A(_09087_), .B(_09496_), .Y(_02827_));
NAND_g _23486_ (.A(_09087_), .B(_09496_), .Y(_02828_));
NAND_g _23487_ (.A(cpuregs[14][0]), .B(_02828_), .Y(_02829_));
NAND_g _23488_ (.A(_09098_), .B(_02827_), .Y(_02830_));
NAND_g _23489_ (.A(_02829_), .B(_02830_), .Y(_00906_));
NAND_g _23490_ (.A(cpuregs[14][1]), .B(_02828_), .Y(_02831_));
NAND_g _23491_ (.A(_09109_), .B(_02827_), .Y(_02832_));
NAND_g _23492_ (.A(_02831_), .B(_02832_), .Y(_00907_));
NAND_g _23493_ (.A(cpuregs[14][2]), .B(_02828_), .Y(_02833_));
NAND_g _23494_ (.A(_09118_), .B(_02827_), .Y(_02834_));
NAND_g _23495_ (.A(_02833_), .B(_02834_), .Y(_00908_));
NAND_g _23496_ (.A(cpuregs[14][3]), .B(_02828_), .Y(_02835_));
NAND_g _23497_ (.A(_09131_), .B(_02827_), .Y(_02836_));
NAND_g _23498_ (.A(_02835_), .B(_02836_), .Y(_00909_));
NAND_g _23499_ (.A(cpuregs[14][4]), .B(_02828_), .Y(_02837_));
NAND_g _23500_ (.A(_09144_), .B(_02827_), .Y(_02838_));
NAND_g _23501_ (.A(_02837_), .B(_02838_), .Y(_00910_));
NAND_g _23502_ (.A(cpuregs[14][5]), .B(_02828_), .Y(_02839_));
NAND_g _23503_ (.A(_09157_), .B(_02827_), .Y(_02840_));
NAND_g _23504_ (.A(_02839_), .B(_02840_), .Y(_00911_));
NAND_g _23505_ (.A(cpuregs[14][6]), .B(_02828_), .Y(_02841_));
NAND_g _23506_ (.A(_09170_), .B(_02827_), .Y(_02842_));
NAND_g _23507_ (.A(_02841_), .B(_02842_), .Y(_00912_));
NAND_g _23508_ (.A(cpuregs[14][7]), .B(_02828_), .Y(_02843_));
NAND_g _23509_ (.A(_09183_), .B(_02827_), .Y(_02844_));
NAND_g _23510_ (.A(_02843_), .B(_02844_), .Y(_00913_));
NAND_g _23511_ (.A(cpuregs[14][8]), .B(_02828_), .Y(_02845_));
NAND_g _23512_ (.A(_09196_), .B(_02827_), .Y(_02846_));
NAND_g _23513_ (.A(_02845_), .B(_02846_), .Y(_00914_));
NAND_g _23514_ (.A(cpuregs[14][9]), .B(_02828_), .Y(_02847_));
NAND_g _23515_ (.A(_09209_), .B(_02827_), .Y(_02848_));
NAND_g _23516_ (.A(_02847_), .B(_02848_), .Y(_00915_));
NAND_g _23517_ (.A(cpuregs[14][10]), .B(_02828_), .Y(_02849_));
NAND_g _23518_ (.A(_09222_), .B(_02827_), .Y(_02850_));
NAND_g _23519_ (.A(_02849_), .B(_02850_), .Y(_00916_));
NAND_g _23520_ (.A(cpuregs[14][11]), .B(_02828_), .Y(_02851_));
NAND_g _23521_ (.A(_09235_), .B(_02827_), .Y(_02852_));
NAND_g _23522_ (.A(_02851_), .B(_02852_), .Y(_00917_));
NAND_g _23523_ (.A(cpuregs[14][12]), .B(_02828_), .Y(_02853_));
NAND_g _23524_ (.A(_09248_), .B(_02827_), .Y(_02854_));
NAND_g _23525_ (.A(_02853_), .B(_02854_), .Y(_00918_));
NAND_g _23526_ (.A(cpuregs[14][13]), .B(_02828_), .Y(_02855_));
NAND_g _23527_ (.A(_09261_), .B(_02827_), .Y(_02856_));
NAND_g _23528_ (.A(_02855_), .B(_02856_), .Y(_00919_));
NAND_g _23529_ (.A(cpuregs[14][14]), .B(_02828_), .Y(_02857_));
NAND_g _23530_ (.A(_09274_), .B(_02827_), .Y(_02858_));
NAND_g _23531_ (.A(_02857_), .B(_02858_), .Y(_00920_));
NAND_g _23532_ (.A(cpuregs[14][15]), .B(_02828_), .Y(_02859_));
NAND_g _23533_ (.A(_09287_), .B(_02827_), .Y(_02860_));
NAND_g _23534_ (.A(_02859_), .B(_02860_), .Y(_00921_));
NOR_g _23535_ (.A(cpuregs[14][16]), .B(_02827_), .Y(_02861_));
NOR_g _23536_ (.A(_09300_), .B(_02828_), .Y(_02862_));
NOR_g _23537_ (.A(_02861_), .B(_02862_), .Y(_00922_));
NOR_g _23538_ (.A(cpuregs[14][17]), .B(_02827_), .Y(_02863_));
NOR_g _23539_ (.A(_09313_), .B(_02828_), .Y(_02864_));
NOR_g _23540_ (.A(_02863_), .B(_02864_), .Y(_00923_));
NOR_g _23541_ (.A(cpuregs[14][18]), .B(_02827_), .Y(_02865_));
NOR_g _23542_ (.A(_09325_), .B(_02828_), .Y(_02866_));
NOR_g _23543_ (.A(_02865_), .B(_02866_), .Y(_00924_));
AND_g _23544_ (.A(_08939_), .B(_02828_), .Y(_02867_));
NOR_g _23545_ (.A(_09338_), .B(_02828_), .Y(_02868_));
NOR_g _23546_ (.A(_02867_), .B(_02868_), .Y(_00925_));
AND_g _23547_ (.A(_08940_), .B(_02828_), .Y(_02869_));
NOR_g _23548_ (.A(_09351_), .B(_02828_), .Y(_02870_));
NOR_g _23549_ (.A(_02869_), .B(_02870_), .Y(_00926_));
NOR_g _23550_ (.A(cpuregs[14][21]), .B(_02827_), .Y(_02871_));
NOR_g _23551_ (.A(_09364_), .B(_02828_), .Y(_02872_));
NOR_g _23552_ (.A(_02871_), .B(_02872_), .Y(_00927_));
NOR_g _23553_ (.A(cpuregs[14][22]), .B(_02827_), .Y(_02873_));
NOR_g _23554_ (.A(_09377_), .B(_02828_), .Y(_02874_));
NOR_g _23555_ (.A(_02873_), .B(_02874_), .Y(_00928_));
NOR_g _23556_ (.A(cpuregs[14][23]), .B(_02827_), .Y(_02875_));
NOR_g _23557_ (.A(_09390_), .B(_02828_), .Y(_02876_));
NOR_g _23558_ (.A(_02875_), .B(_02876_), .Y(_00929_));
NOR_g _23559_ (.A(cpuregs[14][24]), .B(_02827_), .Y(_02877_));
NOR_g _23560_ (.A(_09403_), .B(_02828_), .Y(_02878_));
NOR_g _23561_ (.A(_02877_), .B(_02878_), .Y(_00930_));
NOR_g _23562_ (.A(cpuregs[14][25]), .B(_02827_), .Y(_02879_));
NOR_g _23563_ (.A(_09416_), .B(_02828_), .Y(_02880_));
NOR_g _23564_ (.A(_02879_), .B(_02880_), .Y(_00931_));
NOR_g _23565_ (.A(cpuregs[14][26]), .B(_02827_), .Y(_02881_));
NOR_g _23566_ (.A(_09429_), .B(_02828_), .Y(_02882_));
NOR_g _23567_ (.A(_02881_), .B(_02882_), .Y(_00932_));
NOR_g _23568_ (.A(cpuregs[14][27]), .B(_02827_), .Y(_02883_));
NOR_g _23569_ (.A(_09442_), .B(_02828_), .Y(_02884_));
NOR_g _23570_ (.A(_02883_), .B(_02884_), .Y(_00933_));
NOR_g _23571_ (.A(cpuregs[14][28]), .B(_02827_), .Y(_02885_));
NOR_g _23572_ (.A(_09455_), .B(_02828_), .Y(_02886_));
NOR_g _23573_ (.A(_02885_), .B(_02886_), .Y(_00934_));
NOR_g _23574_ (.A(cpuregs[14][29]), .B(_02827_), .Y(_02887_));
NOR_g _23575_ (.A(_09468_), .B(_02828_), .Y(_02888_));
NOR_g _23576_ (.A(_02887_), .B(_02888_), .Y(_00935_));
NOR_g _23577_ (.A(cpuregs[14][30]), .B(_02827_), .Y(_02889_));
NOR_g _23578_ (.A(_09481_), .B(_02828_), .Y(_02890_));
NOR_g _23579_ (.A(_02889_), .B(_02890_), .Y(_00936_));
NOR_g _23580_ (.A(cpuregs[14][31]), .B(_02827_), .Y(_02891_));
NOR_g _23581_ (.A(_09493_), .B(_02828_), .Y(_02892_));
NOR_g _23582_ (.A(_02891_), .B(_02892_), .Y(_00937_));
AND_g _23583_ (.A(_09825_), .B(_02760_), .Y(_02893_));
NAND_g _23584_ (.A(_09825_), .B(_02760_), .Y(_02894_));
NAND_g _23585_ (.A(_09098_), .B(_02893_), .Y(_02895_));
NAND_g _23586_ (.A(cpuregs[17][0]), .B(_02894_), .Y(_02896_));
NAND_g _23587_ (.A(_02895_), .B(_02896_), .Y(_00938_));
NAND_g _23588_ (.A(_09109_), .B(_02893_), .Y(_02897_));
NAND_g _23589_ (.A(cpuregs[17][1]), .B(_02894_), .Y(_02898_));
NAND_g _23590_ (.A(_02897_), .B(_02898_), .Y(_00939_));
NAND_g _23591_ (.A(_09118_), .B(_02893_), .Y(_02899_));
NAND_g _23592_ (.A(cpuregs[17][2]), .B(_02894_), .Y(_02900_));
NAND_g _23593_ (.A(_02899_), .B(_02900_), .Y(_00940_));
NAND_g _23594_ (.A(_09131_), .B(_02893_), .Y(_02901_));
NAND_g _23595_ (.A(cpuregs[17][3]), .B(_02894_), .Y(_02902_));
NAND_g _23596_ (.A(_02901_), .B(_02902_), .Y(_00941_));
NAND_g _23597_ (.A(_09144_), .B(_02893_), .Y(_02903_));
NAND_g _23598_ (.A(cpuregs[17][4]), .B(_02894_), .Y(_02904_));
NAND_g _23599_ (.A(_02903_), .B(_02904_), .Y(_00942_));
NAND_g _23600_ (.A(_09157_), .B(_02893_), .Y(_02905_));
NAND_g _23601_ (.A(cpuregs[17][5]), .B(_02894_), .Y(_02906_));
NAND_g _23602_ (.A(_02905_), .B(_02906_), .Y(_00943_));
NAND_g _23603_ (.A(_09170_), .B(_02893_), .Y(_02907_));
NAND_g _23604_ (.A(cpuregs[17][6]), .B(_02894_), .Y(_02908_));
NAND_g _23605_ (.A(_02907_), .B(_02908_), .Y(_00944_));
NAND_g _23606_ (.A(_09183_), .B(_02893_), .Y(_02909_));
NAND_g _23607_ (.A(cpuregs[17][7]), .B(_02894_), .Y(_02910_));
NAND_g _23608_ (.A(_02909_), .B(_02910_), .Y(_00945_));
NAND_g _23609_ (.A(_09196_), .B(_02893_), .Y(_02911_));
NAND_g _23610_ (.A(cpuregs[17][8]), .B(_02894_), .Y(_02912_));
NAND_g _23611_ (.A(_02911_), .B(_02912_), .Y(_00946_));
NAND_g _23612_ (.A(_09209_), .B(_02893_), .Y(_02913_));
NAND_g _23613_ (.A(cpuregs[17][9]), .B(_02894_), .Y(_02914_));
NAND_g _23614_ (.A(_02913_), .B(_02914_), .Y(_00947_));
NAND_g _23615_ (.A(_09222_), .B(_02893_), .Y(_02915_));
NAND_g _23616_ (.A(cpuregs[17][10]), .B(_02894_), .Y(_02916_));
NAND_g _23617_ (.A(_02915_), .B(_02916_), .Y(_00948_));
NAND_g _23618_ (.A(_09235_), .B(_02893_), .Y(_02917_));
NAND_g _23619_ (.A(cpuregs[17][11]), .B(_02894_), .Y(_02918_));
NAND_g _23620_ (.A(_02917_), .B(_02918_), .Y(_00949_));
NAND_g _23621_ (.A(_09248_), .B(_02893_), .Y(_02919_));
NAND_g _23622_ (.A(cpuregs[17][12]), .B(_02894_), .Y(_02920_));
NAND_g _23623_ (.A(_02919_), .B(_02920_), .Y(_00950_));
NAND_g _23624_ (.A(_09261_), .B(_02893_), .Y(_02921_));
NAND_g _23625_ (.A(cpuregs[17][13]), .B(_02894_), .Y(_02922_));
NAND_g _23626_ (.A(_02921_), .B(_02922_), .Y(_00951_));
NAND_g _23627_ (.A(_09274_), .B(_02893_), .Y(_02923_));
NAND_g _23628_ (.A(cpuregs[17][14]), .B(_02894_), .Y(_02924_));
NAND_g _23629_ (.A(_02923_), .B(_02924_), .Y(_00952_));
NAND_g _23630_ (.A(_09287_), .B(_02893_), .Y(_02925_));
NAND_g _23631_ (.A(cpuregs[17][15]), .B(_02894_), .Y(_02926_));
NAND_g _23632_ (.A(_02925_), .B(_02926_), .Y(_00953_));
NAND_g _23633_ (.A(_09300_), .B(_02893_), .Y(_02927_));
NAND_g _23634_ (.A(cpuregs[17][16]), .B(_02894_), .Y(_02928_));
NAND_g _23635_ (.A(_02927_), .B(_02928_), .Y(_00954_));
NOR_g _23636_ (.A(cpuregs[17][17]), .B(_02893_), .Y(_02929_));
NOR_g _23637_ (.A(_09313_), .B(_02894_), .Y(_02930_));
NOR_g _23638_ (.A(_02929_), .B(_02930_), .Y(_00955_));
NOR_g _23639_ (.A(cpuregs[17][18]), .B(_02893_), .Y(_02931_));
NOR_g _23640_ (.A(_09325_), .B(_02894_), .Y(_02932_));
NOR_g _23641_ (.A(_02931_), .B(_02932_), .Y(_00956_));
NAND_g _23642_ (.A(_09338_), .B(_02893_), .Y(_02933_));
NAND_g _23643_ (.A(cpuregs[17][19]), .B(_02894_), .Y(_02934_));
NAND_g _23644_ (.A(_02933_), .B(_02934_), .Y(_00957_));
NAND_g _23645_ (.A(_09351_), .B(_02893_), .Y(_02935_));
NAND_g _23646_ (.A(cpuregs[17][20]), .B(_02894_), .Y(_02936_));
NAND_g _23647_ (.A(_02935_), .B(_02936_), .Y(_00958_));
NAND_g _23648_ (.A(_09364_), .B(_02893_), .Y(_02937_));
NAND_g _23649_ (.A(cpuregs[17][21]), .B(_02894_), .Y(_02938_));
NAND_g _23650_ (.A(_02937_), .B(_02938_), .Y(_00959_));
NAND_g _23651_ (.A(_09377_), .B(_02893_), .Y(_02939_));
NAND_g _23652_ (.A(cpuregs[17][22]), .B(_02894_), .Y(_02940_));
NAND_g _23653_ (.A(_02939_), .B(_02940_), .Y(_00960_));
NAND_g _23654_ (.A(_09390_), .B(_02893_), .Y(_02941_));
NAND_g _23655_ (.A(cpuregs[17][23]), .B(_02894_), .Y(_02942_));
NAND_g _23656_ (.A(_02941_), .B(_02942_), .Y(_00961_));
NAND_g _23657_ (.A(_09403_), .B(_02893_), .Y(_02943_));
NAND_g _23658_ (.A(cpuregs[17][24]), .B(_02894_), .Y(_02944_));
NAND_g _23659_ (.A(_02943_), .B(_02944_), .Y(_00962_));
NAND_g _23660_ (.A(_09416_), .B(_02893_), .Y(_02945_));
NAND_g _23661_ (.A(cpuregs[17][25]), .B(_02894_), .Y(_02946_));
NAND_g _23662_ (.A(_02945_), .B(_02946_), .Y(_00963_));
NAND_g _23663_ (.A(_09429_), .B(_02893_), .Y(_02947_));
NAND_g _23664_ (.A(cpuregs[17][26]), .B(_02894_), .Y(_02948_));
NAND_g _23665_ (.A(_02947_), .B(_02948_), .Y(_00964_));
NAND_g _23666_ (.A(_09442_), .B(_02893_), .Y(_02949_));
NAND_g _23667_ (.A(cpuregs[17][27]), .B(_02894_), .Y(_02950_));
NAND_g _23668_ (.A(_02949_), .B(_02950_), .Y(_00965_));
NAND_g _23669_ (.A(_09455_), .B(_02893_), .Y(_02951_));
NAND_g _23670_ (.A(cpuregs[17][28]), .B(_02894_), .Y(_02952_));
NAND_g _23671_ (.A(_02951_), .B(_02952_), .Y(_00966_));
NAND_g _23672_ (.A(_09468_), .B(_02893_), .Y(_02953_));
NAND_g _23673_ (.A(cpuregs[17][29]), .B(_02894_), .Y(_02954_));
NAND_g _23674_ (.A(_02953_), .B(_02954_), .Y(_00967_));
NAND_g _23675_ (.A(_09481_), .B(_02893_), .Y(_02955_));
NAND_g _23676_ (.A(cpuregs[17][30]), .B(_02894_), .Y(_02956_));
NAND_g _23677_ (.A(_02955_), .B(_02956_), .Y(_00968_));
NAND_g _23678_ (.A(_09493_), .B(_02893_), .Y(_02957_));
NAND_g _23679_ (.A(cpuregs[17][31]), .B(_02894_), .Y(_02958_));
NAND_g _23680_ (.A(_02957_), .B(_02958_), .Y(_00969_));
NAND_g _23681_ (.A(_14393_), .B(_00426_), .Y(_02959_));
NAND_g _23682_ (.A(decoded_imm_j[12]), .B(_14394_), .Y(_02960_));
NAND_g _23683_ (.A(_02959_), .B(_02960_), .Y(_00970_));
NAND_g _23684_ (.A(_14393_), .B(_00427_), .Y(_02961_));
NAND_g _23685_ (.A(decoded_imm_j[13]), .B(_14394_), .Y(_02962_));
NAND_g _23686_ (.A(_02961_), .B(_02962_), .Y(_00971_));
NOR_g _23687_ (.A(decoded_imm_j[14]), .B(_14393_), .Y(_02963_));
NOR_g _23688_ (.A(_14457_), .B(_02963_), .Y(_00972_));
NAND_g _23689_ (.A(_14393_), .B(_00429_), .Y(_02964_));
NAND_g _23690_ (.A(decoded_imm_j[15]), .B(_14394_), .Y(_02965_));
NAND_g _23691_ (.A(_02964_), .B(_02965_), .Y(_00973_));
NAND_g _23692_ (.A(_14393_), .B(_00430_), .Y(_02966_));
NAND_g _23693_ (.A(decoded_imm_j[16]), .B(_14394_), .Y(_02967_));
NAND_g _23694_ (.A(_02966_), .B(_02967_), .Y(_00974_));
NAND_g _23695_ (.A(_14393_), .B(_00431_), .Y(_02968_));
NAND_g _23696_ (.A(decoded_imm_j[17]), .B(_14394_), .Y(_02969_));
NAND_g _23697_ (.A(_02968_), .B(_02969_), .Y(_00975_));
NAND_g _23698_ (.A(_14393_), .B(_00432_), .Y(_02970_));
NAND_g _23699_ (.A(decoded_imm_j[18]), .B(_14394_), .Y(_02971_));
NAND_g _23700_ (.A(_02970_), .B(_02971_), .Y(_00976_));
NAND_g _23701_ (.A(_14393_), .B(_00433_), .Y(_02972_));
NAND_g _23702_ (.A(decoded_imm_j[19]), .B(_14394_), .Y(_02973_));
NAND_g _23703_ (.A(_02972_), .B(_02973_), .Y(_00977_));
NAND_g _23704_ (.A(_10595_), .B(_13863_), .Y(_02974_));
AND_g _23705_ (.A(_10601_), .B(_14353_), .Y(_02975_));
NAND_g _23706_ (.A(_14479_), .B(_02975_), .Y(_02976_));
NOT_g _23707_ (.A(_02976_), .Y(_02977_));
NAND_g _23708_ (.A(_13850_), .B(_13860_), .Y(_02978_));
NAND_g _23709_ (.A(_02976_), .B(_02978_), .Y(_02979_));
NAND_g _23710_ (.A(cpu_state[0]), .B(_02979_), .Y(_02980_));
NAND_g _23711_ (.A(_02974_), .B(_02980_), .Y(_02981_));
NOR_g _23712_ (.A(reg_next_pc[0]), .B(reg_pc[1]), .Y(_02982_));
NOT_g _23713_ (.A(_02982_), .Y(_02983_));
NAND_g _23714_ (.A(mem_do_rinst), .B(_02983_), .Y(_02984_));
NAND_g _23715_ (.A(mem_wordsize[0]), .B(_08961_), .Y(_02985_));
NOR_g _23716_ (.A(mem_wordsize[1]), .B(_14264_), .Y(_02986_));
AND_g _23717_ (.A(_02985_), .B(_02986_), .Y(_02987_));
NAND_g _23718_ (.A(_01777_), .B(_02987_), .Y(_02988_));
NAND_g _23719_ (.A(_02984_), .B(_02988_), .Y(_02989_));
NOR_g _23720_ (.A(_08811_), .B(_02989_), .Y(_02990_));
AND_g _23721_ (.A(_02981_), .B(_02990_), .Y(_00978_));
NAND_g _23722_ (.A(is_sb_sh_sw), .B(_11169_), .Y(_02991_));
NAND_g _23723_ (.A(_13850_), .B(_13857_), .Y(_02992_));
NAND_g _23724_ (.A(cpu_state[1]), .B(_02977_), .Y(_02993_));
AND_g _23725_ (.A(_02992_), .B(_02993_), .Y(_02994_));
NAND_g _23726_ (.A(_02991_), .B(_02994_), .Y(_02995_));
AND_g _23727_ (.A(_02990_), .B(_02995_), .Y(_00979_));
NAND_g _23728_ (.A(is_sll_srl_sra), .B(_11169_), .Y(_02996_));
AND_g _23729_ (.A(is_slli_srli_srai), .B(_10595_), .Y(_02997_));
NAND_g _23730_ (.A(_13884_), .B(_02976_), .Y(_02998_));
AND_g _23731_ (.A(cpu_state[2]), .B(_02998_), .Y(_02999_));
NOR_g _23732_ (.A(_02997_), .B(_02999_), .Y(_03000_));
NAND_g _23733_ (.A(_02996_), .B(_03000_), .Y(_03001_));
AND_g _23734_ (.A(_02990_), .B(_03001_), .Y(_00980_));
NOR_g _23735_ (.A(is_sll_srl_sra), .B(is_sb_sh_sw), .Y(_03002_));
NOR_g _23736_ (.A(_10599_), .B(_10753_), .Y(_03003_));
NOT_g _23737_ (.A(_03003_), .Y(_03004_));
NAND_g _23738_ (.A(_03002_), .B(_03004_), .Y(_03005_));
NAND_g _23739_ (.A(_13848_), .B(_14221_), .Y(_03006_));
NAND_g _23740_ (.A(_02976_), .B(_03006_), .Y(_03007_));
AND_g _23741_ (.A(cpu_state[3]), .B(_03007_), .Y(_03008_));
NOR_g _23742_ (.A(_10606_), .B(_03008_), .Y(_03009_));
NAND_g _23743_ (.A(_03005_), .B(_03009_), .Y(_03010_));
AND_g _23744_ (.A(_02990_), .B(_03010_), .Y(_00981_));
NAND_g _23745_ (.A(cpu_state[4]), .B(_02990_), .Y(_03011_));
NOR_g _23746_ (.A(_02976_), .B(_03011_), .Y(_00982_));
NAND_g _23747_ (.A(_09074_), .B(_02976_), .Y(_03012_));
NOR_g _23748_ (.A(cpu_state[5]), .B(_09894_), .Y(_03013_));
NAND_g _23749_ (.A(_02990_), .B(_03012_), .Y(_03014_));
NOR_g _23750_ (.A(_03013_), .B(_03014_), .Y(_00983_));
NAND_g _23751_ (.A(resetn), .B(_02989_), .Y(_03015_));
NAND_g _23752_ (.A(cpu_state[6]), .B(_02977_), .Y(_03016_));
AND_g _23753_ (.A(resetn), .B(_13891_), .Y(_03017_));
NAND_g _23754_ (.A(_14355_), .B(_03017_), .Y(_03018_));
NOR_g _23755_ (.A(_13889_), .B(_03018_), .Y(_03019_));
AND_g _23756_ (.A(_13861_), .B(_03019_), .Y(_03020_));
NAND_g _23757_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(_13848_), .Y(_03021_));
NAND_g _23758_ (.A(_14214_), .B(_03021_), .Y(_03022_));
AND_g _23759_ (.A(_03020_), .B(_03022_), .Y(_03023_));
NAND_g _23760_ (.A(_03016_), .B(_03023_), .Y(_03024_));
AND_g _23761_ (.A(_03015_), .B(_03024_), .Y(_00984_));
AND_g _23762_ (.A(resetn), .B(_10595_), .Y(_03025_));
NAND_g _23763_ (.A(_10749_), .B(_03025_), .Y(_03026_));
AND_g _23764_ (.A(_09822_), .B(_03015_), .Y(_03027_));
NAND_g _23765_ (.A(_03026_), .B(_03027_), .Y(_00985_));
AND_g _23766_ (.A(_09825_), .B(_02494_), .Y(_03028_));
NAND_g _23767_ (.A(_09825_), .B(_02494_), .Y(_03029_));
NAND_g _23768_ (.A(_09098_), .B(_03028_), .Y(_03030_));
NAND_g _23769_ (.A(cpuregs[5][0]), .B(_03029_), .Y(_03031_));
NAND_g _23770_ (.A(_03030_), .B(_03031_), .Y(_00986_));
NAND_g _23771_ (.A(_09109_), .B(_03028_), .Y(_03032_));
NAND_g _23772_ (.A(cpuregs[5][1]), .B(_03029_), .Y(_03033_));
NAND_g _23773_ (.A(_03032_), .B(_03033_), .Y(_00987_));
NAND_g _23774_ (.A(_09118_), .B(_03028_), .Y(_03034_));
NAND_g _23775_ (.A(cpuregs[5][2]), .B(_03029_), .Y(_03035_));
NAND_g _23776_ (.A(_03034_), .B(_03035_), .Y(_00988_));
NAND_g _23777_ (.A(_09131_), .B(_03028_), .Y(_03036_));
NAND_g _23778_ (.A(cpuregs[5][3]), .B(_03029_), .Y(_03037_));
NAND_g _23779_ (.A(_03036_), .B(_03037_), .Y(_00989_));
NAND_g _23780_ (.A(_09144_), .B(_03028_), .Y(_03038_));
NAND_g _23781_ (.A(cpuregs[5][4]), .B(_03029_), .Y(_03039_));
NAND_g _23782_ (.A(_03038_), .B(_03039_), .Y(_00990_));
NAND_g _23783_ (.A(_09157_), .B(_03028_), .Y(_03040_));
NAND_g _23784_ (.A(cpuregs[5][5]), .B(_03029_), .Y(_03041_));
NAND_g _23785_ (.A(_03040_), .B(_03041_), .Y(_00991_));
NAND_g _23786_ (.A(_09170_), .B(_03028_), .Y(_03042_));
NAND_g _23787_ (.A(cpuregs[5][6]), .B(_03029_), .Y(_03043_));
NAND_g _23788_ (.A(_03042_), .B(_03043_), .Y(_00992_));
NAND_g _23789_ (.A(_09183_), .B(_03028_), .Y(_03044_));
NAND_g _23790_ (.A(cpuregs[5][7]), .B(_03029_), .Y(_03045_));
NAND_g _23791_ (.A(_03044_), .B(_03045_), .Y(_00993_));
NAND_g _23792_ (.A(_09196_), .B(_03028_), .Y(_03046_));
NAND_g _23793_ (.A(cpuregs[5][8]), .B(_03029_), .Y(_03047_));
NAND_g _23794_ (.A(_03046_), .B(_03047_), .Y(_00994_));
NAND_g _23795_ (.A(_09209_), .B(_03028_), .Y(_03048_));
NAND_g _23796_ (.A(cpuregs[5][9]), .B(_03029_), .Y(_03049_));
NAND_g _23797_ (.A(_03048_), .B(_03049_), .Y(_00995_));
NAND_g _23798_ (.A(_09222_), .B(_03028_), .Y(_03050_));
NAND_g _23799_ (.A(cpuregs[5][10]), .B(_03029_), .Y(_03051_));
NAND_g _23800_ (.A(_03050_), .B(_03051_), .Y(_00996_));
NAND_g _23801_ (.A(_09235_), .B(_03028_), .Y(_03052_));
NAND_g _23802_ (.A(cpuregs[5][11]), .B(_03029_), .Y(_03053_));
NAND_g _23803_ (.A(_03052_), .B(_03053_), .Y(_00997_));
NAND_g _23804_ (.A(_09248_), .B(_03028_), .Y(_03054_));
NAND_g _23805_ (.A(cpuregs[5][12]), .B(_03029_), .Y(_03055_));
NAND_g _23806_ (.A(_03054_), .B(_03055_), .Y(_00998_));
NAND_g _23807_ (.A(_09261_), .B(_03028_), .Y(_03056_));
NAND_g _23808_ (.A(cpuregs[5][13]), .B(_03029_), .Y(_03057_));
NAND_g _23809_ (.A(_03056_), .B(_03057_), .Y(_00999_));
NAND_g _23810_ (.A(_09274_), .B(_03028_), .Y(_03058_));
NAND_g _23811_ (.A(cpuregs[5][14]), .B(_03029_), .Y(_03059_));
NAND_g _23812_ (.A(_03058_), .B(_03059_), .Y(_01000_));
NAND_g _23813_ (.A(_09287_), .B(_03028_), .Y(_03060_));
NAND_g _23814_ (.A(cpuregs[5][15]), .B(_03029_), .Y(_03061_));
NAND_g _23815_ (.A(_03060_), .B(_03061_), .Y(_01001_));
NAND_g _23816_ (.A(_09300_), .B(_03028_), .Y(_03062_));
NAND_g _23817_ (.A(cpuregs[5][16]), .B(_03029_), .Y(_03063_));
NAND_g _23818_ (.A(_03062_), .B(_03063_), .Y(_01002_));
NOR_g _23819_ (.A(cpuregs[5][17]), .B(_03028_), .Y(_03064_));
NOR_g _23820_ (.A(_09313_), .B(_03029_), .Y(_03065_));
NOR_g _23821_ (.A(_03064_), .B(_03065_), .Y(_01003_));
AND_g _23822_ (.A(_08955_), .B(_03029_), .Y(_03066_));
NOR_g _23823_ (.A(_09325_), .B(_03029_), .Y(_03067_));
NOR_g _23824_ (.A(_03066_), .B(_03067_), .Y(_01004_));
NAND_g _23825_ (.A(_09338_), .B(_03028_), .Y(_03068_));
NAND_g _23826_ (.A(cpuregs[5][19]), .B(_03029_), .Y(_03069_));
NAND_g _23827_ (.A(_03068_), .B(_03069_), .Y(_01005_));
NAND_g _23828_ (.A(_09351_), .B(_03028_), .Y(_03070_));
NAND_g _23829_ (.A(cpuregs[5][20]), .B(_03029_), .Y(_03071_));
NAND_g _23830_ (.A(_03070_), .B(_03071_), .Y(_01006_));
NAND_g _23831_ (.A(_09364_), .B(_03028_), .Y(_03072_));
NAND_g _23832_ (.A(cpuregs[5][21]), .B(_03029_), .Y(_03073_));
NAND_g _23833_ (.A(_03072_), .B(_03073_), .Y(_01007_));
NAND_g _23834_ (.A(_09377_), .B(_03028_), .Y(_03074_));
NAND_g _23835_ (.A(cpuregs[5][22]), .B(_03029_), .Y(_03075_));
NAND_g _23836_ (.A(_03074_), .B(_03075_), .Y(_01008_));
NAND_g _23837_ (.A(_09390_), .B(_03028_), .Y(_03076_));
NAND_g _23838_ (.A(cpuregs[5][23]), .B(_03029_), .Y(_03077_));
NAND_g _23839_ (.A(_03076_), .B(_03077_), .Y(_01009_));
NAND_g _23840_ (.A(_09403_), .B(_03028_), .Y(_03078_));
NAND_g _23841_ (.A(cpuregs[5][24]), .B(_03029_), .Y(_03079_));
NAND_g _23842_ (.A(_03078_), .B(_03079_), .Y(_01010_));
NAND_g _23843_ (.A(_09416_), .B(_03028_), .Y(_03080_));
NAND_g _23844_ (.A(cpuregs[5][25]), .B(_03029_), .Y(_03081_));
NAND_g _23845_ (.A(_03080_), .B(_03081_), .Y(_01011_));
NAND_g _23846_ (.A(_09429_), .B(_03028_), .Y(_03082_));
NAND_g _23847_ (.A(cpuregs[5][26]), .B(_03029_), .Y(_03083_));
NAND_g _23848_ (.A(_03082_), .B(_03083_), .Y(_01012_));
NAND_g _23849_ (.A(_09442_), .B(_03028_), .Y(_03084_));
NAND_g _23850_ (.A(cpuregs[5][27]), .B(_03029_), .Y(_03085_));
NAND_g _23851_ (.A(_03084_), .B(_03085_), .Y(_01013_));
NAND_g _23852_ (.A(_09455_), .B(_03028_), .Y(_03086_));
NAND_g _23853_ (.A(cpuregs[5][28]), .B(_03029_), .Y(_03087_));
NAND_g _23854_ (.A(_03086_), .B(_03087_), .Y(_01014_));
NAND_g _23855_ (.A(_09468_), .B(_03028_), .Y(_03088_));
NAND_g _23856_ (.A(cpuregs[5][29]), .B(_03029_), .Y(_03089_));
NAND_g _23857_ (.A(_03088_), .B(_03089_), .Y(_01015_));
NAND_g _23858_ (.A(_09481_), .B(_03028_), .Y(_03090_));
NAND_g _23859_ (.A(cpuregs[5][30]), .B(_03029_), .Y(_03091_));
NAND_g _23860_ (.A(_03090_), .B(_03091_), .Y(_01016_));
NAND_g _23861_ (.A(_09493_), .B(_03028_), .Y(_03092_));
NAND_g _23862_ (.A(cpuregs[5][31]), .B(_03029_), .Y(_03093_));
NAND_g _23863_ (.A(_03092_), .B(_03093_), .Y(_01017_));
NOR_g _23864_ (.A(pcpi_rs1[0]), .B(_14488_), .Y(_03094_));
NAND_g _23865_ (.A(reg_next_pc[0]), .B(_14617_), .Y(_03095_));
NAND_g _23866_ (.A(_08963_), .B(_00008_[2]), .Y(_03096_));
NOR_g _23867_ (.A(cpuregs[3][0]), .B(_00008_[2]), .Y(_03097_));
NOR_g _23868_ (.A(_09030_), .B(_03097_), .Y(_03098_));
NAND_g _23869_ (.A(_03096_), .B(_03098_), .Y(_03099_));
NOR_g _23870_ (.A(cpuregs[2][0]), .B(_00008_[2]), .Y(_03100_));
AND_g _23871_ (.A(_09003_), .B(_00008_[2]), .Y(_03101_));
NOR_g _23872_ (.A(_03100_), .B(_03101_), .Y(_03102_));
NAND_g _23873_ (.A(_09030_), .B(_03102_), .Y(_03103_));
NAND_g _23874_ (.A(_03099_), .B(_03103_), .Y(_03104_));
NAND_g _23875_ (.A(_00008_[1]), .B(_03104_), .Y(_03105_));
NAND_g _23876_ (.A(_08946_), .B(_00008_[2]), .Y(_03106_));
NOR_g _23877_ (.A(cpuregs[1][0]), .B(_00008_[2]), .Y(_03107_));
NOR_g _23878_ (.A(_09030_), .B(_03107_), .Y(_03108_));
NAND_g _23879_ (.A(_03106_), .B(_03108_), .Y(_03109_));
NOR_g _23880_ (.A(cpuregs[0][0]), .B(_00008_[2]), .Y(_03110_));
AND_g _23881_ (.A(_08904_), .B(_00008_[2]), .Y(_03111_));
NOR_g _23882_ (.A(_03110_), .B(_03111_), .Y(_03112_));
NAND_g _23883_ (.A(_09030_), .B(_03112_), .Y(_03113_));
NAND_g _23884_ (.A(_03109_), .B(_03113_), .Y(_03114_));
NAND_g _23885_ (.A(_09031_), .B(_03114_), .Y(_03115_));
NAND_g _23886_ (.A(_03105_), .B(_03115_), .Y(_03116_));
NAND_g _23887_ (.A(_09033_), .B(_03116_), .Y(_03117_));
NAND_g _23888_ (.A(cpuregs[13][0]), .B(_00008_[0]), .Y(_03118_));
NAND_g _23889_ (.A(cpuregs[12][0]), .B(_09030_), .Y(_03119_));
AND_g _23890_ (.A(_00008_[2]), .B(_03119_), .Y(_03120_));
NAND_g _23891_ (.A(_03118_), .B(_03120_), .Y(_03121_));
NAND_g _23892_ (.A(cpuregs[9][0]), .B(_00008_[0]), .Y(_03122_));
NAND_g _23893_ (.A(cpuregs[8][0]), .B(_09030_), .Y(_03123_));
AND_g _23894_ (.A(_09032_), .B(_03123_), .Y(_03124_));
NAND_g _23895_ (.A(_03122_), .B(_03124_), .Y(_03125_));
AND_g _23896_ (.A(_09031_), .B(_03125_), .Y(_03126_));
NAND_g _23897_ (.A(_03121_), .B(_03126_), .Y(_03127_));
NAND_g _23898_ (.A(cpuregs[15][0]), .B(_00008_[0]), .Y(_03128_));
NAND_g _23899_ (.A(cpuregs[14][0]), .B(_09030_), .Y(_03129_));
AND_g _23900_ (.A(_00008_[2]), .B(_03129_), .Y(_03130_));
NAND_g _23901_ (.A(_03128_), .B(_03130_), .Y(_03131_));
NAND_g _23902_ (.A(cpuregs[11][0]), .B(_00008_[0]), .Y(_03132_));
NAND_g _23903_ (.A(cpuregs[10][0]), .B(_09030_), .Y(_03133_));
AND_g _23904_ (.A(_09032_), .B(_03133_), .Y(_03134_));
NAND_g _23905_ (.A(_03132_), .B(_03134_), .Y(_03135_));
AND_g _23906_ (.A(_00008_[1]), .B(_03135_), .Y(_03136_));
NAND_g _23907_ (.A(_03131_), .B(_03136_), .Y(_03137_));
NAND_g _23908_ (.A(_03127_), .B(_03137_), .Y(_03138_));
AND_g _23909_ (.A(_00008_[3]), .B(_03138_), .Y(_03139_));
NOR_g _23910_ (.A(_00008_[4]), .B(_03139_), .Y(_03140_));
NAND_g _23911_ (.A(_03117_), .B(_03140_), .Y(_03141_));
NAND_g _23912_ (.A(cpuregs[26][0]), .B(_09032_), .Y(_03142_));
NAND_g _23913_ (.A(cpuregs[30][0]), .B(_00008_[2]), .Y(_03143_));
AND_g _23914_ (.A(_09030_), .B(_03143_), .Y(_03144_));
NAND_g _23915_ (.A(_03142_), .B(_03144_), .Y(_03145_));
NAND_g _23916_ (.A(cpuregs[31][0]), .B(_00008_[2]), .Y(_03146_));
NAND_g _23917_ (.A(cpuregs[27][0]), .B(_09032_), .Y(_03147_));
AND_g _23918_ (.A(_00008_[0]), .B(_03147_), .Y(_03148_));
NAND_g _23919_ (.A(_03146_), .B(_03148_), .Y(_03149_));
NAND_g _23920_ (.A(_03145_), .B(_03149_), .Y(_03150_));
NAND_g _23921_ (.A(_00008_[3]), .B(_03150_), .Y(_03151_));
NAND_g _23922_ (.A(cpuregs[18][0]), .B(_09032_), .Y(_03152_));
NAND_g _23923_ (.A(cpuregs[22][0]), .B(_00008_[2]), .Y(_03153_));
AND_g _23924_ (.A(_09030_), .B(_03153_), .Y(_03154_));
NAND_g _23925_ (.A(_03152_), .B(_03154_), .Y(_03155_));
NAND_g _23926_ (.A(cpuregs[19][0]), .B(_09032_), .Y(_03156_));
NAND_g _23927_ (.A(cpuregs[23][0]), .B(_00008_[2]), .Y(_03157_));
AND_g _23928_ (.A(_00008_[0]), .B(_03157_), .Y(_03158_));
NAND_g _23929_ (.A(_03156_), .B(_03158_), .Y(_03159_));
NAND_g _23930_ (.A(_03155_), .B(_03159_), .Y(_03160_));
NAND_g _23931_ (.A(_09033_), .B(_03160_), .Y(_03161_));
AND_g _23932_ (.A(_03151_), .B(_03161_), .Y(_03162_));
NAND_g _23933_ (.A(cpuregs[24][0]), .B(_09032_), .Y(_03163_));
NAND_g _23934_ (.A(cpuregs[28][0]), .B(_00008_[2]), .Y(_03164_));
AND_g _23935_ (.A(_09030_), .B(_03164_), .Y(_03165_));
NAND_g _23936_ (.A(_03163_), .B(_03165_), .Y(_03166_));
NAND_g _23937_ (.A(cpuregs[29][0]), .B(_00008_[2]), .Y(_03167_));
NAND_g _23938_ (.A(cpuregs[25][0]), .B(_09032_), .Y(_03168_));
AND_g _23939_ (.A(_00008_[0]), .B(_03168_), .Y(_03169_));
NAND_g _23940_ (.A(_03167_), .B(_03169_), .Y(_03170_));
NAND_g _23941_ (.A(_03166_), .B(_03170_), .Y(_03171_));
NAND_g _23942_ (.A(_00008_[3]), .B(_03171_), .Y(_03172_));
NAND_g _23943_ (.A(cpuregs[16][0]), .B(_09032_), .Y(_03173_));
NAND_g _23944_ (.A(cpuregs[20][0]), .B(_00008_[2]), .Y(_03174_));
AND_g _23945_ (.A(_09030_), .B(_03174_), .Y(_03175_));
NAND_g _23946_ (.A(_03173_), .B(_03175_), .Y(_03176_));
NAND_g _23947_ (.A(cpuregs[17][0]), .B(_09032_), .Y(_03177_));
NAND_g _23948_ (.A(cpuregs[21][0]), .B(_00008_[2]), .Y(_03178_));
AND_g _23949_ (.A(_00008_[0]), .B(_03178_), .Y(_03179_));
NAND_g _23950_ (.A(_03177_), .B(_03179_), .Y(_03180_));
NAND_g _23951_ (.A(_03176_), .B(_03180_), .Y(_03181_));
NAND_g _23952_ (.A(_09033_), .B(_03181_), .Y(_03182_));
AND_g _23953_ (.A(_03172_), .B(_03182_), .Y(_03183_));
NAND_g _23954_ (.A(_00008_[1]), .B(_03162_), .Y(_03184_));
NAND_g _23955_ (.A(_09031_), .B(_03183_), .Y(_03185_));
AND_g _23956_ (.A(_00008_[4]), .B(_03184_), .Y(_03186_));
NAND_g _23957_ (.A(_03185_), .B(_03186_), .Y(_03187_));
AND_g _23958_ (.A(_03141_), .B(_03187_), .Y(_03188_));
NAND_g _23959_ (.A(_14624_), .B(_03188_), .Y(_03189_));
NAND_g _23960_ (.A(_03095_), .B(_03189_), .Y(_03190_));
NAND_g _23961_ (.A(_10595_), .B(_03190_), .Y(_03191_));
NAND_g _23962_ (.A(pcpi_rs1[4]), .B(_13880_), .Y(_03192_));
NAND_g _23963_ (.A(pcpi_rs1[1]), .B(_13879_), .Y(_03193_));
NAND_g _23964_ (.A(_03192_), .B(_03193_), .Y(_03194_));
AND_g _23965_ (.A(_14482_), .B(_03194_), .Y(_03195_));
AND_g _23966_ (.A(_13883_), .B(_03195_), .Y(_03196_));
NOR_g _23967_ (.A(decoded_imm[0]), .B(pcpi_rs1[0]), .Y(_03197_));
NAND_g _23968_ (.A(_14549_), .B(_14614_), .Y(_03198_));
AND_g _23969_ (.A(_14488_), .B(_03198_), .Y(_03199_));
NOR_g _23970_ (.A(_03197_), .B(_03199_), .Y(_03200_));
NOR_g _23971_ (.A(_03196_), .B(_03200_), .Y(_03201_));
AND_g _23972_ (.A(_03191_), .B(_03201_), .Y(_03202_));
NOR_g _23973_ (.A(_03094_), .B(_03202_), .Y(_01018_));
NAND_g _23974_ (.A(reg_pc[1]), .B(_14617_), .Y(_03203_));
NAND_g _23975_ (.A(cpuregs[22][1]), .B(_00008_[2]), .Y(_03204_));
NAND_g _23976_ (.A(cpuregs[18][1]), .B(_09032_), .Y(_03205_));
AND_g _23977_ (.A(_03204_), .B(_03205_), .Y(_03206_));
NOR_g _23978_ (.A(_00008_[0]), .B(_03206_), .Y(_03207_));
NAND_g _23979_ (.A(_08885_), .B(_00008_[2]), .Y(_03208_));
NOR_g _23980_ (.A(cpuregs[19][1]), .B(_00008_[2]), .Y(_03209_));
NOR_g _23981_ (.A(_09030_), .B(_03209_), .Y(_03210_));
AND_g _23982_ (.A(_03208_), .B(_03210_), .Y(_03211_));
NOR_g _23983_ (.A(_03207_), .B(_03211_), .Y(_03212_));
NAND_g _23984_ (.A(_00008_[1]), .B(_03212_), .Y(_03213_));
NAND_g _23985_ (.A(cpuregs[20][1]), .B(_00008_[2]), .Y(_03214_));
NAND_g _23986_ (.A(cpuregs[16][1]), .B(_09032_), .Y(_03215_));
AND_g _23987_ (.A(_03214_), .B(_03215_), .Y(_03216_));
NOR_g _23988_ (.A(_00008_[0]), .B(_03216_), .Y(_03217_));
NAND_g _23989_ (.A(_08982_), .B(_00008_[2]), .Y(_03218_));
NOR_g _23990_ (.A(cpuregs[17][1]), .B(_00008_[2]), .Y(_03219_));
NOR_g _23991_ (.A(_09030_), .B(_03219_), .Y(_03220_));
NAND_g _23992_ (.A(_03218_), .B(_03220_), .Y(_03221_));
NAND_g _23993_ (.A(_09031_), .B(_03221_), .Y(_03222_));
NOR_g _23994_ (.A(_03217_), .B(_03222_), .Y(_03223_));
NAND_g _23995_ (.A(cpuregs[27][1]), .B(_00008_[0]), .Y(_03224_));
NAND_g _23996_ (.A(cpuregs[26][1]), .B(_09030_), .Y(_03225_));
AND_g _23997_ (.A(_09032_), .B(_03225_), .Y(_03226_));
NAND_g _23998_ (.A(_03224_), .B(_03226_), .Y(_03227_));
NAND_g _23999_ (.A(cpuregs[31][1]), .B(_00008_[0]), .Y(_03228_));
NAND_g _24000_ (.A(cpuregs[30][1]), .B(_09030_), .Y(_03229_));
AND_g _24001_ (.A(_00008_[2]), .B(_03229_), .Y(_03230_));
NAND_g _24002_ (.A(_03228_), .B(_03230_), .Y(_03231_));
NAND_g _24003_ (.A(_03227_), .B(_03231_), .Y(_03232_));
NAND_g _24004_ (.A(_00008_[1]), .B(_03232_), .Y(_03233_));
NAND_g _24005_ (.A(cpuregs[25][1]), .B(_00008_[0]), .Y(_03234_));
NAND_g _24006_ (.A(cpuregs[24][1]), .B(_09030_), .Y(_03235_));
AND_g _24007_ (.A(_09032_), .B(_03235_), .Y(_03236_));
NAND_g _24008_ (.A(_03234_), .B(_03236_), .Y(_03237_));
NAND_g _24009_ (.A(cpuregs[29][1]), .B(_00008_[0]), .Y(_03238_));
NAND_g _24010_ (.A(cpuregs[28][1]), .B(_09030_), .Y(_03239_));
AND_g _24011_ (.A(_00008_[2]), .B(_03239_), .Y(_03240_));
NAND_g _24012_ (.A(_03238_), .B(_03240_), .Y(_03241_));
NAND_g _24013_ (.A(_03237_), .B(_03241_), .Y(_03242_));
NAND_g _24014_ (.A(_09031_), .B(_03242_), .Y(_03243_));
AND_g _24015_ (.A(_00008_[3]), .B(_03233_), .Y(_03244_));
NAND_g _24016_ (.A(_03243_), .B(_03244_), .Y(_03245_));
NOR_g _24017_ (.A(_00008_[3]), .B(_03223_), .Y(_03246_));
NAND_g _24018_ (.A(_03213_), .B(_03246_), .Y(_03247_));
AND_g _24019_ (.A(_00008_[4]), .B(_03247_), .Y(_03248_));
AND_g _24020_ (.A(_03245_), .B(_03248_), .Y(_03249_));
NAND_g _24021_ (.A(cpuregs[9][1]), .B(_09032_), .Y(_03250_));
NAND_g _24022_ (.A(cpuregs[13][1]), .B(_00008_[2]), .Y(_03251_));
AND_g _24023_ (.A(_09031_), .B(_03251_), .Y(_03252_));
NAND_g _24024_ (.A(_03250_), .B(_03252_), .Y(_03253_));
NAND_g _24025_ (.A(cpuregs[15][1]), .B(_00008_[2]), .Y(_03254_));
NAND_g _24026_ (.A(cpuregs[11][1]), .B(_09032_), .Y(_03255_));
AND_g _24027_ (.A(_00008_[1]), .B(_03255_), .Y(_03256_));
NAND_g _24028_ (.A(_03254_), .B(_03256_), .Y(_03257_));
NAND_g _24029_ (.A(_03253_), .B(_03257_), .Y(_03258_));
NAND_g _24030_ (.A(_00008_[0]), .B(_03258_), .Y(_03259_));
NAND_g _24031_ (.A(cpuregs[8][1]), .B(_09032_), .Y(_03260_));
NAND_g _24032_ (.A(cpuregs[12][1]), .B(_00008_[2]), .Y(_03261_));
AND_g _24033_ (.A(_09031_), .B(_03261_), .Y(_03262_));
NAND_g _24034_ (.A(_03260_), .B(_03262_), .Y(_03263_));
NAND_g _24035_ (.A(cpuregs[10][1]), .B(_09032_), .Y(_03264_));
NAND_g _24036_ (.A(cpuregs[14][1]), .B(_00008_[2]), .Y(_03265_));
AND_g _24037_ (.A(_00008_[1]), .B(_03265_), .Y(_03266_));
NAND_g _24038_ (.A(_03264_), .B(_03266_), .Y(_03267_));
NAND_g _24039_ (.A(_03263_), .B(_03267_), .Y(_03268_));
NAND_g _24040_ (.A(_09030_), .B(_03268_), .Y(_03269_));
NAND_g _24041_ (.A(_03259_), .B(_03269_), .Y(_03270_));
NAND_g _24042_ (.A(_00008_[3]), .B(_03270_), .Y(_03271_));
NAND_g _24043_ (.A(cpuregs[1][1]), .B(_09031_), .Y(_03272_));
NAND_g _24044_ (.A(cpuregs[3][1]), .B(_00008_[1]), .Y(_03273_));
AND_g _24045_ (.A(_09032_), .B(_03273_), .Y(_03274_));
NAND_g _24046_ (.A(_03272_), .B(_03274_), .Y(_03275_));
NAND_g _24047_ (.A(cpuregs[5][1]), .B(_09031_), .Y(_03276_));
NAND_g _24048_ (.A(cpuregs[7][1]), .B(_00008_[1]), .Y(_03277_));
AND_g _24049_ (.A(_00008_[2]), .B(_03277_), .Y(_03278_));
NAND_g _24050_ (.A(_03276_), .B(_03278_), .Y(_03279_));
NAND_g _24051_ (.A(_03275_), .B(_03279_), .Y(_03280_));
NAND_g _24052_ (.A(_00008_[0]), .B(_03280_), .Y(_03281_));
NAND_g _24053_ (.A(cpuregs[0][1]), .B(_09031_), .Y(_03282_));
NAND_g _24054_ (.A(cpuregs[2][1]), .B(_00008_[1]), .Y(_03283_));
AND_g _24055_ (.A(_09032_), .B(_03283_), .Y(_03284_));
NAND_g _24056_ (.A(_03282_), .B(_03284_), .Y(_03285_));
NAND_g _24057_ (.A(cpuregs[4][1]), .B(_09031_), .Y(_03286_));
NAND_g _24058_ (.A(cpuregs[6][1]), .B(_00008_[1]), .Y(_03287_));
AND_g _24059_ (.A(_00008_[2]), .B(_03287_), .Y(_03288_));
NAND_g _24060_ (.A(_03286_), .B(_03288_), .Y(_03289_));
NAND_g _24061_ (.A(_03285_), .B(_03289_), .Y(_03290_));
NAND_g _24062_ (.A(_09030_), .B(_03290_), .Y(_03291_));
NAND_g _24063_ (.A(_03281_), .B(_03291_), .Y(_03292_));
NAND_g _24064_ (.A(_09033_), .B(_03292_), .Y(_03293_));
AND_g _24065_ (.A(_03271_), .B(_03293_), .Y(_03294_));
NOR_g _24066_ (.A(_00008_[4]), .B(_03294_), .Y(_03295_));
NOR_g _24067_ (.A(_03249_), .B(_03295_), .Y(_03296_));
NAND_g _24068_ (.A(_14624_), .B(_03296_), .Y(_03297_));
NAND_g _24069_ (.A(_03203_), .B(_03297_), .Y(_03298_));
NAND_g _24070_ (.A(_10595_), .B(_03298_), .Y(_03299_));
XNOR_g _24071_ (.A(_14549_), .B(_14550_), .Y(_03300_));
NAND_g _24072_ (.A(_14614_), .B(_03300_), .Y(_03301_));
NAND_g _24073_ (.A(pcpi_rs1[2]), .B(_14482_), .Y(_03302_));
NAND_g _24074_ (.A(pcpi_rs1[0]), .B(_14481_), .Y(_03303_));
NAND_g _24075_ (.A(pcpi_rs1[5]), .B(_14482_), .Y(_03304_));
AND_g _24076_ (.A(_13879_), .B(_03303_), .Y(_03305_));
NAND_g _24077_ (.A(_03302_), .B(_03305_), .Y(_03306_));
NAND_g _24078_ (.A(_13880_), .B(_03304_), .Y(_03307_));
AND_g _24079_ (.A(_13883_), .B(_03306_), .Y(_03308_));
NAND_g _24080_ (.A(_03307_), .B(_03308_), .Y(_03309_));
AND_g _24081_ (.A(_14488_), .B(_03309_), .Y(_03310_));
AND_g _24082_ (.A(_03301_), .B(_03310_), .Y(_03311_));
AND_g _24083_ (.A(_03299_), .B(_03311_), .Y(_03312_));
NOR_g _24084_ (.A(pcpi_rs1[1]), .B(_14488_), .Y(_03313_));
NOR_g _24085_ (.A(_03312_), .B(_03313_), .Y(_01019_));
NAND_g _24086_ (.A(reg_pc[2]), .B(_14617_), .Y(_03314_));
NAND_g _24087_ (.A(cpuregs[20][2]), .B(_00008_[2]), .Y(_03315_));
NAND_g _24088_ (.A(cpuregs[16][2]), .B(_09032_), .Y(_03316_));
AND_g _24089_ (.A(_03315_), .B(_03316_), .Y(_03317_));
NOR_g _24090_ (.A(_00008_[0]), .B(_03317_), .Y(_03318_));
NAND_g _24091_ (.A(_08983_), .B(_00008_[2]), .Y(_03319_));
NOR_g _24092_ (.A(cpuregs[17][2]), .B(_00008_[2]), .Y(_03320_));
NOR_g _24093_ (.A(_09030_), .B(_03320_), .Y(_03321_));
NAND_g _24094_ (.A(_03319_), .B(_03321_), .Y(_03322_));
NAND_g _24095_ (.A(_09031_), .B(_03322_), .Y(_03323_));
NOR_g _24096_ (.A(_03318_), .B(_03323_), .Y(_03324_));
NAND_g _24097_ (.A(cpuregs[22][2]), .B(_00008_[2]), .Y(_03325_));
NAND_g _24098_ (.A(cpuregs[18][2]), .B(_09032_), .Y(_03326_));
AND_g _24099_ (.A(_03325_), .B(_03326_), .Y(_03327_));
NOR_g _24100_ (.A(_00008_[0]), .B(_03327_), .Y(_03328_));
NAND_g _24101_ (.A(cpuregs[23][2]), .B(_00008_[2]), .Y(_03329_));
NAND_g _24102_ (.A(cpuregs[19][2]), .B(_09032_), .Y(_03330_));
NAND_g _24103_ (.A(_03329_), .B(_03330_), .Y(_03331_));
AND_g _24104_ (.A(_00008_[0]), .B(_03331_), .Y(_03332_));
NOR_g _24105_ (.A(_03328_), .B(_03332_), .Y(_03333_));
NAND_g _24106_ (.A(_00008_[1]), .B(_03333_), .Y(_03334_));
NAND_g _24107_ (.A(cpuregs[27][2]), .B(_00008_[0]), .Y(_03335_));
NAND_g _24108_ (.A(cpuregs[26][2]), .B(_09030_), .Y(_03336_));
AND_g _24109_ (.A(_09032_), .B(_03336_), .Y(_03337_));
NAND_g _24110_ (.A(_03335_), .B(_03337_), .Y(_03338_));
NAND_g _24111_ (.A(cpuregs[31][2]), .B(_00008_[0]), .Y(_03339_));
NAND_g _24112_ (.A(cpuregs[30][2]), .B(_09030_), .Y(_03340_));
AND_g _24113_ (.A(_00008_[2]), .B(_03340_), .Y(_03341_));
NAND_g _24114_ (.A(_03339_), .B(_03341_), .Y(_03342_));
NAND_g _24115_ (.A(_03338_), .B(_03342_), .Y(_03343_));
NAND_g _24116_ (.A(_00008_[1]), .B(_03343_), .Y(_03344_));
NAND_g _24117_ (.A(cpuregs[25][2]), .B(_00008_[0]), .Y(_03345_));
NAND_g _24118_ (.A(cpuregs[24][2]), .B(_09030_), .Y(_03346_));
AND_g _24119_ (.A(_09032_), .B(_03346_), .Y(_03347_));
NAND_g _24120_ (.A(_03345_), .B(_03347_), .Y(_03348_));
NAND_g _24121_ (.A(cpuregs[29][2]), .B(_00008_[0]), .Y(_03349_));
NAND_g _24122_ (.A(cpuregs[28][2]), .B(_09030_), .Y(_03350_));
AND_g _24123_ (.A(_00008_[2]), .B(_03350_), .Y(_03351_));
NAND_g _24124_ (.A(_03349_), .B(_03351_), .Y(_03352_));
NAND_g _24125_ (.A(_03348_), .B(_03352_), .Y(_03353_));
NAND_g _24126_ (.A(_09031_), .B(_03353_), .Y(_03354_));
AND_g _24127_ (.A(_00008_[3]), .B(_03344_), .Y(_03355_));
NAND_g _24128_ (.A(_03354_), .B(_03355_), .Y(_03356_));
NOR_g _24129_ (.A(_00008_[3]), .B(_03324_), .Y(_03357_));
NAND_g _24130_ (.A(_03334_), .B(_03357_), .Y(_03358_));
AND_g _24131_ (.A(_00008_[4]), .B(_03358_), .Y(_03359_));
AND_g _24132_ (.A(_03356_), .B(_03359_), .Y(_03360_));
NAND_g _24133_ (.A(cpuregs[9][2]), .B(_09032_), .Y(_03361_));
NAND_g _24134_ (.A(cpuregs[13][2]), .B(_00008_[2]), .Y(_03362_));
AND_g _24135_ (.A(_09031_), .B(_03362_), .Y(_03363_));
NAND_g _24136_ (.A(_03361_), .B(_03363_), .Y(_03364_));
NAND_g _24137_ (.A(cpuregs[15][2]), .B(_00008_[2]), .Y(_03365_));
NAND_g _24138_ (.A(cpuregs[11][2]), .B(_09032_), .Y(_03366_));
AND_g _24139_ (.A(_00008_[1]), .B(_03366_), .Y(_03367_));
NAND_g _24140_ (.A(_03365_), .B(_03367_), .Y(_03368_));
NAND_g _24141_ (.A(_03364_), .B(_03368_), .Y(_03369_));
NAND_g _24142_ (.A(_00008_[0]), .B(_03369_), .Y(_03370_));
NAND_g _24143_ (.A(cpuregs[8][2]), .B(_09032_), .Y(_03371_));
NAND_g _24144_ (.A(cpuregs[12][2]), .B(_00008_[2]), .Y(_03372_));
AND_g _24145_ (.A(_09031_), .B(_03372_), .Y(_03373_));
NAND_g _24146_ (.A(_03371_), .B(_03373_), .Y(_03374_));
NAND_g _24147_ (.A(cpuregs[10][2]), .B(_09032_), .Y(_03375_));
NAND_g _24148_ (.A(cpuregs[14][2]), .B(_00008_[2]), .Y(_03376_));
AND_g _24149_ (.A(_00008_[1]), .B(_03376_), .Y(_03377_));
NAND_g _24150_ (.A(_03375_), .B(_03377_), .Y(_03378_));
NAND_g _24151_ (.A(_03374_), .B(_03378_), .Y(_03379_));
NAND_g _24152_ (.A(_09030_), .B(_03379_), .Y(_03380_));
NAND_g _24153_ (.A(_03370_), .B(_03380_), .Y(_03381_));
NAND_g _24154_ (.A(_00008_[3]), .B(_03381_), .Y(_03382_));
NAND_g _24155_ (.A(cpuregs[1][2]), .B(_09031_), .Y(_03383_));
NAND_g _24156_ (.A(cpuregs[3][2]), .B(_00008_[1]), .Y(_03384_));
AND_g _24157_ (.A(_09032_), .B(_03384_), .Y(_03385_));
NAND_g _24158_ (.A(_03383_), .B(_03385_), .Y(_03386_));
NAND_g _24159_ (.A(cpuregs[5][2]), .B(_09031_), .Y(_03387_));
NAND_g _24160_ (.A(cpuregs[7][2]), .B(_00008_[1]), .Y(_03388_));
AND_g _24161_ (.A(_00008_[2]), .B(_03388_), .Y(_03389_));
NAND_g _24162_ (.A(_03387_), .B(_03389_), .Y(_03390_));
NAND_g _24163_ (.A(_03386_), .B(_03390_), .Y(_03391_));
NAND_g _24164_ (.A(_00008_[0]), .B(_03391_), .Y(_03392_));
NAND_g _24165_ (.A(cpuregs[0][2]), .B(_09031_), .Y(_03393_));
NAND_g _24166_ (.A(cpuregs[2][2]), .B(_00008_[1]), .Y(_03394_));
AND_g _24167_ (.A(_09032_), .B(_03394_), .Y(_03395_));
NAND_g _24168_ (.A(_03393_), .B(_03395_), .Y(_03396_));
NAND_g _24169_ (.A(cpuregs[4][2]), .B(_09031_), .Y(_03397_));
NAND_g _24170_ (.A(cpuregs[6][2]), .B(_00008_[1]), .Y(_03398_));
AND_g _24171_ (.A(_00008_[2]), .B(_03398_), .Y(_03399_));
NAND_g _24172_ (.A(_03397_), .B(_03399_), .Y(_03400_));
NAND_g _24173_ (.A(_03396_), .B(_03400_), .Y(_03401_));
NAND_g _24174_ (.A(_09030_), .B(_03401_), .Y(_03402_));
NAND_g _24175_ (.A(_03392_), .B(_03402_), .Y(_03403_));
NAND_g _24176_ (.A(_09033_), .B(_03403_), .Y(_03404_));
AND_g _24177_ (.A(_03382_), .B(_03404_), .Y(_03405_));
NOR_g _24178_ (.A(_00008_[4]), .B(_03405_), .Y(_03406_));
NOR_g _24179_ (.A(_03360_), .B(_03406_), .Y(_03407_));
NAND_g _24180_ (.A(_14624_), .B(_03407_), .Y(_03408_));
NAND_g _24181_ (.A(_03314_), .B(_03408_), .Y(_03409_));
NAND_g _24182_ (.A(_10595_), .B(_03409_), .Y(_03410_));
XOR_g _24183_ (.A(_14552_), .B(_14553_), .Y(_03411_));
NAND_g _24184_ (.A(_14614_), .B(_03411_), .Y(_03412_));
NAND_g _24185_ (.A(pcpi_rs1[3]), .B(_14482_), .Y(_03413_));
NAND_g _24186_ (.A(pcpi_rs1[1]), .B(_14481_), .Y(_03414_));
NAND_g _24187_ (.A(pcpi_rs1[6]), .B(_14482_), .Y(_03415_));
AND_g _24188_ (.A(_13879_), .B(_03414_), .Y(_03416_));
NAND_g _24189_ (.A(_03413_), .B(_03416_), .Y(_03417_));
NAND_g _24190_ (.A(_13880_), .B(_03415_), .Y(_03418_));
AND_g _24191_ (.A(_13883_), .B(_03417_), .Y(_03419_));
NAND_g _24192_ (.A(_03418_), .B(_03419_), .Y(_03420_));
AND_g _24193_ (.A(_14488_), .B(_03420_), .Y(_03421_));
AND_g _24194_ (.A(_03412_), .B(_03421_), .Y(_03422_));
AND_g _24195_ (.A(_03410_), .B(_03422_), .Y(_03423_));
NOR_g _24196_ (.A(pcpi_rs1[2]), .B(_14488_), .Y(_03424_));
NOR_g _24197_ (.A(_03423_), .B(_03424_), .Y(_01020_));
NAND_g _24198_ (.A(reg_pc[3]), .B(_14617_), .Y(_03425_));
NAND_g _24199_ (.A(cpuregs[9][3]), .B(_09032_), .Y(_03426_));
NAND_g _24200_ (.A(cpuregs[13][3]), .B(_00008_[2]), .Y(_03427_));
NAND_g _24201_ (.A(_03426_), .B(_03427_), .Y(_03428_));
NAND_g _24202_ (.A(_00008_[0]), .B(_03428_), .Y(_03429_));
NAND_g _24203_ (.A(cpuregs[12][3]), .B(_00008_[2]), .Y(_03430_));
NAND_g _24204_ (.A(cpuregs[8][3]), .B(_09032_), .Y(_03431_));
NAND_g _24205_ (.A(_03430_), .B(_03431_), .Y(_03432_));
NAND_g _24206_ (.A(_09030_), .B(_03432_), .Y(_03433_));
NAND_g _24207_ (.A(_03429_), .B(_03433_), .Y(_03434_));
NAND_g _24208_ (.A(_00008_[3]), .B(_03434_), .Y(_03435_));
NAND_g _24209_ (.A(cpuregs[5][3]), .B(_00008_[2]), .Y(_03436_));
NAND_g _24210_ (.A(cpuregs[1][3]), .B(_09032_), .Y(_03437_));
AND_g _24211_ (.A(_03436_), .B(_03437_), .Y(_03438_));
NAND_g _24212_ (.A(cpuregs[4][3]), .B(_00008_[2]), .Y(_03439_));
NAND_g _24213_ (.A(cpuregs[0][3]), .B(_09032_), .Y(_03440_));
AND_g _24214_ (.A(_03439_), .B(_03440_), .Y(_03441_));
NAND_g _24215_ (.A(_00008_[0]), .B(_03438_), .Y(_03442_));
NAND_g _24216_ (.A(_09030_), .B(_03441_), .Y(_03443_));
AND_g _24217_ (.A(_03442_), .B(_03443_), .Y(_03444_));
NAND_g _24218_ (.A(_09033_), .B(_03444_), .Y(_03445_));
NAND_g _24219_ (.A(_03435_), .B(_03445_), .Y(_03446_));
AND_g _24220_ (.A(_09031_), .B(_03446_), .Y(_03447_));
NAND_g _24221_ (.A(cpuregs[7][3]), .B(_00008_[0]), .Y(_03448_));
NAND_g _24222_ (.A(cpuregs[6][3]), .B(_09030_), .Y(_03449_));
AND_g _24223_ (.A(_00008_[2]), .B(_03449_), .Y(_03450_));
NAND_g _24224_ (.A(_03448_), .B(_03450_), .Y(_03451_));
NAND_g _24225_ (.A(cpuregs[3][3]), .B(_00008_[0]), .Y(_03452_));
NAND_g _24226_ (.A(cpuregs[2][3]), .B(_09030_), .Y(_03453_));
AND_g _24227_ (.A(_09032_), .B(_03453_), .Y(_03454_));
NAND_g _24228_ (.A(_03452_), .B(_03454_), .Y(_03455_));
AND_g _24229_ (.A(_09033_), .B(_03455_), .Y(_03456_));
NAND_g _24230_ (.A(_03451_), .B(_03456_), .Y(_03457_));
NAND_g _24231_ (.A(cpuregs[15][3]), .B(_00008_[0]), .Y(_03458_));
NAND_g _24232_ (.A(cpuregs[14][3]), .B(_09030_), .Y(_03459_));
AND_g _24233_ (.A(_00008_[2]), .B(_03459_), .Y(_03460_));
NAND_g _24234_ (.A(_03458_), .B(_03460_), .Y(_03461_));
NAND_g _24235_ (.A(cpuregs[11][3]), .B(_00008_[0]), .Y(_03462_));
NAND_g _24236_ (.A(cpuregs[10][3]), .B(_09030_), .Y(_03463_));
AND_g _24237_ (.A(_09032_), .B(_03463_), .Y(_03464_));
NAND_g _24238_ (.A(_03462_), .B(_03464_), .Y(_03465_));
AND_g _24239_ (.A(_00008_[3]), .B(_03465_), .Y(_03466_));
NAND_g _24240_ (.A(_03461_), .B(_03466_), .Y(_03467_));
NAND_g _24241_ (.A(_03457_), .B(_03467_), .Y(_03468_));
NAND_g _24242_ (.A(_00008_[1]), .B(_03468_), .Y(_03469_));
NOR_g _24243_ (.A(_00008_[4]), .B(_03447_), .Y(_03470_));
NAND_g _24244_ (.A(_03469_), .B(_03470_), .Y(_03471_));
NAND_g _24245_ (.A(cpuregs[25][3]), .B(_09032_), .Y(_03472_));
NAND_g _24246_ (.A(cpuregs[29][3]), .B(_00008_[2]), .Y(_03473_));
AND_g _24247_ (.A(_09031_), .B(_03473_), .Y(_03474_));
NAND_g _24248_ (.A(_03472_), .B(_03474_), .Y(_03475_));
NAND_g _24249_ (.A(cpuregs[31][3]), .B(_00008_[2]), .Y(_03476_));
NAND_g _24250_ (.A(cpuregs[27][3]), .B(_09032_), .Y(_03477_));
AND_g _24251_ (.A(_00008_[1]), .B(_03477_), .Y(_03478_));
NAND_g _24252_ (.A(_03476_), .B(_03478_), .Y(_03479_));
NAND_g _24253_ (.A(_03475_), .B(_03479_), .Y(_03480_));
NAND_g _24254_ (.A(_00008_[0]), .B(_03480_), .Y(_03481_));
NAND_g _24255_ (.A(cpuregs[24][3]), .B(_09032_), .Y(_03482_));
NAND_g _24256_ (.A(cpuregs[28][3]), .B(_00008_[2]), .Y(_03483_));
AND_g _24257_ (.A(_09031_), .B(_03483_), .Y(_03484_));
NAND_g _24258_ (.A(_03482_), .B(_03484_), .Y(_03485_));
NAND_g _24259_ (.A(cpuregs[26][3]), .B(_09032_), .Y(_03486_));
NAND_g _24260_ (.A(cpuregs[30][3]), .B(_00008_[2]), .Y(_03487_));
AND_g _24261_ (.A(_00008_[1]), .B(_03487_), .Y(_03488_));
NAND_g _24262_ (.A(_03486_), .B(_03488_), .Y(_03489_));
NAND_g _24263_ (.A(_03485_), .B(_03489_), .Y(_03490_));
NAND_g _24264_ (.A(_09030_), .B(_03490_), .Y(_03491_));
NAND_g _24265_ (.A(_03481_), .B(_03491_), .Y(_03492_));
NAND_g _24266_ (.A(_00008_[3]), .B(_03492_), .Y(_03493_));
NAND_g _24267_ (.A(cpuregs[17][3]), .B(_09031_), .Y(_03494_));
NAND_g _24268_ (.A(cpuregs[19][3]), .B(_00008_[1]), .Y(_03495_));
AND_g _24269_ (.A(_09032_), .B(_03495_), .Y(_03496_));
NAND_g _24270_ (.A(_03494_), .B(_03496_), .Y(_03497_));
NAND_g _24271_ (.A(cpuregs[21][3]), .B(_09031_), .Y(_03498_));
NAND_g _24272_ (.A(cpuregs[23][3]), .B(_00008_[1]), .Y(_03499_));
AND_g _24273_ (.A(_00008_[2]), .B(_03499_), .Y(_03500_));
NAND_g _24274_ (.A(_03498_), .B(_03500_), .Y(_03501_));
NAND_g _24275_ (.A(_03497_), .B(_03501_), .Y(_03502_));
NAND_g _24276_ (.A(_00008_[0]), .B(_03502_), .Y(_03503_));
NAND_g _24277_ (.A(cpuregs[16][3]), .B(_09031_), .Y(_03504_));
NAND_g _24278_ (.A(cpuregs[18][3]), .B(_00008_[1]), .Y(_03505_));
AND_g _24279_ (.A(_09032_), .B(_03505_), .Y(_03506_));
NAND_g _24280_ (.A(_03504_), .B(_03506_), .Y(_03507_));
NAND_g _24281_ (.A(cpuregs[20][3]), .B(_09031_), .Y(_03508_));
NAND_g _24282_ (.A(cpuregs[22][3]), .B(_00008_[1]), .Y(_03509_));
AND_g _24283_ (.A(_00008_[2]), .B(_03509_), .Y(_03510_));
NAND_g _24284_ (.A(_03508_), .B(_03510_), .Y(_03511_));
NAND_g _24285_ (.A(_03507_), .B(_03511_), .Y(_03512_));
NAND_g _24286_ (.A(_09030_), .B(_03512_), .Y(_03513_));
NAND_g _24287_ (.A(_03503_), .B(_03513_), .Y(_03514_));
AND_g _24288_ (.A(_09033_), .B(_03514_), .Y(_03515_));
NOT_g _24289_ (.A(_03515_), .Y(_03516_));
NAND_g _24290_ (.A(_03493_), .B(_03516_), .Y(_03517_));
NAND_g _24291_ (.A(_00008_[4]), .B(_03517_), .Y(_03518_));
AND_g _24292_ (.A(_03471_), .B(_03518_), .Y(_03519_));
NAND_g _24293_ (.A(_14624_), .B(_03519_), .Y(_03520_));
NAND_g _24294_ (.A(_03425_), .B(_03520_), .Y(_03521_));
NAND_g _24295_ (.A(_10595_), .B(_03521_), .Y(_03522_));
XOR_g _24296_ (.A(decoded_imm[3]), .B(pcpi_rs1[3]), .Y(_03523_));
XNOR_g _24297_ (.A(_14555_), .B(_03523_), .Y(_03524_));
NAND_g _24298_ (.A(_14614_), .B(_03524_), .Y(_03525_));
NAND_g _24299_ (.A(pcpi_rs1[7]), .B(_14482_), .Y(_03526_));
NAND_g _24300_ (.A(_13880_), .B(_03526_), .Y(_03527_));
NAND_g _24301_ (.A(pcpi_rs1[4]), .B(_14482_), .Y(_03528_));
NAND_g _24302_ (.A(pcpi_rs1[2]), .B(_14481_), .Y(_03529_));
AND_g _24303_ (.A(_13879_), .B(_03528_), .Y(_03530_));
NAND_g _24304_ (.A(_03529_), .B(_03530_), .Y(_03531_));
AND_g _24305_ (.A(_03527_), .B(_03531_), .Y(_03532_));
NAND_g _24306_ (.A(_13883_), .B(_03532_), .Y(_03533_));
AND_g _24307_ (.A(_14488_), .B(_03525_), .Y(_03534_));
AND_g _24308_ (.A(_03533_), .B(_03534_), .Y(_03535_));
AND_g _24309_ (.A(_03522_), .B(_03535_), .Y(_03536_));
NOR_g _24310_ (.A(pcpi_rs1[3]), .B(_14488_), .Y(_03537_));
NOR_g _24311_ (.A(_03536_), .B(_03537_), .Y(_01021_));
NAND_g _24312_ (.A(reg_pc[4]), .B(_14617_), .Y(_03538_));
NAND_g _24313_ (.A(cpuregs[7][4]), .B(_00008_[2]), .Y(_03539_));
NAND_g _24314_ (.A(cpuregs[3][4]), .B(_09032_), .Y(_03540_));
NAND_g _24315_ (.A(_03539_), .B(_03540_), .Y(_03541_));
AND_g _24316_ (.A(_00008_[0]), .B(_03541_), .Y(_03542_));
NAND_g _24317_ (.A(cpuregs[6][4]), .B(_00008_[2]), .Y(_03543_));
NAND_g _24318_ (.A(cpuregs[2][4]), .B(_09032_), .Y(_03544_));
AND_g _24319_ (.A(_03543_), .B(_03544_), .Y(_03545_));
NOR_g _24320_ (.A(_00008_[0]), .B(_03545_), .Y(_03546_));
NOR_g _24321_ (.A(_03542_), .B(_03546_), .Y(_03547_));
NAND_g _24322_ (.A(cpuregs[5][4]), .B(_00008_[2]), .Y(_03548_));
NAND_g _24323_ (.A(cpuregs[1][4]), .B(_09032_), .Y(_03549_));
NAND_g _24324_ (.A(_03548_), .B(_03549_), .Y(_03550_));
NAND_g _24325_ (.A(_00008_[0]), .B(_03550_), .Y(_03551_));
NAND_g _24326_ (.A(cpuregs[4][4]), .B(_00008_[2]), .Y(_03552_));
NAND_g _24327_ (.A(cpuregs[0][4]), .B(_09032_), .Y(_03553_));
AND_g _24328_ (.A(_03552_), .B(_03553_), .Y(_03554_));
NOR_g _24329_ (.A(_00008_[0]), .B(_03554_), .Y(_03555_));
NAND_g _24330_ (.A(_00008_[1]), .B(_03547_), .Y(_03556_));
NOR_g _24331_ (.A(_00008_[1]), .B(_03555_), .Y(_03557_));
NAND_g _24332_ (.A(_03551_), .B(_03557_), .Y(_03558_));
AND_g _24333_ (.A(_03556_), .B(_03558_), .Y(_03559_));
NAND_g _24334_ (.A(_09033_), .B(_03559_), .Y(_03560_));
NAND_g _24335_ (.A(cpuregs[13][4]), .B(_00008_[0]), .Y(_03561_));
NAND_g _24336_ (.A(cpuregs[12][4]), .B(_09030_), .Y(_03562_));
AND_g _24337_ (.A(_00008_[2]), .B(_03562_), .Y(_03563_));
NAND_g _24338_ (.A(_03561_), .B(_03563_), .Y(_03564_));
NAND_g _24339_ (.A(cpuregs[9][4]), .B(_00008_[0]), .Y(_03565_));
NAND_g _24340_ (.A(cpuregs[8][4]), .B(_09030_), .Y(_03566_));
AND_g _24341_ (.A(_09032_), .B(_03566_), .Y(_03567_));
NAND_g _24342_ (.A(_03565_), .B(_03567_), .Y(_03568_));
AND_g _24343_ (.A(_09031_), .B(_03568_), .Y(_03569_));
NAND_g _24344_ (.A(_03564_), .B(_03569_), .Y(_03570_));
NAND_g _24345_ (.A(cpuregs[15][4]), .B(_00008_[0]), .Y(_03571_));
NAND_g _24346_ (.A(cpuregs[14][4]), .B(_09030_), .Y(_03572_));
AND_g _24347_ (.A(_00008_[2]), .B(_03572_), .Y(_03573_));
NAND_g _24348_ (.A(_03571_), .B(_03573_), .Y(_03574_));
NAND_g _24349_ (.A(cpuregs[11][4]), .B(_00008_[0]), .Y(_03575_));
NAND_g _24350_ (.A(cpuregs[10][4]), .B(_09030_), .Y(_03576_));
AND_g _24351_ (.A(_09032_), .B(_03576_), .Y(_03577_));
NAND_g _24352_ (.A(_03575_), .B(_03577_), .Y(_03578_));
AND_g _24353_ (.A(_00008_[1]), .B(_03578_), .Y(_03579_));
NAND_g _24354_ (.A(_03574_), .B(_03579_), .Y(_03580_));
NAND_g _24355_ (.A(_03570_), .B(_03580_), .Y(_03581_));
AND_g _24356_ (.A(_00008_[3]), .B(_03581_), .Y(_03582_));
NOR_g _24357_ (.A(_00008_[4]), .B(_03582_), .Y(_03583_));
NAND_g _24358_ (.A(_03560_), .B(_03583_), .Y(_03584_));
NAND_g _24359_ (.A(cpuregs[25][4]), .B(_09032_), .Y(_03585_));
NAND_g _24360_ (.A(cpuregs[29][4]), .B(_00008_[2]), .Y(_03586_));
AND_g _24361_ (.A(_09031_), .B(_03586_), .Y(_03587_));
NAND_g _24362_ (.A(_03585_), .B(_03587_), .Y(_03588_));
NAND_g _24363_ (.A(cpuregs[31][4]), .B(_00008_[2]), .Y(_03589_));
NAND_g _24364_ (.A(cpuregs[27][4]), .B(_09032_), .Y(_03590_));
AND_g _24365_ (.A(_00008_[1]), .B(_03590_), .Y(_03591_));
NAND_g _24366_ (.A(_03589_), .B(_03591_), .Y(_03592_));
NAND_g _24367_ (.A(_03588_), .B(_03592_), .Y(_03593_));
NAND_g _24368_ (.A(_00008_[0]), .B(_03593_), .Y(_03594_));
NAND_g _24369_ (.A(cpuregs[24][4]), .B(_09032_), .Y(_03595_));
NAND_g _24370_ (.A(cpuregs[28][4]), .B(_00008_[2]), .Y(_03596_));
AND_g _24371_ (.A(_09031_), .B(_03596_), .Y(_03597_));
NAND_g _24372_ (.A(_03595_), .B(_03597_), .Y(_03598_));
NAND_g _24373_ (.A(cpuregs[26][4]), .B(_09032_), .Y(_03599_));
NAND_g _24374_ (.A(cpuregs[30][4]), .B(_00008_[2]), .Y(_03600_));
AND_g _24375_ (.A(_00008_[1]), .B(_03600_), .Y(_03601_));
NAND_g _24376_ (.A(_03599_), .B(_03601_), .Y(_03602_));
NAND_g _24377_ (.A(_03598_), .B(_03602_), .Y(_03603_));
NAND_g _24378_ (.A(_09030_), .B(_03603_), .Y(_03604_));
NAND_g _24379_ (.A(_03594_), .B(_03604_), .Y(_03605_));
NAND_g _24380_ (.A(_00008_[3]), .B(_03605_), .Y(_03606_));
NAND_g _24381_ (.A(cpuregs[17][4]), .B(_09031_), .Y(_03607_));
NAND_g _24382_ (.A(cpuregs[19][4]), .B(_00008_[1]), .Y(_03608_));
AND_g _24383_ (.A(_09032_), .B(_03608_), .Y(_03609_));
NAND_g _24384_ (.A(_03607_), .B(_03609_), .Y(_03610_));
NAND_g _24385_ (.A(cpuregs[21][4]), .B(_09031_), .Y(_03611_));
NAND_g _24386_ (.A(cpuregs[23][4]), .B(_00008_[1]), .Y(_03612_));
AND_g _24387_ (.A(_00008_[2]), .B(_03612_), .Y(_03613_));
NAND_g _24388_ (.A(_03611_), .B(_03613_), .Y(_03614_));
NAND_g _24389_ (.A(_03610_), .B(_03614_), .Y(_03615_));
NAND_g _24390_ (.A(_00008_[0]), .B(_03615_), .Y(_03616_));
NAND_g _24391_ (.A(cpuregs[16][4]), .B(_09031_), .Y(_03617_));
NAND_g _24392_ (.A(cpuregs[18][4]), .B(_00008_[1]), .Y(_03618_));
AND_g _24393_ (.A(_09032_), .B(_03618_), .Y(_03619_));
NAND_g _24394_ (.A(_03617_), .B(_03619_), .Y(_03620_));
NAND_g _24395_ (.A(cpuregs[20][4]), .B(_09031_), .Y(_03621_));
NAND_g _24396_ (.A(cpuregs[22][4]), .B(_00008_[1]), .Y(_03622_));
AND_g _24397_ (.A(_00008_[2]), .B(_03622_), .Y(_03623_));
NAND_g _24398_ (.A(_03621_), .B(_03623_), .Y(_03624_));
NAND_g _24399_ (.A(_03620_), .B(_03624_), .Y(_03625_));
NAND_g _24400_ (.A(_09030_), .B(_03625_), .Y(_03626_));
NAND_g _24401_ (.A(_03616_), .B(_03626_), .Y(_03627_));
AND_g _24402_ (.A(_09033_), .B(_03627_), .Y(_03628_));
NOT_g _24403_ (.A(_03628_), .Y(_03629_));
NAND_g _24404_ (.A(_03606_), .B(_03629_), .Y(_03630_));
NAND_g _24405_ (.A(_00008_[4]), .B(_03630_), .Y(_03631_));
AND_g _24406_ (.A(_14624_), .B(_03631_), .Y(_03632_));
NAND_g _24407_ (.A(_03584_), .B(_03632_), .Y(_03633_));
NAND_g _24408_ (.A(_03538_), .B(_03633_), .Y(_03634_));
NAND_g _24409_ (.A(_10595_), .B(_03634_), .Y(_03635_));
XOR_g _24410_ (.A(_14543_), .B(_14557_), .Y(_03636_));
NAND_g _24411_ (.A(_14614_), .B(_03636_), .Y(_03637_));
NAND_g _24412_ (.A(pcpi_rs1[3]), .B(_14481_), .Y(_03638_));
AND_g _24413_ (.A(_03304_), .B(_03638_), .Y(_03639_));
NAND_g _24414_ (.A(_13879_), .B(_03639_), .Y(_03640_));
NAND_g _24415_ (.A(pcpi_rs1[8]), .B(_14482_), .Y(_03641_));
AND_g _24416_ (.A(_03303_), .B(_03641_), .Y(_03642_));
NAND_g _24417_ (.A(_13880_), .B(_03642_), .Y(_03643_));
AND_g _24418_ (.A(_03640_), .B(_03643_), .Y(_03644_));
NAND_g _24419_ (.A(_13883_), .B(_03644_), .Y(_03645_));
AND_g _24420_ (.A(_03637_), .B(_03645_), .Y(_03646_));
AND_g _24421_ (.A(_14488_), .B(_03646_), .Y(_03647_));
AND_g _24422_ (.A(_03635_), .B(_03647_), .Y(_03648_));
NOR_g _24423_ (.A(pcpi_rs1[4]), .B(_14488_), .Y(_03649_));
NOR_g _24424_ (.A(_03648_), .B(_03649_), .Y(_01022_));
NOR_g _24425_ (.A(pcpi_rs1[5]), .B(_14488_), .Y(_03650_));
AND_g _24426_ (.A(reg_pc[5]), .B(_14617_), .Y(_03651_));
NAND_g _24427_ (.A(cpuregs[26][5]), .B(_09032_), .Y(_03652_));
NAND_g _24428_ (.A(cpuregs[30][5]), .B(_00008_[2]), .Y(_03653_));
AND_g _24429_ (.A(_09030_), .B(_03653_), .Y(_03654_));
NAND_g _24430_ (.A(_03652_), .B(_03654_), .Y(_03655_));
NAND_g _24431_ (.A(cpuregs[31][5]), .B(_00008_[2]), .Y(_03656_));
NAND_g _24432_ (.A(cpuregs[27][5]), .B(_09032_), .Y(_03657_));
AND_g _24433_ (.A(_00008_[0]), .B(_03657_), .Y(_03658_));
NAND_g _24434_ (.A(_03656_), .B(_03658_), .Y(_03659_));
NAND_g _24435_ (.A(_03655_), .B(_03659_), .Y(_03660_));
NAND_g _24436_ (.A(_00008_[3]), .B(_03660_), .Y(_03661_));
NAND_g _24437_ (.A(cpuregs[18][5]), .B(_09032_), .Y(_03662_));
NAND_g _24438_ (.A(cpuregs[22][5]), .B(_00008_[2]), .Y(_03663_));
AND_g _24439_ (.A(_09030_), .B(_03663_), .Y(_03664_));
NAND_g _24440_ (.A(_03662_), .B(_03664_), .Y(_03665_));
NAND_g _24441_ (.A(cpuregs[19][5]), .B(_09032_), .Y(_03666_));
NAND_g _24442_ (.A(cpuregs[23][5]), .B(_00008_[2]), .Y(_03667_));
AND_g _24443_ (.A(_00008_[0]), .B(_03667_), .Y(_03668_));
NAND_g _24444_ (.A(_03666_), .B(_03668_), .Y(_03669_));
NAND_g _24445_ (.A(_03665_), .B(_03669_), .Y(_03670_));
NAND_g _24446_ (.A(_09033_), .B(_03670_), .Y(_03671_));
NAND_g _24447_ (.A(cpuregs[16][5]), .B(_09032_), .Y(_03672_));
NAND_g _24448_ (.A(cpuregs[20][5]), .B(_00008_[2]), .Y(_03673_));
AND_g _24449_ (.A(_09030_), .B(_03673_), .Y(_03674_));
NAND_g _24450_ (.A(_03672_), .B(_03674_), .Y(_03675_));
NAND_g _24451_ (.A(cpuregs[17][5]), .B(_09032_), .Y(_03676_));
NAND_g _24452_ (.A(cpuregs[21][5]), .B(_00008_[2]), .Y(_03677_));
AND_g _24453_ (.A(_00008_[0]), .B(_03677_), .Y(_03678_));
NAND_g _24454_ (.A(_03676_), .B(_03678_), .Y(_03679_));
NAND_g _24455_ (.A(_03675_), .B(_03679_), .Y(_03680_));
NAND_g _24456_ (.A(_09033_), .B(_03680_), .Y(_03681_));
NAND_g _24457_ (.A(cpuregs[24][5]), .B(_09032_), .Y(_03682_));
NAND_g _24458_ (.A(cpuregs[28][5]), .B(_00008_[2]), .Y(_03683_));
AND_g _24459_ (.A(_09030_), .B(_03683_), .Y(_03684_));
NAND_g _24460_ (.A(_03682_), .B(_03684_), .Y(_03685_));
NAND_g _24461_ (.A(cpuregs[25][5]), .B(_09032_), .Y(_03686_));
NAND_g _24462_ (.A(cpuregs[29][5]), .B(_00008_[2]), .Y(_03687_));
AND_g _24463_ (.A(_00008_[0]), .B(_03687_), .Y(_03688_));
NAND_g _24464_ (.A(_03686_), .B(_03688_), .Y(_03689_));
NAND_g _24465_ (.A(_03685_), .B(_03689_), .Y(_03690_));
NAND_g _24466_ (.A(_00008_[3]), .B(_03690_), .Y(_03691_));
AND_g _24467_ (.A(_00008_[1]), .B(_03671_), .Y(_03692_));
NAND_g _24468_ (.A(_03661_), .B(_03692_), .Y(_03693_));
AND_g _24469_ (.A(_09031_), .B(_03691_), .Y(_03694_));
NAND_g _24470_ (.A(_03681_), .B(_03694_), .Y(_03695_));
AND_g _24471_ (.A(_00008_[4]), .B(_03695_), .Y(_03696_));
NAND_g _24472_ (.A(_03693_), .B(_03696_), .Y(_03697_));
NAND_g _24473_ (.A(cpuregs[9][5]), .B(_09032_), .Y(_03698_));
NAND_g _24474_ (.A(cpuregs[13][5]), .B(_00008_[2]), .Y(_03699_));
AND_g _24475_ (.A(_09031_), .B(_03699_), .Y(_03700_));
NAND_g _24476_ (.A(_03698_), .B(_03700_), .Y(_03701_));
NAND_g _24477_ (.A(cpuregs[15][5]), .B(_00008_[2]), .Y(_03702_));
NAND_g _24478_ (.A(cpuregs[11][5]), .B(_09032_), .Y(_03703_));
AND_g _24479_ (.A(_00008_[1]), .B(_03703_), .Y(_03704_));
NAND_g _24480_ (.A(_03702_), .B(_03704_), .Y(_03705_));
NAND_g _24481_ (.A(_03701_), .B(_03705_), .Y(_03706_));
NAND_g _24482_ (.A(_00008_[0]), .B(_03706_), .Y(_03707_));
NAND_g _24483_ (.A(cpuregs[8][5]), .B(_09032_), .Y(_03708_));
NAND_g _24484_ (.A(cpuregs[12][5]), .B(_00008_[2]), .Y(_03709_));
AND_g _24485_ (.A(_09031_), .B(_03709_), .Y(_03710_));
NAND_g _24486_ (.A(_03708_), .B(_03710_), .Y(_03711_));
NAND_g _24487_ (.A(cpuregs[10][5]), .B(_09032_), .Y(_03712_));
NAND_g _24488_ (.A(cpuregs[14][5]), .B(_00008_[2]), .Y(_03713_));
AND_g _24489_ (.A(_00008_[1]), .B(_03713_), .Y(_03714_));
NAND_g _24490_ (.A(_03712_), .B(_03714_), .Y(_03715_));
NAND_g _24491_ (.A(_03711_), .B(_03715_), .Y(_03716_));
NAND_g _24492_ (.A(_09030_), .B(_03716_), .Y(_03717_));
NAND_g _24493_ (.A(_03707_), .B(_03717_), .Y(_03718_));
NAND_g _24494_ (.A(_00008_[3]), .B(_03718_), .Y(_03719_));
NAND_g _24495_ (.A(cpuregs[1][5]), .B(_09031_), .Y(_03720_));
NAND_g _24496_ (.A(cpuregs[3][5]), .B(_00008_[1]), .Y(_03721_));
AND_g _24497_ (.A(_09032_), .B(_03721_), .Y(_03722_));
NAND_g _24498_ (.A(_03720_), .B(_03722_), .Y(_03723_));
NAND_g _24499_ (.A(cpuregs[5][5]), .B(_09031_), .Y(_03724_));
NAND_g _24500_ (.A(cpuregs[7][5]), .B(_00008_[1]), .Y(_03725_));
AND_g _24501_ (.A(_00008_[2]), .B(_03725_), .Y(_03726_));
NAND_g _24502_ (.A(_03724_), .B(_03726_), .Y(_03727_));
NAND_g _24503_ (.A(_03723_), .B(_03727_), .Y(_03728_));
NAND_g _24504_ (.A(_00008_[0]), .B(_03728_), .Y(_03729_));
NAND_g _24505_ (.A(cpuregs[0][5]), .B(_09031_), .Y(_03730_));
NAND_g _24506_ (.A(cpuregs[2][5]), .B(_00008_[1]), .Y(_03731_));
AND_g _24507_ (.A(_09032_), .B(_03731_), .Y(_03732_));
NAND_g _24508_ (.A(_03730_), .B(_03732_), .Y(_03733_));
NAND_g _24509_ (.A(cpuregs[4][5]), .B(_09031_), .Y(_03734_));
NAND_g _24510_ (.A(cpuregs[6][5]), .B(_00008_[1]), .Y(_03735_));
AND_g _24511_ (.A(_00008_[2]), .B(_03735_), .Y(_03736_));
NAND_g _24512_ (.A(_03734_), .B(_03736_), .Y(_03737_));
NAND_g _24513_ (.A(_03733_), .B(_03737_), .Y(_03738_));
NAND_g _24514_ (.A(_09030_), .B(_03738_), .Y(_03739_));
NAND_g _24515_ (.A(_03729_), .B(_03739_), .Y(_03740_));
NAND_g _24516_ (.A(_09033_), .B(_03740_), .Y(_03741_));
AND_g _24517_ (.A(_03719_), .B(_03741_), .Y(_03742_));
NOR_g _24518_ (.A(_00008_[4]), .B(_03742_), .Y(_03743_));
NAND_g _24519_ (.A(_14624_), .B(_03697_), .Y(_03744_));
NOR_g _24520_ (.A(_03743_), .B(_03744_), .Y(_03745_));
NOR_g _24521_ (.A(_03651_), .B(_03745_), .Y(_03746_));
NOR_g _24522_ (.A(_10596_), .B(_03746_), .Y(_03747_));
XOR_g _24523_ (.A(_14559_), .B(_14560_), .Y(_03748_));
NAND_g _24524_ (.A(_14614_), .B(_03748_), .Y(_03749_));
NAND_g _24525_ (.A(pcpi_rs1[4]), .B(_14481_), .Y(_03750_));
AND_g _24526_ (.A(_13879_), .B(_03750_), .Y(_03751_));
NAND_g _24527_ (.A(_03415_), .B(_03751_), .Y(_03752_));
NAND_g _24528_ (.A(pcpi_rs1[9]), .B(_14482_), .Y(_03753_));
AND_g _24529_ (.A(_03414_), .B(_03753_), .Y(_03754_));
NAND_g _24530_ (.A(_13880_), .B(_03754_), .Y(_03755_));
AND_g _24531_ (.A(_03752_), .B(_03755_), .Y(_03756_));
NAND_g _24532_ (.A(_13883_), .B(_03756_), .Y(_03757_));
AND_g _24533_ (.A(_14488_), .B(_03757_), .Y(_03758_));
NAND_g _24534_ (.A(_03749_), .B(_03758_), .Y(_03759_));
NOR_g _24535_ (.A(_03747_), .B(_03759_), .Y(_03760_));
NOR_g _24536_ (.A(_03650_), .B(_03760_), .Y(_01023_));
NOR_g _24537_ (.A(pcpi_rs1[6]), .B(_14488_), .Y(_03761_));
NAND_g _24538_ (.A(reg_pc[6]), .B(_14617_), .Y(_03762_));
NAND_g _24539_ (.A(cpuregs[7][6]), .B(_00008_[2]), .Y(_03763_));
NAND_g _24540_ (.A(cpuregs[3][6]), .B(_09032_), .Y(_03764_));
NAND_g _24541_ (.A(_03763_), .B(_03764_), .Y(_03765_));
NAND_g _24542_ (.A(_00008_[0]), .B(_03765_), .Y(_03766_));
NAND_g _24543_ (.A(cpuregs[6][6]), .B(_00008_[2]), .Y(_03767_));
NAND_g _24544_ (.A(cpuregs[2][6]), .B(_09032_), .Y(_03768_));
NAND_g _24545_ (.A(_03767_), .B(_03768_), .Y(_03769_));
NAND_g _24546_ (.A(_09030_), .B(_03769_), .Y(_03770_));
AND_g _24547_ (.A(_03766_), .B(_03770_), .Y(_03771_));
NAND_g _24548_ (.A(_08905_), .B(_00008_[2]), .Y(_03772_));
NOR_g _24549_ (.A(cpuregs[0][6]), .B(_00008_[2]), .Y(_03773_));
NOR_g _24550_ (.A(_00008_[0]), .B(_03773_), .Y(_03774_));
NAND_g _24551_ (.A(_03772_), .B(_03774_), .Y(_03775_));
NAND_g _24552_ (.A(_08947_), .B(_00008_[2]), .Y(_03776_));
NOR_g _24553_ (.A(cpuregs[1][6]), .B(_00008_[2]), .Y(_03777_));
NOR_g _24554_ (.A(_09030_), .B(_03777_), .Y(_03778_));
NAND_g _24555_ (.A(_03776_), .B(_03778_), .Y(_03779_));
AND_g _24556_ (.A(_03775_), .B(_03779_), .Y(_03780_));
NAND_g _24557_ (.A(cpuregs[11][6]), .B(_09032_), .Y(_03781_));
NAND_g _24558_ (.A(cpuregs[15][6]), .B(_00008_[2]), .Y(_03782_));
NAND_g _24559_ (.A(_03781_), .B(_03782_), .Y(_03783_));
AND_g _24560_ (.A(_00008_[0]), .B(_03783_), .Y(_03784_));
NAND_g _24561_ (.A(cpuregs[14][6]), .B(_00008_[2]), .Y(_03785_));
NAND_g _24562_ (.A(cpuregs[10][6]), .B(_09032_), .Y(_03786_));
AND_g _24563_ (.A(_03785_), .B(_03786_), .Y(_03787_));
NOR_g _24564_ (.A(_00008_[0]), .B(_03787_), .Y(_03788_));
NOR_g _24565_ (.A(_03784_), .B(_03788_), .Y(_03789_));
NAND_g _24566_ (.A(_08880_), .B(_00008_[2]), .Y(_03790_));
NOR_g _24567_ (.A(cpuregs[8][6]), .B(_00008_[2]), .Y(_03791_));
NOR_g _24568_ (.A(_00008_[0]), .B(_03791_), .Y(_03792_));
AND_g _24569_ (.A(_03790_), .B(_03792_), .Y(_03793_));
NOR_g _24570_ (.A(cpuregs[9][6]), .B(_00008_[2]), .Y(_03794_));
NAND_g _24571_ (.A(_08928_), .B(_00008_[2]), .Y(_03795_));
NAND_g _24572_ (.A(_00008_[0]), .B(_03795_), .Y(_03796_));
NOR_g _24573_ (.A(_03794_), .B(_03796_), .Y(_03797_));
NOR_g _24574_ (.A(_03793_), .B(_03797_), .Y(_03798_));
AND_g _24575_ (.A(_09033_), .B(_03780_), .Y(_03799_));
NOT_g _24576_ (.A(_03799_), .Y(_03800_));
NAND_g _24577_ (.A(_00008_[3]), .B(_03798_), .Y(_03801_));
AND_g _24578_ (.A(_09031_), .B(_03801_), .Y(_03802_));
NAND_g _24579_ (.A(_03800_), .B(_03802_), .Y(_03803_));
NAND_g _24580_ (.A(_00008_[3]), .B(_03789_), .Y(_03804_));
NAND_g _24581_ (.A(_09033_), .B(_03771_), .Y(_03805_));
AND_g _24582_ (.A(_03804_), .B(_03805_), .Y(_03806_));
AND_g _24583_ (.A(_00008_[1]), .B(_03806_), .Y(_03807_));
NOR_g _24584_ (.A(_00008_[4]), .B(_03807_), .Y(_03808_));
NAND_g _24585_ (.A(_03803_), .B(_03808_), .Y(_03809_));
NAND_g _24586_ (.A(_08886_), .B(_00008_[2]), .Y(_03810_));
NOR_g _24587_ (.A(cpuregs[19][6]), .B(_00008_[2]), .Y(_03811_));
NOR_g _24588_ (.A(cpuregs[18][6]), .B(_00008_[2]), .Y(_03812_));
AND_g _24589_ (.A(_08918_), .B(_00008_[2]), .Y(_03813_));
NOR_g _24590_ (.A(_03812_), .B(_03813_), .Y(_03814_));
NOR_g _24591_ (.A(_09030_), .B(_03811_), .Y(_03815_));
NAND_g _24592_ (.A(_03810_), .B(_03815_), .Y(_03816_));
NAND_g _24593_ (.A(_09030_), .B(_03814_), .Y(_03817_));
AND_g _24594_ (.A(_03816_), .B(_03817_), .Y(_03818_));
NAND_g _24595_ (.A(_00008_[1]), .B(_03818_), .Y(_03819_));
NOR_g _24596_ (.A(cpuregs[17][6]), .B(_00008_[2]), .Y(_03820_));
NAND_g _24597_ (.A(_08985_), .B(_00008_[2]), .Y(_03821_));
NOR_g _24598_ (.A(cpuregs[16][6]), .B(_00008_[2]), .Y(_03822_));
AND_g _24599_ (.A(_08844_), .B(_00008_[2]), .Y(_03823_));
NOR_g _24600_ (.A(_03822_), .B(_03823_), .Y(_03824_));
NOR_g _24601_ (.A(_09030_), .B(_03820_), .Y(_03825_));
NAND_g _24602_ (.A(_03821_), .B(_03825_), .Y(_03826_));
NAND_g _24603_ (.A(_09030_), .B(_03824_), .Y(_03827_));
AND_g _24604_ (.A(_03826_), .B(_03827_), .Y(_03828_));
NAND_g _24605_ (.A(_09031_), .B(_03828_), .Y(_03829_));
NAND_g _24606_ (.A(_03819_), .B(_03829_), .Y(_03830_));
NAND_g _24607_ (.A(_09033_), .B(_03830_), .Y(_03831_));
NAND_g _24608_ (.A(cpuregs[25][6]), .B(_09031_), .Y(_03832_));
NAND_g _24609_ (.A(cpuregs[27][6]), .B(_00008_[1]), .Y(_03833_));
AND_g _24610_ (.A(_09032_), .B(_03833_), .Y(_03834_));
NAND_g _24611_ (.A(_03832_), .B(_03834_), .Y(_03835_));
NAND_g _24612_ (.A(cpuregs[29][6]), .B(_09031_), .Y(_03836_));
NAND_g _24613_ (.A(cpuregs[31][6]), .B(_00008_[1]), .Y(_03837_));
AND_g _24614_ (.A(_00008_[2]), .B(_03837_), .Y(_03838_));
NAND_g _24615_ (.A(_03836_), .B(_03838_), .Y(_03839_));
NAND_g _24616_ (.A(_03835_), .B(_03839_), .Y(_03840_));
NAND_g _24617_ (.A(_00008_[0]), .B(_03840_), .Y(_03841_));
NAND_g _24618_ (.A(cpuregs[24][6]), .B(_09031_), .Y(_03842_));
NAND_g _24619_ (.A(cpuregs[26][6]), .B(_00008_[1]), .Y(_03843_));
AND_g _24620_ (.A(_09032_), .B(_03843_), .Y(_03844_));
NAND_g _24621_ (.A(_03842_), .B(_03844_), .Y(_03845_));
NAND_g _24622_ (.A(cpuregs[28][6]), .B(_09031_), .Y(_03846_));
NAND_g _24623_ (.A(cpuregs[30][6]), .B(_00008_[1]), .Y(_03847_));
AND_g _24624_ (.A(_00008_[2]), .B(_03847_), .Y(_03848_));
NAND_g _24625_ (.A(_03846_), .B(_03848_), .Y(_03849_));
NAND_g _24626_ (.A(_03845_), .B(_03849_), .Y(_03850_));
NAND_g _24627_ (.A(_09030_), .B(_03850_), .Y(_03851_));
NAND_g _24628_ (.A(_03841_), .B(_03851_), .Y(_03852_));
NAND_g _24629_ (.A(_00008_[3]), .B(_03852_), .Y(_03853_));
NAND_g _24630_ (.A(_03831_), .B(_03853_), .Y(_03854_));
NAND_g _24631_ (.A(_00008_[4]), .B(_03854_), .Y(_03855_));
AND_g _24632_ (.A(_14624_), .B(_03809_), .Y(_03856_));
NAND_g _24633_ (.A(_03855_), .B(_03856_), .Y(_03857_));
NAND_g _24634_ (.A(_03762_), .B(_03857_), .Y(_03858_));
NAND_g _24635_ (.A(_10595_), .B(_03858_), .Y(_03859_));
NAND_g _24636_ (.A(pcpi_rs1[5]), .B(_14481_), .Y(_03860_));
AND_g _24637_ (.A(_03526_), .B(_03860_), .Y(_03861_));
NAND_g _24638_ (.A(pcpi_rs1[10]), .B(_14482_), .Y(_03862_));
AND_g _24639_ (.A(_03529_), .B(_03862_), .Y(_03863_));
NAND_g _24640_ (.A(_13880_), .B(_03863_), .Y(_03864_));
NAND_g _24641_ (.A(_13879_), .B(_03861_), .Y(_03865_));
AND_g _24642_ (.A(_13883_), .B(_03864_), .Y(_03866_));
NAND_g _24643_ (.A(_03865_), .B(_03866_), .Y(_03867_));
AND_g _24644_ (.A(_14488_), .B(_03867_), .Y(_03868_));
AND_g _24645_ (.A(_03859_), .B(_03868_), .Y(_03869_));
XOR_g _24646_ (.A(_14540_), .B(_14562_), .Y(_03870_));
NAND_g _24647_ (.A(_14614_), .B(_03870_), .Y(_03871_));
AND_g _24648_ (.A(_03869_), .B(_03871_), .Y(_03872_));
NOR_g _24649_ (.A(_03761_), .B(_03872_), .Y(_01024_));
XOR_g _24650_ (.A(decoded_imm[7]), .B(pcpi_rs1[7]), .Y(_03873_));
XNOR_g _24651_ (.A(_14564_), .B(_03873_), .Y(_03874_));
NAND_g _24652_ (.A(_14614_), .B(_03874_), .Y(_03875_));
NAND_g _24653_ (.A(reg_pc[7]), .B(_14617_), .Y(_03876_));
NAND_g _24654_ (.A(cpuregs[27][7]), .B(_00008_[0]), .Y(_03877_));
NAND_g _24655_ (.A(cpuregs[26][7]), .B(_09030_), .Y(_03878_));
AND_g _24656_ (.A(_09032_), .B(_03878_), .Y(_03879_));
NAND_g _24657_ (.A(_03877_), .B(_03879_), .Y(_03880_));
NAND_g _24658_ (.A(cpuregs[31][7]), .B(_00008_[0]), .Y(_03881_));
NAND_g _24659_ (.A(cpuregs[30][7]), .B(_09030_), .Y(_03882_));
AND_g _24660_ (.A(_00008_[2]), .B(_03882_), .Y(_03883_));
NAND_g _24661_ (.A(_03881_), .B(_03883_), .Y(_03884_));
NAND_g _24662_ (.A(_03880_), .B(_03884_), .Y(_03885_));
NAND_g _24663_ (.A(_00008_[1]), .B(_03885_), .Y(_03886_));
NAND_g _24664_ (.A(cpuregs[25][7]), .B(_00008_[0]), .Y(_03887_));
NAND_g _24665_ (.A(cpuregs[24][7]), .B(_09030_), .Y(_03888_));
AND_g _24666_ (.A(_09032_), .B(_03888_), .Y(_03889_));
NAND_g _24667_ (.A(_03887_), .B(_03889_), .Y(_03890_));
NAND_g _24668_ (.A(cpuregs[29][7]), .B(_00008_[0]), .Y(_03891_));
NAND_g _24669_ (.A(cpuregs[28][7]), .B(_09030_), .Y(_03892_));
AND_g _24670_ (.A(_00008_[2]), .B(_03892_), .Y(_03893_));
NAND_g _24671_ (.A(_03891_), .B(_03893_), .Y(_03894_));
NAND_g _24672_ (.A(_03890_), .B(_03894_), .Y(_03895_));
NAND_g _24673_ (.A(_09031_), .B(_03895_), .Y(_03896_));
NAND_g _24674_ (.A(_03886_), .B(_03896_), .Y(_03897_));
NAND_g _24675_ (.A(_00008_[3]), .B(_03897_), .Y(_03898_));
NAND_g _24676_ (.A(cpuregs[22][7]), .B(_00008_[2]), .Y(_03899_));
NAND_g _24677_ (.A(cpuregs[18][7]), .B(_09032_), .Y(_03900_));
AND_g _24678_ (.A(_03899_), .B(_03900_), .Y(_03901_));
NOR_g _24679_ (.A(_00008_[0]), .B(_03901_), .Y(_03902_));
NAND_g _24680_ (.A(cpuregs[23][7]), .B(_00008_[2]), .Y(_03903_));
NAND_g _24681_ (.A(cpuregs[19][7]), .B(_09032_), .Y(_03904_));
NAND_g _24682_ (.A(_03903_), .B(_03904_), .Y(_03905_));
AND_g _24683_ (.A(_00008_[0]), .B(_03905_), .Y(_03906_));
NOR_g _24684_ (.A(_03902_), .B(_03906_), .Y(_03907_));
NAND_g _24685_ (.A(_00008_[1]), .B(_03907_), .Y(_03908_));
NAND_g _24686_ (.A(cpuregs[20][7]), .B(_00008_[2]), .Y(_03909_));
NAND_g _24687_ (.A(cpuregs[16][7]), .B(_09032_), .Y(_03910_));
NAND_g _24688_ (.A(_03909_), .B(_03910_), .Y(_03911_));
NAND_g _24689_ (.A(_09030_), .B(_03911_), .Y(_03912_));
NAND_g _24690_ (.A(cpuregs[21][7]), .B(_00008_[2]), .Y(_03913_));
NAND_g _24691_ (.A(cpuregs[17][7]), .B(_09032_), .Y(_03914_));
NAND_g _24692_ (.A(_03913_), .B(_03914_), .Y(_03915_));
NAND_g _24693_ (.A(_00008_[0]), .B(_03915_), .Y(_03916_));
AND_g _24694_ (.A(_03912_), .B(_03916_), .Y(_03917_));
NAND_g _24695_ (.A(_09031_), .B(_03917_), .Y(_03918_));
NAND_g _24696_ (.A(_03908_), .B(_03918_), .Y(_03919_));
NAND_g _24697_ (.A(_09033_), .B(_03919_), .Y(_03920_));
AND_g _24698_ (.A(_00008_[4]), .B(_03920_), .Y(_03921_));
NAND_g _24699_ (.A(_03898_), .B(_03921_), .Y(_03922_));
NAND_g _24700_ (.A(cpuregs[1][7]), .B(_09031_), .Y(_03923_));
NAND_g _24701_ (.A(cpuregs[3][7]), .B(_00008_[1]), .Y(_03924_));
AND_g _24702_ (.A(_09032_), .B(_03924_), .Y(_03925_));
NAND_g _24703_ (.A(_03923_), .B(_03925_), .Y(_03926_));
NAND_g _24704_ (.A(cpuregs[5][7]), .B(_09031_), .Y(_03927_));
NAND_g _24705_ (.A(cpuregs[7][7]), .B(_00008_[1]), .Y(_03928_));
AND_g _24706_ (.A(_00008_[2]), .B(_03928_), .Y(_03929_));
NAND_g _24707_ (.A(_03927_), .B(_03929_), .Y(_03930_));
NAND_g _24708_ (.A(_03926_), .B(_03930_), .Y(_03931_));
NAND_g _24709_ (.A(_00008_[0]), .B(_03931_), .Y(_03932_));
NAND_g _24710_ (.A(cpuregs[0][7]), .B(_09031_), .Y(_03933_));
NAND_g _24711_ (.A(cpuregs[2][7]), .B(_00008_[1]), .Y(_03934_));
AND_g _24712_ (.A(_09032_), .B(_03934_), .Y(_03935_));
NAND_g _24713_ (.A(_03933_), .B(_03935_), .Y(_03936_));
NAND_g _24714_ (.A(cpuregs[4][7]), .B(_09031_), .Y(_03937_));
NAND_g _24715_ (.A(cpuregs[6][7]), .B(_00008_[1]), .Y(_03938_));
AND_g _24716_ (.A(_00008_[2]), .B(_03938_), .Y(_03939_));
NAND_g _24717_ (.A(_03937_), .B(_03939_), .Y(_03940_));
NAND_g _24718_ (.A(_03936_), .B(_03940_), .Y(_03941_));
NAND_g _24719_ (.A(_09030_), .B(_03941_), .Y(_03942_));
NAND_g _24720_ (.A(_03932_), .B(_03942_), .Y(_03943_));
NAND_g _24721_ (.A(_09033_), .B(_03943_), .Y(_03944_));
NAND_g _24722_ (.A(cpuregs[9][7]), .B(_09032_), .Y(_03945_));
NAND_g _24723_ (.A(cpuregs[13][7]), .B(_00008_[2]), .Y(_03946_));
AND_g _24724_ (.A(_09031_), .B(_03946_), .Y(_03947_));
NAND_g _24725_ (.A(_03945_), .B(_03947_), .Y(_03948_));
NAND_g _24726_ (.A(cpuregs[15][7]), .B(_00008_[2]), .Y(_03949_));
NAND_g _24727_ (.A(cpuregs[11][7]), .B(_09032_), .Y(_03950_));
AND_g _24728_ (.A(_00008_[1]), .B(_03950_), .Y(_03951_));
NAND_g _24729_ (.A(_03949_), .B(_03951_), .Y(_03952_));
NAND_g _24730_ (.A(_03948_), .B(_03952_), .Y(_03953_));
NAND_g _24731_ (.A(_00008_[0]), .B(_03953_), .Y(_03954_));
NAND_g _24732_ (.A(cpuregs[8][7]), .B(_09032_), .Y(_03955_));
NAND_g _24733_ (.A(cpuregs[12][7]), .B(_00008_[2]), .Y(_03956_));
AND_g _24734_ (.A(_09031_), .B(_03956_), .Y(_03957_));
NAND_g _24735_ (.A(_03955_), .B(_03957_), .Y(_03958_));
NAND_g _24736_ (.A(cpuregs[10][7]), .B(_09032_), .Y(_03959_));
NAND_g _24737_ (.A(cpuregs[14][7]), .B(_00008_[2]), .Y(_03960_));
AND_g _24738_ (.A(_00008_[1]), .B(_03960_), .Y(_03961_));
NAND_g _24739_ (.A(_03959_), .B(_03961_), .Y(_03962_));
NAND_g _24740_ (.A(_03958_), .B(_03962_), .Y(_03963_));
NAND_g _24741_ (.A(_09030_), .B(_03963_), .Y(_03964_));
NAND_g _24742_ (.A(_03954_), .B(_03964_), .Y(_03965_));
AND_g _24743_ (.A(_00008_[3]), .B(_03965_), .Y(_03966_));
NOR_g _24744_ (.A(_00008_[4]), .B(_03966_), .Y(_03967_));
NAND_g _24745_ (.A(_03944_), .B(_03967_), .Y(_03968_));
NAND_g _24746_ (.A(_03922_), .B(_03968_), .Y(_03969_));
NAND_g _24747_ (.A(_14624_), .B(_03969_), .Y(_03970_));
NAND_g _24748_ (.A(_03876_), .B(_03970_), .Y(_03971_));
NAND_g _24749_ (.A(_10595_), .B(_03971_), .Y(_03972_));
NAND_g _24750_ (.A(pcpi_rs1[6]), .B(_14481_), .Y(_03973_));
AND_g _24751_ (.A(_03641_), .B(_03973_), .Y(_03974_));
NAND_g _24752_ (.A(pcpi_rs1[11]), .B(_14482_), .Y(_03975_));
AND_g _24753_ (.A(_03638_), .B(_03975_), .Y(_03976_));
NAND_g _24754_ (.A(_13880_), .B(_03976_), .Y(_03977_));
NAND_g _24755_ (.A(_13879_), .B(_03974_), .Y(_03978_));
AND_g _24756_ (.A(_13883_), .B(_03978_), .Y(_03979_));
NAND_g _24757_ (.A(_03977_), .B(_03979_), .Y(_03980_));
AND_g _24758_ (.A(_03972_), .B(_03980_), .Y(_03981_));
AND_g _24759_ (.A(_03875_), .B(_03981_), .Y(_03982_));
NOR_g _24760_ (.A(pcpi_rs1[7]), .B(_14488_), .Y(_03983_));
AND_g _24761_ (.A(_14488_), .B(_03982_), .Y(_03984_));
NOR_g _24762_ (.A(_03983_), .B(_03984_), .Y(_01025_));
XOR_g _24763_ (.A(_14536_), .B(_14566_), .Y(_03985_));
NAND_g _24764_ (.A(_14614_), .B(_03985_), .Y(_03986_));
NAND_g _24765_ (.A(reg_pc[8]), .B(_14617_), .Y(_03987_));
NAND_g _24766_ (.A(cpuregs[13][8]), .B(_00008_[2]), .Y(_03988_));
NAND_g _24767_ (.A(cpuregs[9][8]), .B(_09032_), .Y(_03989_));
NAND_g _24768_ (.A(_03988_), .B(_03989_), .Y(_03990_));
NAND_g _24769_ (.A(_00008_[0]), .B(_03990_), .Y(_03991_));
NAND_g _24770_ (.A(cpuregs[12][8]), .B(_00008_[2]), .Y(_03992_));
NAND_g _24771_ (.A(cpuregs[8][8]), .B(_09032_), .Y(_03993_));
AND_g _24772_ (.A(_03992_), .B(_03993_), .Y(_03994_));
NOR_g _24773_ (.A(_00008_[0]), .B(_03994_), .Y(_03995_));
NAND_g _24774_ (.A(_08906_), .B(_00008_[2]), .Y(_03996_));
NOR_g _24775_ (.A(cpuregs[0][8]), .B(_00008_[2]), .Y(_03997_));
NOR_g _24776_ (.A(_00008_[0]), .B(_03997_), .Y(_03998_));
NAND_g _24777_ (.A(_03996_), .B(_03998_), .Y(_03999_));
NAND_g _24778_ (.A(_08948_), .B(_00008_[2]), .Y(_04000_));
NOR_g _24779_ (.A(cpuregs[1][8]), .B(_00008_[2]), .Y(_04001_));
NOR_g _24780_ (.A(_09030_), .B(_04001_), .Y(_04002_));
NAND_g _24781_ (.A(_04000_), .B(_04002_), .Y(_04003_));
NAND_g _24782_ (.A(cpuregs[11][8]), .B(_09032_), .Y(_04004_));
NAND_g _24783_ (.A(cpuregs[15][8]), .B(_00008_[2]), .Y(_04005_));
NAND_g _24784_ (.A(_04004_), .B(_04005_), .Y(_04006_));
AND_g _24785_ (.A(_00008_[0]), .B(_04006_), .Y(_04007_));
NAND_g _24786_ (.A(cpuregs[14][8]), .B(_00008_[2]), .Y(_04008_));
NAND_g _24787_ (.A(cpuregs[10][8]), .B(_09032_), .Y(_04009_));
AND_g _24788_ (.A(_04008_), .B(_04009_), .Y(_04010_));
NOR_g _24789_ (.A(_00008_[0]), .B(_04010_), .Y(_04011_));
NOR_g _24790_ (.A(_04007_), .B(_04011_), .Y(_04012_));
NAND_g _24791_ (.A(_09005_), .B(_00008_[2]), .Y(_04013_));
NOR_g _24792_ (.A(cpuregs[2][8]), .B(_00008_[2]), .Y(_04014_));
NOR_g _24793_ (.A(_00008_[0]), .B(_04014_), .Y(_04015_));
NAND_g _24794_ (.A(_04013_), .B(_04015_), .Y(_04016_));
NAND_g _24795_ (.A(_08965_), .B(_00008_[2]), .Y(_04017_));
NOR_g _24796_ (.A(cpuregs[3][8]), .B(_00008_[2]), .Y(_04018_));
NOR_g _24797_ (.A(_09030_), .B(_04018_), .Y(_04019_));
NAND_g _24798_ (.A(_04017_), .B(_04019_), .Y(_04020_));
AND_g _24799_ (.A(_04016_), .B(_04020_), .Y(_04021_));
AND_g _24800_ (.A(_09031_), .B(_03999_), .Y(_04022_));
NAND_g _24801_ (.A(_04003_), .B(_04022_), .Y(_04023_));
NAND_g _24802_ (.A(_00008_[1]), .B(_04021_), .Y(_04024_));
AND_g _24803_ (.A(_04023_), .B(_04024_), .Y(_04025_));
NAND_g _24804_ (.A(_09033_), .B(_04025_), .Y(_04026_));
NAND_g _24805_ (.A(_00008_[1]), .B(_04012_), .Y(_04027_));
NOR_g _24806_ (.A(_00008_[1]), .B(_03995_), .Y(_04028_));
NAND_g _24807_ (.A(_03991_), .B(_04028_), .Y(_04029_));
AND_g _24808_ (.A(_00008_[3]), .B(_04029_), .Y(_04030_));
AND_g _24809_ (.A(_04027_), .B(_04030_), .Y(_04031_));
NOR_g _24810_ (.A(_00008_[4]), .B(_04031_), .Y(_04032_));
NAND_g _24811_ (.A(_04026_), .B(_04032_), .Y(_04033_));
NAND_g _24812_ (.A(_08887_), .B(_00008_[2]), .Y(_04034_));
NOR_g _24813_ (.A(cpuregs[19][8]), .B(_00008_[2]), .Y(_04035_));
NOR_g _24814_ (.A(cpuregs[18][8]), .B(_00008_[2]), .Y(_04036_));
NOR_g _24815_ (.A(cpuregs[22][8]), .B(_09032_), .Y(_04037_));
NOR_g _24816_ (.A(_04036_), .B(_04037_), .Y(_04038_));
NOR_g _24817_ (.A(_09030_), .B(_04035_), .Y(_04039_));
NAND_g _24818_ (.A(_04034_), .B(_04039_), .Y(_04040_));
NAND_g _24819_ (.A(_09030_), .B(_04038_), .Y(_04041_));
AND_g _24820_ (.A(_04040_), .B(_04041_), .Y(_04042_));
NAND_g _24821_ (.A(_00008_[1]), .B(_04042_), .Y(_04043_));
NOR_g _24822_ (.A(cpuregs[17][8]), .B(_00008_[2]), .Y(_04044_));
NAND_g _24823_ (.A(_08986_), .B(_00008_[2]), .Y(_04045_));
NOR_g _24824_ (.A(cpuregs[16][8]), .B(_00008_[2]), .Y(_04046_));
NOR_g _24825_ (.A(cpuregs[20][8]), .B(_09032_), .Y(_04047_));
NOR_g _24826_ (.A(_04046_), .B(_04047_), .Y(_04048_));
NOR_g _24827_ (.A(_09030_), .B(_04044_), .Y(_04049_));
NAND_g _24828_ (.A(_04045_), .B(_04049_), .Y(_04050_));
NAND_g _24829_ (.A(_09030_), .B(_04048_), .Y(_04051_));
AND_g _24830_ (.A(_04050_), .B(_04051_), .Y(_04052_));
NAND_g _24831_ (.A(_09031_), .B(_04052_), .Y(_04053_));
NAND_g _24832_ (.A(_04043_), .B(_04053_), .Y(_04054_));
NAND_g _24833_ (.A(_09033_), .B(_04054_), .Y(_04055_));
NAND_g _24834_ (.A(cpuregs[25][8]), .B(_09031_), .Y(_04056_));
NAND_g _24835_ (.A(cpuregs[27][8]), .B(_00008_[1]), .Y(_04057_));
AND_g _24836_ (.A(_09032_), .B(_04057_), .Y(_04058_));
NAND_g _24837_ (.A(_04056_), .B(_04058_), .Y(_04059_));
NAND_g _24838_ (.A(cpuregs[29][8]), .B(_09031_), .Y(_04060_));
NAND_g _24839_ (.A(cpuregs[31][8]), .B(_00008_[1]), .Y(_04061_));
AND_g _24840_ (.A(_00008_[2]), .B(_04061_), .Y(_04062_));
NAND_g _24841_ (.A(_04060_), .B(_04062_), .Y(_04063_));
NAND_g _24842_ (.A(_04059_), .B(_04063_), .Y(_04064_));
NAND_g _24843_ (.A(_00008_[0]), .B(_04064_), .Y(_04065_));
NAND_g _24844_ (.A(cpuregs[24][8]), .B(_09031_), .Y(_04066_));
NAND_g _24845_ (.A(cpuregs[26][8]), .B(_00008_[1]), .Y(_04067_));
AND_g _24846_ (.A(_09032_), .B(_04067_), .Y(_04068_));
NAND_g _24847_ (.A(_04066_), .B(_04068_), .Y(_04069_));
NAND_g _24848_ (.A(cpuregs[28][8]), .B(_09031_), .Y(_04070_));
NAND_g _24849_ (.A(cpuregs[30][8]), .B(_00008_[1]), .Y(_04071_));
AND_g _24850_ (.A(_00008_[2]), .B(_04071_), .Y(_04072_));
NAND_g _24851_ (.A(_04070_), .B(_04072_), .Y(_04073_));
NAND_g _24852_ (.A(_04069_), .B(_04073_), .Y(_04074_));
NAND_g _24853_ (.A(_09030_), .B(_04074_), .Y(_04075_));
NAND_g _24854_ (.A(_04065_), .B(_04075_), .Y(_04076_));
NAND_g _24855_ (.A(_00008_[3]), .B(_04076_), .Y(_04077_));
NAND_g _24856_ (.A(_04055_), .B(_04077_), .Y(_04078_));
NAND_g _24857_ (.A(_00008_[4]), .B(_04078_), .Y(_04079_));
AND_g _24858_ (.A(_14624_), .B(_04033_), .Y(_04080_));
NAND_g _24859_ (.A(_04079_), .B(_04080_), .Y(_04081_));
NAND_g _24860_ (.A(_03987_), .B(_04081_), .Y(_04082_));
NAND_g _24861_ (.A(_10595_), .B(_04082_), .Y(_04083_));
NAND_g _24862_ (.A(pcpi_rs1[7]), .B(_14481_), .Y(_04084_));
AND_g _24863_ (.A(_03753_), .B(_04084_), .Y(_04085_));
NAND_g _24864_ (.A(pcpi_rs1[12]), .B(_14482_), .Y(_04086_));
AND_g _24865_ (.A(_03750_), .B(_04086_), .Y(_04087_));
NAND_g _24866_ (.A(_13880_), .B(_04087_), .Y(_04088_));
NAND_g _24867_ (.A(_13879_), .B(_04085_), .Y(_04089_));
NOR_g _24868_ (.A(pcpi_rs1[8]), .B(_14488_), .Y(_04090_));
AND_g _24869_ (.A(_13883_), .B(_04088_), .Y(_04091_));
NAND_g _24870_ (.A(_04089_), .B(_04091_), .Y(_04092_));
AND_g _24871_ (.A(_04083_), .B(_04092_), .Y(_04093_));
AND_g _24872_ (.A(_14488_), .B(_04093_), .Y(_04094_));
AND_g _24873_ (.A(_03986_), .B(_04094_), .Y(_04095_));
NOR_g _24874_ (.A(_04090_), .B(_04095_), .Y(_01026_));
NOR_g _24875_ (.A(pcpi_rs1[9]), .B(_14488_), .Y(_04096_));
NAND_g _24876_ (.A(reg_pc[9]), .B(_14617_), .Y(_04097_));
NAND_g _24877_ (.A(cpuregs[13][9]), .B(_00008_[2]), .Y(_04098_));
NAND_g _24878_ (.A(cpuregs[9][9]), .B(_09032_), .Y(_04099_));
NAND_g _24879_ (.A(_04098_), .B(_04099_), .Y(_04100_));
NAND_g _24880_ (.A(_00008_[0]), .B(_04100_), .Y(_04101_));
NAND_g _24881_ (.A(cpuregs[12][9]), .B(_00008_[2]), .Y(_04102_));
NAND_g _24882_ (.A(cpuregs[8][9]), .B(_09032_), .Y(_04103_));
AND_g _24883_ (.A(_04102_), .B(_04103_), .Y(_04104_));
NOR_g _24884_ (.A(_00008_[0]), .B(_04104_), .Y(_04105_));
NAND_g _24885_ (.A(_08907_), .B(_00008_[2]), .Y(_04106_));
NOR_g _24886_ (.A(cpuregs[0][9]), .B(_00008_[2]), .Y(_04107_));
NOR_g _24887_ (.A(_00008_[0]), .B(_04107_), .Y(_04108_));
NAND_g _24888_ (.A(_04106_), .B(_04108_), .Y(_04109_));
NAND_g _24889_ (.A(_08949_), .B(_00008_[2]), .Y(_04110_));
NOR_g _24890_ (.A(cpuregs[1][9]), .B(_00008_[2]), .Y(_04111_));
NOR_g _24891_ (.A(_09030_), .B(_04111_), .Y(_04112_));
NAND_g _24892_ (.A(_04110_), .B(_04112_), .Y(_04113_));
NAND_g _24893_ (.A(cpuregs[11][9]), .B(_09032_), .Y(_04114_));
NAND_g _24894_ (.A(cpuregs[15][9]), .B(_00008_[2]), .Y(_04115_));
NAND_g _24895_ (.A(_04114_), .B(_04115_), .Y(_04116_));
AND_g _24896_ (.A(_00008_[0]), .B(_04116_), .Y(_04117_));
NAND_g _24897_ (.A(cpuregs[14][9]), .B(_00008_[2]), .Y(_04118_));
NAND_g _24898_ (.A(cpuregs[10][9]), .B(_09032_), .Y(_04119_));
AND_g _24899_ (.A(_04118_), .B(_04119_), .Y(_04120_));
NOR_g _24900_ (.A(_00008_[0]), .B(_04120_), .Y(_04121_));
NOR_g _24901_ (.A(_04117_), .B(_04121_), .Y(_04122_));
NAND_g _24902_ (.A(_09006_), .B(_00008_[2]), .Y(_04123_));
NOR_g _24903_ (.A(cpuregs[2][9]), .B(_00008_[2]), .Y(_04124_));
NOR_g _24904_ (.A(_00008_[0]), .B(_04124_), .Y(_04125_));
NAND_g _24905_ (.A(_04123_), .B(_04125_), .Y(_04126_));
NAND_g _24906_ (.A(_08966_), .B(_00008_[2]), .Y(_04127_));
NOR_g _24907_ (.A(cpuregs[3][9]), .B(_00008_[2]), .Y(_04128_));
NOR_g _24908_ (.A(_09030_), .B(_04128_), .Y(_04129_));
NAND_g _24909_ (.A(_04127_), .B(_04129_), .Y(_04130_));
AND_g _24910_ (.A(_04126_), .B(_04130_), .Y(_04131_));
AND_g _24911_ (.A(_09031_), .B(_04109_), .Y(_04132_));
NAND_g _24912_ (.A(_04113_), .B(_04132_), .Y(_04133_));
NAND_g _24913_ (.A(_00008_[1]), .B(_04131_), .Y(_04134_));
AND_g _24914_ (.A(_04133_), .B(_04134_), .Y(_04135_));
NAND_g _24915_ (.A(_09033_), .B(_04135_), .Y(_04136_));
NAND_g _24916_ (.A(_00008_[1]), .B(_04122_), .Y(_04137_));
NOR_g _24917_ (.A(_00008_[1]), .B(_04105_), .Y(_04138_));
NAND_g _24918_ (.A(_04101_), .B(_04138_), .Y(_04139_));
AND_g _24919_ (.A(_00008_[3]), .B(_04139_), .Y(_04140_));
AND_g _24920_ (.A(_04137_), .B(_04140_), .Y(_04141_));
NOR_g _24921_ (.A(_00008_[4]), .B(_04141_), .Y(_04142_));
NAND_g _24922_ (.A(_04136_), .B(_04142_), .Y(_04143_));
NAND_g _24923_ (.A(_08888_), .B(_00008_[2]), .Y(_04144_));
NOR_g _24924_ (.A(cpuregs[19][9]), .B(_00008_[2]), .Y(_04145_));
NOR_g _24925_ (.A(cpuregs[18][9]), .B(_00008_[2]), .Y(_04146_));
NOR_g _24926_ (.A(cpuregs[22][9]), .B(_09032_), .Y(_04147_));
NOR_g _24927_ (.A(_04146_), .B(_04147_), .Y(_04148_));
NOR_g _24928_ (.A(_09030_), .B(_04145_), .Y(_04149_));
NAND_g _24929_ (.A(_04144_), .B(_04149_), .Y(_04150_));
NAND_g _24930_ (.A(_09030_), .B(_04148_), .Y(_04151_));
AND_g _24931_ (.A(_04150_), .B(_04151_), .Y(_04152_));
NAND_g _24932_ (.A(_00008_[1]), .B(_04152_), .Y(_04153_));
NOR_g _24933_ (.A(cpuregs[17][9]), .B(_00008_[2]), .Y(_04154_));
NAND_g _24934_ (.A(_08987_), .B(_00008_[2]), .Y(_04155_));
NOR_g _24935_ (.A(cpuregs[16][9]), .B(_00008_[2]), .Y(_04156_));
NOR_g _24936_ (.A(cpuregs[20][9]), .B(_09032_), .Y(_04157_));
NOR_g _24937_ (.A(_04156_), .B(_04157_), .Y(_04158_));
NOR_g _24938_ (.A(_09030_), .B(_04154_), .Y(_04159_));
NAND_g _24939_ (.A(_04155_), .B(_04159_), .Y(_04160_));
NAND_g _24940_ (.A(_09030_), .B(_04158_), .Y(_04161_));
AND_g _24941_ (.A(_04160_), .B(_04161_), .Y(_04162_));
NAND_g _24942_ (.A(_09031_), .B(_04162_), .Y(_04163_));
NAND_g _24943_ (.A(_04153_), .B(_04163_), .Y(_04164_));
NAND_g _24944_ (.A(_09033_), .B(_04164_), .Y(_04165_));
NAND_g _24945_ (.A(cpuregs[25][9]), .B(_09031_), .Y(_04166_));
NAND_g _24946_ (.A(cpuregs[27][9]), .B(_00008_[1]), .Y(_04167_));
AND_g _24947_ (.A(_09032_), .B(_04167_), .Y(_04168_));
NAND_g _24948_ (.A(_04166_), .B(_04168_), .Y(_04169_));
NAND_g _24949_ (.A(cpuregs[29][9]), .B(_09031_), .Y(_04170_));
NAND_g _24950_ (.A(cpuregs[31][9]), .B(_00008_[1]), .Y(_04171_));
AND_g _24951_ (.A(_00008_[2]), .B(_04171_), .Y(_04172_));
NAND_g _24952_ (.A(_04170_), .B(_04172_), .Y(_04173_));
NAND_g _24953_ (.A(_04169_), .B(_04173_), .Y(_04174_));
NAND_g _24954_ (.A(_00008_[0]), .B(_04174_), .Y(_04175_));
NAND_g _24955_ (.A(cpuregs[24][9]), .B(_09031_), .Y(_04176_));
NAND_g _24956_ (.A(cpuregs[26][9]), .B(_00008_[1]), .Y(_04177_));
AND_g _24957_ (.A(_09032_), .B(_04177_), .Y(_04178_));
NAND_g _24958_ (.A(_04176_), .B(_04178_), .Y(_04179_));
NAND_g _24959_ (.A(cpuregs[28][9]), .B(_09031_), .Y(_04180_));
NAND_g _24960_ (.A(cpuregs[30][9]), .B(_00008_[1]), .Y(_04181_));
AND_g _24961_ (.A(_00008_[2]), .B(_04181_), .Y(_04182_));
NAND_g _24962_ (.A(_04180_), .B(_04182_), .Y(_04183_));
NAND_g _24963_ (.A(_04179_), .B(_04183_), .Y(_04184_));
NAND_g _24964_ (.A(_09030_), .B(_04184_), .Y(_04185_));
NAND_g _24965_ (.A(_04175_), .B(_04185_), .Y(_04186_));
NAND_g _24966_ (.A(_00008_[3]), .B(_04186_), .Y(_04187_));
NAND_g _24967_ (.A(_04165_), .B(_04187_), .Y(_04188_));
NAND_g _24968_ (.A(_00008_[4]), .B(_04188_), .Y(_04189_));
AND_g _24969_ (.A(_14624_), .B(_04143_), .Y(_04190_));
NAND_g _24970_ (.A(_04189_), .B(_04190_), .Y(_04191_));
NAND_g _24971_ (.A(_04097_), .B(_04191_), .Y(_04192_));
NAND_g _24972_ (.A(_10595_), .B(_04192_), .Y(_04193_));
NAND_g _24973_ (.A(pcpi_rs1[8]), .B(_14481_), .Y(_04194_));
NAND_g _24974_ (.A(_03862_), .B(_04194_), .Y(_04195_));
NAND_g _24975_ (.A(_13879_), .B(_04195_), .Y(_04196_));
NAND_g _24976_ (.A(pcpi_rs1[13]), .B(_14482_), .Y(_04197_));
NAND_g _24977_ (.A(_03860_), .B(_04197_), .Y(_04198_));
NAND_g _24978_ (.A(_13880_), .B(_04198_), .Y(_04199_));
NAND_g _24979_ (.A(_04196_), .B(_04199_), .Y(_04200_));
NAND_g _24980_ (.A(_13883_), .B(_04200_), .Y(_04201_));
AND_g _24981_ (.A(_14488_), .B(_04201_), .Y(_04202_));
AND_g _24982_ (.A(_04193_), .B(_04202_), .Y(_04203_));
XOR_g _24983_ (.A(decoded_imm[9]), .B(pcpi_rs1[9]), .Y(_04204_));
XNOR_g _24984_ (.A(_14568_), .B(_04204_), .Y(_04205_));
NAND_g _24985_ (.A(_14614_), .B(_04205_), .Y(_04206_));
AND_g _24986_ (.A(_04203_), .B(_04206_), .Y(_04207_));
NOR_g _24987_ (.A(_04096_), .B(_04207_), .Y(_01027_));
NOR_g _24988_ (.A(pcpi_rs1[10]), .B(_14488_), .Y(_04208_));
XOR_g _24989_ (.A(_14532_), .B(_14570_), .Y(_04209_));
NAND_g _24990_ (.A(_14614_), .B(_04209_), .Y(_04210_));
NAND_g _24991_ (.A(reg_pc[10]), .B(_14617_), .Y(_04211_));
NAND_g _24992_ (.A(cpuregs[7][10]), .B(_00008_[2]), .Y(_04212_));
NAND_g _24993_ (.A(cpuregs[3][10]), .B(_09032_), .Y(_04213_));
NAND_g _24994_ (.A(_04212_), .B(_04213_), .Y(_04214_));
NAND_g _24995_ (.A(_00008_[0]), .B(_04214_), .Y(_04215_));
NAND_g _24996_ (.A(cpuregs[6][10]), .B(_00008_[2]), .Y(_04216_));
NAND_g _24997_ (.A(cpuregs[2][10]), .B(_09032_), .Y(_04217_));
NAND_g _24998_ (.A(_04216_), .B(_04217_), .Y(_04218_));
NAND_g _24999_ (.A(_09030_), .B(_04218_), .Y(_04219_));
AND_g _25000_ (.A(_04215_), .B(_04219_), .Y(_04220_));
NAND_g _25001_ (.A(cpuregs[4][10]), .B(_00008_[2]), .Y(_04221_));
NAND_g _25002_ (.A(cpuregs[0][10]), .B(_09032_), .Y(_04222_));
AND_g _25003_ (.A(_04221_), .B(_04222_), .Y(_04223_));
NAND_g _25004_ (.A(_09030_), .B(_04223_), .Y(_04224_));
NAND_g _25005_ (.A(cpuregs[5][10]), .B(_00008_[2]), .Y(_04225_));
NAND_g _25006_ (.A(cpuregs[1][10]), .B(_09032_), .Y(_04226_));
AND_g _25007_ (.A(_00008_[0]), .B(_04226_), .Y(_04227_));
NAND_g _25008_ (.A(_04225_), .B(_04227_), .Y(_04228_));
NAND_g _25009_ (.A(cpuregs[11][10]), .B(_09032_), .Y(_04229_));
NAND_g _25010_ (.A(cpuregs[15][10]), .B(_00008_[2]), .Y(_04230_));
NAND_g _25011_ (.A(_04229_), .B(_04230_), .Y(_04231_));
AND_g _25012_ (.A(_00008_[0]), .B(_04231_), .Y(_04232_));
NAND_g _25013_ (.A(cpuregs[14][10]), .B(_00008_[2]), .Y(_04233_));
NAND_g _25014_ (.A(cpuregs[10][10]), .B(_09032_), .Y(_04234_));
AND_g _25015_ (.A(_04233_), .B(_04234_), .Y(_04235_));
NOR_g _25016_ (.A(_00008_[0]), .B(_04235_), .Y(_04236_));
NOR_g _25017_ (.A(_04232_), .B(_04236_), .Y(_04237_));
NAND_g _25018_ (.A(_08881_), .B(_00008_[2]), .Y(_04238_));
NOR_g _25019_ (.A(cpuregs[8][10]), .B(_00008_[2]), .Y(_04239_));
NOR_g _25020_ (.A(_00008_[0]), .B(_04239_), .Y(_04240_));
NAND_g _25021_ (.A(_04238_), .B(_04240_), .Y(_04241_));
NAND_g _25022_ (.A(_08980_), .B(_09032_), .Y(_04242_));
NAND_g _25023_ (.A(_08929_), .B(_00008_[2]), .Y(_04243_));
AND_g _25024_ (.A(_00008_[0]), .B(_04243_), .Y(_04244_));
NAND_g _25025_ (.A(_04242_), .B(_04244_), .Y(_04245_));
NAND_g _25026_ (.A(_04241_), .B(_04245_), .Y(_04246_));
NAND_g _25027_ (.A(_00008_[3]), .B(_04246_), .Y(_04247_));
AND_g _25028_ (.A(_09033_), .B(_04228_), .Y(_04248_));
NAND_g _25029_ (.A(_04224_), .B(_04248_), .Y(_04249_));
NAND_g _25030_ (.A(_04247_), .B(_04249_), .Y(_04250_));
NAND_g _25031_ (.A(_09031_), .B(_04250_), .Y(_04251_));
NAND_g _25032_ (.A(_00008_[3]), .B(_04237_), .Y(_04252_));
NAND_g _25033_ (.A(_09033_), .B(_04220_), .Y(_04253_));
AND_g _25034_ (.A(_04252_), .B(_04253_), .Y(_04254_));
AND_g _25035_ (.A(_00008_[1]), .B(_04254_), .Y(_04255_));
NOR_g _25036_ (.A(_00008_[4]), .B(_04255_), .Y(_04256_));
NAND_g _25037_ (.A(_04251_), .B(_04256_), .Y(_04257_));
NAND_g _25038_ (.A(cpuregs[25][10]), .B(_09032_), .Y(_04258_));
NAND_g _25039_ (.A(cpuregs[29][10]), .B(_00008_[2]), .Y(_04259_));
AND_g _25040_ (.A(_09031_), .B(_04259_), .Y(_04260_));
NAND_g _25041_ (.A(_04258_), .B(_04260_), .Y(_04261_));
NAND_g _25042_ (.A(cpuregs[31][10]), .B(_00008_[2]), .Y(_04262_));
NAND_g _25043_ (.A(cpuregs[27][10]), .B(_09032_), .Y(_04263_));
AND_g _25044_ (.A(_00008_[1]), .B(_04263_), .Y(_04264_));
NAND_g _25045_ (.A(_04262_), .B(_04264_), .Y(_04265_));
NAND_g _25046_ (.A(_04261_), .B(_04265_), .Y(_04266_));
NAND_g _25047_ (.A(_00008_[0]), .B(_04266_), .Y(_04267_));
NAND_g _25048_ (.A(cpuregs[24][10]), .B(_09032_), .Y(_04268_));
NAND_g _25049_ (.A(cpuregs[28][10]), .B(_00008_[2]), .Y(_04269_));
AND_g _25050_ (.A(_09031_), .B(_04269_), .Y(_04270_));
NAND_g _25051_ (.A(_04268_), .B(_04270_), .Y(_04271_));
NAND_g _25052_ (.A(cpuregs[26][10]), .B(_09032_), .Y(_04272_));
NAND_g _25053_ (.A(cpuregs[30][10]), .B(_00008_[2]), .Y(_04273_));
AND_g _25054_ (.A(_00008_[1]), .B(_04273_), .Y(_04274_));
NAND_g _25055_ (.A(_04272_), .B(_04274_), .Y(_04275_));
NAND_g _25056_ (.A(_04271_), .B(_04275_), .Y(_04276_));
NAND_g _25057_ (.A(_09030_), .B(_04276_), .Y(_04277_));
NAND_g _25058_ (.A(_04267_), .B(_04277_), .Y(_04278_));
NAND_g _25059_ (.A(_00008_[3]), .B(_04278_), .Y(_04279_));
NAND_g _25060_ (.A(cpuregs[17][10]), .B(_09031_), .Y(_04280_));
NAND_g _25061_ (.A(cpuregs[19][10]), .B(_00008_[1]), .Y(_04281_));
AND_g _25062_ (.A(_09032_), .B(_04281_), .Y(_04282_));
NAND_g _25063_ (.A(_04280_), .B(_04282_), .Y(_04283_));
NAND_g _25064_ (.A(cpuregs[21][10]), .B(_09031_), .Y(_04284_));
NAND_g _25065_ (.A(cpuregs[23][10]), .B(_00008_[1]), .Y(_04285_));
AND_g _25066_ (.A(_00008_[2]), .B(_04285_), .Y(_04286_));
NAND_g _25067_ (.A(_04284_), .B(_04286_), .Y(_04287_));
NAND_g _25068_ (.A(_04283_), .B(_04287_), .Y(_04288_));
NAND_g _25069_ (.A(_00008_[0]), .B(_04288_), .Y(_04289_));
NAND_g _25070_ (.A(cpuregs[16][10]), .B(_09031_), .Y(_04290_));
NAND_g _25071_ (.A(cpuregs[18][10]), .B(_00008_[1]), .Y(_04291_));
AND_g _25072_ (.A(_09032_), .B(_04291_), .Y(_04292_));
NAND_g _25073_ (.A(_04290_), .B(_04292_), .Y(_04293_));
NAND_g _25074_ (.A(cpuregs[20][10]), .B(_09031_), .Y(_04294_));
NAND_g _25075_ (.A(cpuregs[22][10]), .B(_00008_[1]), .Y(_04295_));
AND_g _25076_ (.A(_00008_[2]), .B(_04295_), .Y(_04296_));
NAND_g _25077_ (.A(_04294_), .B(_04296_), .Y(_04297_));
NAND_g _25078_ (.A(_04293_), .B(_04297_), .Y(_04298_));
NAND_g _25079_ (.A(_09030_), .B(_04298_), .Y(_04299_));
NAND_g _25080_ (.A(_04289_), .B(_04299_), .Y(_04300_));
AND_g _25081_ (.A(_09033_), .B(_04300_), .Y(_04301_));
NOT_g _25082_ (.A(_04301_), .Y(_04302_));
NAND_g _25083_ (.A(_04279_), .B(_04302_), .Y(_04303_));
NAND_g _25084_ (.A(_00008_[4]), .B(_04303_), .Y(_04304_));
AND_g _25085_ (.A(_14624_), .B(_04257_), .Y(_04305_));
NAND_g _25086_ (.A(_04304_), .B(_04305_), .Y(_04306_));
NAND_g _25087_ (.A(_04211_), .B(_04306_), .Y(_04307_));
NAND_g _25088_ (.A(_10595_), .B(_04307_), .Y(_04308_));
NAND_g _25089_ (.A(pcpi_rs1[9]), .B(_14481_), .Y(_04309_));
AND_g _25090_ (.A(_03975_), .B(_04309_), .Y(_04310_));
NAND_g _25091_ (.A(_13879_), .B(_04310_), .Y(_04311_));
NAND_g _25092_ (.A(pcpi_rs1[14]), .B(_14482_), .Y(_04312_));
AND_g _25093_ (.A(_03973_), .B(_04312_), .Y(_04313_));
NAND_g _25094_ (.A(_13880_), .B(_04313_), .Y(_04314_));
AND_g _25095_ (.A(_04311_), .B(_04314_), .Y(_04315_));
NAND_g _25096_ (.A(_13883_), .B(_04315_), .Y(_04316_));
AND_g _25097_ (.A(_14488_), .B(_04308_), .Y(_04317_));
AND_g _25098_ (.A(_04316_), .B(_04317_), .Y(_04318_));
AND_g _25099_ (.A(_04210_), .B(_04318_), .Y(_04319_));
NOR_g _25100_ (.A(_04208_), .B(_04319_), .Y(_01028_));
NOR_g _25101_ (.A(pcpi_rs1[11]), .B(_14488_), .Y(_04320_));
XOR_g _25102_ (.A(decoded_imm[11]), .B(pcpi_rs1[11]), .Y(_04321_));
XNOR_g _25103_ (.A(_14572_), .B(_04321_), .Y(_04322_));
NAND_g _25104_ (.A(_14614_), .B(_04322_), .Y(_04323_));
NAND_g _25105_ (.A(reg_pc[11]), .B(_14617_), .Y(_04324_));
NAND_g _25106_ (.A(cpuregs[13][11]), .B(_00008_[2]), .Y(_04325_));
NAND_g _25107_ (.A(cpuregs[9][11]), .B(_09032_), .Y(_04326_));
NAND_g _25108_ (.A(_04325_), .B(_04326_), .Y(_04327_));
NAND_g _25109_ (.A(_00008_[0]), .B(_04327_), .Y(_04328_));
NAND_g _25110_ (.A(cpuregs[12][11]), .B(_00008_[2]), .Y(_04329_));
NAND_g _25111_ (.A(cpuregs[8][11]), .B(_09032_), .Y(_04330_));
AND_g _25112_ (.A(_04329_), .B(_04330_), .Y(_04331_));
NOR_g _25113_ (.A(_00008_[0]), .B(_04331_), .Y(_04332_));
NAND_g _25114_ (.A(_08908_), .B(_00008_[2]), .Y(_04333_));
NOR_g _25115_ (.A(cpuregs[0][11]), .B(_00008_[2]), .Y(_04334_));
NOR_g _25116_ (.A(_00008_[0]), .B(_04334_), .Y(_04335_));
NAND_g _25117_ (.A(_04333_), .B(_04335_), .Y(_04336_));
NAND_g _25118_ (.A(_08950_), .B(_00008_[2]), .Y(_04337_));
NOR_g _25119_ (.A(cpuregs[1][11]), .B(_00008_[2]), .Y(_04338_));
NOR_g _25120_ (.A(_09030_), .B(_04338_), .Y(_04339_));
NAND_g _25121_ (.A(_04337_), .B(_04339_), .Y(_04340_));
NAND_g _25122_ (.A(cpuregs[11][11]), .B(_09032_), .Y(_04341_));
NAND_g _25123_ (.A(cpuregs[15][11]), .B(_00008_[2]), .Y(_04342_));
NAND_g _25124_ (.A(_04341_), .B(_04342_), .Y(_04343_));
AND_g _25125_ (.A(_00008_[0]), .B(_04343_), .Y(_04344_));
NAND_g _25126_ (.A(cpuregs[14][11]), .B(_00008_[2]), .Y(_04345_));
NAND_g _25127_ (.A(cpuregs[10][11]), .B(_09032_), .Y(_04346_));
AND_g _25128_ (.A(_04345_), .B(_04346_), .Y(_04347_));
NOR_g _25129_ (.A(_00008_[0]), .B(_04347_), .Y(_04348_));
NOR_g _25130_ (.A(_04344_), .B(_04348_), .Y(_04349_));
NAND_g _25131_ (.A(_09007_), .B(_00008_[2]), .Y(_04350_));
NOR_g _25132_ (.A(cpuregs[2][11]), .B(_00008_[2]), .Y(_04351_));
NOR_g _25133_ (.A(_00008_[0]), .B(_04351_), .Y(_04352_));
NAND_g _25134_ (.A(_04350_), .B(_04352_), .Y(_04353_));
NAND_g _25135_ (.A(_08967_), .B(_00008_[2]), .Y(_04354_));
NOR_g _25136_ (.A(cpuregs[3][11]), .B(_00008_[2]), .Y(_04355_));
NOR_g _25137_ (.A(_09030_), .B(_04355_), .Y(_04356_));
NAND_g _25138_ (.A(_04354_), .B(_04356_), .Y(_04357_));
AND_g _25139_ (.A(_04353_), .B(_04357_), .Y(_04358_));
AND_g _25140_ (.A(_09031_), .B(_04336_), .Y(_04359_));
NAND_g _25141_ (.A(_04340_), .B(_04359_), .Y(_04360_));
NAND_g _25142_ (.A(_00008_[1]), .B(_04358_), .Y(_04361_));
AND_g _25143_ (.A(_04360_), .B(_04361_), .Y(_04362_));
NAND_g _25144_ (.A(_09033_), .B(_04362_), .Y(_04363_));
NAND_g _25145_ (.A(_00008_[1]), .B(_04349_), .Y(_04364_));
NOR_g _25146_ (.A(_00008_[1]), .B(_04332_), .Y(_04365_));
NAND_g _25147_ (.A(_04328_), .B(_04365_), .Y(_04366_));
AND_g _25148_ (.A(_00008_[3]), .B(_04366_), .Y(_04367_));
AND_g _25149_ (.A(_04364_), .B(_04367_), .Y(_04368_));
NOR_g _25150_ (.A(_00008_[4]), .B(_04368_), .Y(_04369_));
NAND_g _25151_ (.A(_04363_), .B(_04369_), .Y(_04370_));
NAND_g _25152_ (.A(_08890_), .B(_00008_[2]), .Y(_04371_));
NOR_g _25153_ (.A(cpuregs[19][11]), .B(_00008_[2]), .Y(_04372_));
NOR_g _25154_ (.A(cpuregs[18][11]), .B(_00008_[2]), .Y(_04373_));
AND_g _25155_ (.A(_08919_), .B(_00008_[2]), .Y(_04374_));
NOR_g _25156_ (.A(_04373_), .B(_04374_), .Y(_04375_));
NOR_g _25157_ (.A(_09030_), .B(_04372_), .Y(_04376_));
NAND_g _25158_ (.A(_04371_), .B(_04376_), .Y(_04377_));
NAND_g _25159_ (.A(_09030_), .B(_04375_), .Y(_04378_));
AND_g _25160_ (.A(_04377_), .B(_04378_), .Y(_04379_));
NAND_g _25161_ (.A(_00008_[1]), .B(_04379_), .Y(_04380_));
NOR_g _25162_ (.A(cpuregs[17][11]), .B(_00008_[2]), .Y(_04381_));
NAND_g _25163_ (.A(_08989_), .B(_00008_[2]), .Y(_04382_));
NOR_g _25164_ (.A(cpuregs[16][11]), .B(_00008_[2]), .Y(_04383_));
AND_g _25165_ (.A(_08845_), .B(_00008_[2]), .Y(_04384_));
NOR_g _25166_ (.A(_04383_), .B(_04384_), .Y(_04385_));
NOR_g _25167_ (.A(_09030_), .B(_04381_), .Y(_04386_));
NAND_g _25168_ (.A(_04382_), .B(_04386_), .Y(_04387_));
NAND_g _25169_ (.A(_09030_), .B(_04385_), .Y(_04388_));
AND_g _25170_ (.A(_04387_), .B(_04388_), .Y(_04389_));
NAND_g _25171_ (.A(_09031_), .B(_04389_), .Y(_04390_));
NAND_g _25172_ (.A(_04380_), .B(_04390_), .Y(_04391_));
NAND_g _25173_ (.A(_09033_), .B(_04391_), .Y(_04392_));
NAND_g _25174_ (.A(cpuregs[25][11]), .B(_09031_), .Y(_04393_));
NAND_g _25175_ (.A(cpuregs[27][11]), .B(_00008_[1]), .Y(_04394_));
AND_g _25176_ (.A(_09032_), .B(_04394_), .Y(_04395_));
NAND_g _25177_ (.A(_04393_), .B(_04395_), .Y(_04396_));
NAND_g _25178_ (.A(cpuregs[29][11]), .B(_09031_), .Y(_04397_));
NAND_g _25179_ (.A(cpuregs[31][11]), .B(_00008_[1]), .Y(_04398_));
AND_g _25180_ (.A(_00008_[2]), .B(_04398_), .Y(_04399_));
NAND_g _25181_ (.A(_04397_), .B(_04399_), .Y(_04400_));
NAND_g _25182_ (.A(_04396_), .B(_04400_), .Y(_04401_));
NAND_g _25183_ (.A(_00008_[0]), .B(_04401_), .Y(_04402_));
NAND_g _25184_ (.A(cpuregs[24][11]), .B(_09031_), .Y(_04403_));
NAND_g _25185_ (.A(cpuregs[26][11]), .B(_00008_[1]), .Y(_04404_));
AND_g _25186_ (.A(_09032_), .B(_04404_), .Y(_04405_));
NAND_g _25187_ (.A(_04403_), .B(_04405_), .Y(_04406_));
NAND_g _25188_ (.A(cpuregs[28][11]), .B(_09031_), .Y(_04407_));
NAND_g _25189_ (.A(cpuregs[30][11]), .B(_00008_[1]), .Y(_04408_));
AND_g _25190_ (.A(_00008_[2]), .B(_04408_), .Y(_04409_));
NAND_g _25191_ (.A(_04407_), .B(_04409_), .Y(_04410_));
NAND_g _25192_ (.A(_04406_), .B(_04410_), .Y(_04411_));
NAND_g _25193_ (.A(_09030_), .B(_04411_), .Y(_04412_));
NAND_g _25194_ (.A(_04402_), .B(_04412_), .Y(_04413_));
NAND_g _25195_ (.A(_00008_[3]), .B(_04413_), .Y(_04414_));
NAND_g _25196_ (.A(_04392_), .B(_04414_), .Y(_04415_));
NAND_g _25197_ (.A(_00008_[4]), .B(_04415_), .Y(_04416_));
AND_g _25198_ (.A(_14624_), .B(_04370_), .Y(_04417_));
NAND_g _25199_ (.A(_04416_), .B(_04417_), .Y(_04418_));
NAND_g _25200_ (.A(_04324_), .B(_04418_), .Y(_04419_));
NAND_g _25201_ (.A(_10595_), .B(_04419_), .Y(_04420_));
NAND_g _25202_ (.A(pcpi_rs1[10]), .B(_14481_), .Y(_04421_));
AND_g _25203_ (.A(_04086_), .B(_04421_), .Y(_04422_));
NAND_g _25204_ (.A(pcpi_rs1[15]), .B(_14482_), .Y(_04423_));
AND_g _25205_ (.A(_04084_), .B(_04423_), .Y(_04424_));
NAND_g _25206_ (.A(_13880_), .B(_04424_), .Y(_04425_));
NAND_g _25207_ (.A(_13879_), .B(_04422_), .Y(_04426_));
AND_g _25208_ (.A(_13883_), .B(_04425_), .Y(_04427_));
NAND_g _25209_ (.A(_04426_), .B(_04427_), .Y(_04428_));
AND_g _25210_ (.A(_14488_), .B(_04428_), .Y(_04429_));
AND_g _25211_ (.A(_04420_), .B(_04429_), .Y(_04430_));
AND_g _25212_ (.A(_04323_), .B(_04430_), .Y(_04431_));
NOR_g _25213_ (.A(_04320_), .B(_04431_), .Y(_01029_));
NOR_g _25214_ (.A(pcpi_rs1[12]), .B(_14488_), .Y(_04432_));
XOR_g _25215_ (.A(_14528_), .B(_14574_), .Y(_04433_));
NAND_g _25216_ (.A(_14614_), .B(_04433_), .Y(_04434_));
NAND_g _25217_ (.A(reg_pc[12]), .B(_14617_), .Y(_04435_));
NAND_g _25218_ (.A(_08968_), .B(_00008_[2]), .Y(_04436_));
NOR_g _25219_ (.A(cpuregs[3][12]), .B(_00008_[2]), .Y(_04437_));
NOR_g _25220_ (.A(_09030_), .B(_04437_), .Y(_04438_));
NAND_g _25221_ (.A(_04436_), .B(_04438_), .Y(_04439_));
NOR_g _25222_ (.A(cpuregs[2][12]), .B(_00008_[2]), .Y(_04440_));
AND_g _25223_ (.A(_09008_), .B(_00008_[2]), .Y(_04441_));
NOR_g _25224_ (.A(_04440_), .B(_04441_), .Y(_04442_));
NAND_g _25225_ (.A(_09030_), .B(_04442_), .Y(_04443_));
AND_g _25226_ (.A(_04439_), .B(_04443_), .Y(_04444_));
NAND_g _25227_ (.A(_08951_), .B(_00008_[2]), .Y(_04445_));
NOR_g _25228_ (.A(cpuregs[1][12]), .B(_00008_[2]), .Y(_04446_));
NOR_g _25229_ (.A(_09030_), .B(_04446_), .Y(_04447_));
NAND_g _25230_ (.A(_04445_), .B(_04447_), .Y(_04448_));
NOR_g _25231_ (.A(cpuregs[0][12]), .B(_00008_[2]), .Y(_04449_));
AND_g _25232_ (.A(_08909_), .B(_00008_[2]), .Y(_04450_));
NOR_g _25233_ (.A(_04449_), .B(_04450_), .Y(_04451_));
NAND_g _25234_ (.A(_09030_), .B(_04451_), .Y(_04452_));
AND_g _25235_ (.A(_04448_), .B(_04452_), .Y(_04453_));
NAND_g _25236_ (.A(_00008_[1]), .B(_04444_), .Y(_04454_));
NAND_g _25237_ (.A(_09031_), .B(_04453_), .Y(_04455_));
AND_g _25238_ (.A(_04454_), .B(_04455_), .Y(_04456_));
NAND_g _25239_ (.A(_09033_), .B(_04456_), .Y(_04457_));
NAND_g _25240_ (.A(cpuregs[13][12]), .B(_00008_[0]), .Y(_04458_));
NAND_g _25241_ (.A(cpuregs[12][12]), .B(_09030_), .Y(_04459_));
AND_g _25242_ (.A(_00008_[2]), .B(_04459_), .Y(_04460_));
NAND_g _25243_ (.A(_04458_), .B(_04460_), .Y(_04461_));
NAND_g _25244_ (.A(cpuregs[9][12]), .B(_00008_[0]), .Y(_04462_));
NAND_g _25245_ (.A(cpuregs[8][12]), .B(_09030_), .Y(_04463_));
AND_g _25246_ (.A(_09032_), .B(_04463_), .Y(_04464_));
NAND_g _25247_ (.A(_04462_), .B(_04464_), .Y(_04465_));
AND_g _25248_ (.A(_09031_), .B(_04465_), .Y(_04466_));
NAND_g _25249_ (.A(_04461_), .B(_04466_), .Y(_04467_));
NAND_g _25250_ (.A(cpuregs[15][12]), .B(_00008_[0]), .Y(_04468_));
NAND_g _25251_ (.A(cpuregs[14][12]), .B(_09030_), .Y(_04469_));
AND_g _25252_ (.A(_00008_[2]), .B(_04469_), .Y(_04470_));
NAND_g _25253_ (.A(_04468_), .B(_04470_), .Y(_04471_));
NAND_g _25254_ (.A(cpuregs[11][12]), .B(_00008_[0]), .Y(_04472_));
NAND_g _25255_ (.A(cpuregs[10][12]), .B(_09030_), .Y(_04473_));
AND_g _25256_ (.A(_09032_), .B(_04473_), .Y(_04474_));
NAND_g _25257_ (.A(_04472_), .B(_04474_), .Y(_04475_));
AND_g _25258_ (.A(_00008_[1]), .B(_04475_), .Y(_04476_));
NAND_g _25259_ (.A(_04471_), .B(_04476_), .Y(_04477_));
NAND_g _25260_ (.A(_04467_), .B(_04477_), .Y(_04478_));
AND_g _25261_ (.A(_00008_[3]), .B(_04478_), .Y(_04479_));
NOR_g _25262_ (.A(_00008_[4]), .B(_04479_), .Y(_04480_));
NAND_g _25263_ (.A(_04457_), .B(_04480_), .Y(_04481_));
NAND_g _25264_ (.A(cpuregs[25][12]), .B(_09032_), .Y(_04482_));
NAND_g _25265_ (.A(cpuregs[29][12]), .B(_00008_[2]), .Y(_04483_));
AND_g _25266_ (.A(_09031_), .B(_04483_), .Y(_04484_));
NAND_g _25267_ (.A(_04482_), .B(_04484_), .Y(_04485_));
NAND_g _25268_ (.A(cpuregs[31][12]), .B(_00008_[2]), .Y(_04486_));
NAND_g _25269_ (.A(cpuregs[27][12]), .B(_09032_), .Y(_04487_));
AND_g _25270_ (.A(_00008_[1]), .B(_04487_), .Y(_04488_));
NAND_g _25271_ (.A(_04486_), .B(_04488_), .Y(_04489_));
NAND_g _25272_ (.A(_04485_), .B(_04489_), .Y(_04490_));
NAND_g _25273_ (.A(_00008_[0]), .B(_04490_), .Y(_04491_));
NAND_g _25274_ (.A(cpuregs[24][12]), .B(_09032_), .Y(_04492_));
NAND_g _25275_ (.A(cpuregs[28][12]), .B(_00008_[2]), .Y(_04493_));
AND_g _25276_ (.A(_09031_), .B(_04493_), .Y(_04494_));
NAND_g _25277_ (.A(_04492_), .B(_04494_), .Y(_04495_));
NAND_g _25278_ (.A(cpuregs[26][12]), .B(_09032_), .Y(_04496_));
NAND_g _25279_ (.A(cpuregs[30][12]), .B(_00008_[2]), .Y(_04497_));
AND_g _25280_ (.A(_00008_[1]), .B(_04497_), .Y(_04498_));
NAND_g _25281_ (.A(_04496_), .B(_04498_), .Y(_04499_));
NAND_g _25282_ (.A(_04495_), .B(_04499_), .Y(_04500_));
NAND_g _25283_ (.A(_09030_), .B(_04500_), .Y(_04501_));
NAND_g _25284_ (.A(_04491_), .B(_04501_), .Y(_04502_));
NAND_g _25285_ (.A(_00008_[3]), .B(_04502_), .Y(_04503_));
NAND_g _25286_ (.A(cpuregs[17][12]), .B(_09031_), .Y(_04504_));
NAND_g _25287_ (.A(cpuregs[19][12]), .B(_00008_[1]), .Y(_04505_));
AND_g _25288_ (.A(_09032_), .B(_04505_), .Y(_04506_));
NAND_g _25289_ (.A(_04504_), .B(_04506_), .Y(_04507_));
NAND_g _25290_ (.A(cpuregs[21][12]), .B(_09031_), .Y(_04508_));
NAND_g _25291_ (.A(cpuregs[23][12]), .B(_00008_[1]), .Y(_04509_));
AND_g _25292_ (.A(_00008_[2]), .B(_04509_), .Y(_04510_));
NAND_g _25293_ (.A(_04508_), .B(_04510_), .Y(_04511_));
NAND_g _25294_ (.A(_04507_), .B(_04511_), .Y(_04512_));
NAND_g _25295_ (.A(_00008_[0]), .B(_04512_), .Y(_04513_));
NAND_g _25296_ (.A(cpuregs[16][12]), .B(_09031_), .Y(_04514_));
NAND_g _25297_ (.A(cpuregs[18][12]), .B(_00008_[1]), .Y(_04515_));
AND_g _25298_ (.A(_09032_), .B(_04515_), .Y(_04516_));
NAND_g _25299_ (.A(_04514_), .B(_04516_), .Y(_04517_));
NAND_g _25300_ (.A(cpuregs[20][12]), .B(_09031_), .Y(_04518_));
NAND_g _25301_ (.A(cpuregs[22][12]), .B(_00008_[1]), .Y(_04519_));
AND_g _25302_ (.A(_00008_[2]), .B(_04519_), .Y(_04520_));
NAND_g _25303_ (.A(_04518_), .B(_04520_), .Y(_04521_));
NAND_g _25304_ (.A(_04517_), .B(_04521_), .Y(_04522_));
NAND_g _25305_ (.A(_09030_), .B(_04522_), .Y(_04523_));
NAND_g _25306_ (.A(_04513_), .B(_04523_), .Y(_04524_));
AND_g _25307_ (.A(_09033_), .B(_04524_), .Y(_04525_));
NOT_g _25308_ (.A(_04525_), .Y(_04526_));
NAND_g _25309_ (.A(_04503_), .B(_04526_), .Y(_04527_));
NAND_g _25310_ (.A(_00008_[4]), .B(_04527_), .Y(_04528_));
AND_g _25311_ (.A(_14624_), .B(_04528_), .Y(_04529_));
NAND_g _25312_ (.A(_04481_), .B(_04529_), .Y(_04530_));
NAND_g _25313_ (.A(_04435_), .B(_04530_), .Y(_04531_));
NAND_g _25314_ (.A(_10595_), .B(_04531_), .Y(_04532_));
NAND_g _25315_ (.A(pcpi_rs1[11]), .B(_14481_), .Y(_04533_));
AND_g _25316_ (.A(_04197_), .B(_04533_), .Y(_04534_));
NAND_g _25317_ (.A(_13879_), .B(_04534_), .Y(_04535_));
NAND_g _25318_ (.A(pcpi_rs1[16]), .B(_14482_), .Y(_04536_));
AND_g _25319_ (.A(_04194_), .B(_04536_), .Y(_04537_));
NAND_g _25320_ (.A(_13880_), .B(_04537_), .Y(_04538_));
AND_g _25321_ (.A(_04535_), .B(_04538_), .Y(_04539_));
NAND_g _25322_ (.A(_13883_), .B(_04539_), .Y(_04540_));
AND_g _25323_ (.A(_14488_), .B(_04532_), .Y(_04541_));
AND_g _25324_ (.A(_04540_), .B(_04541_), .Y(_04542_));
AND_g _25325_ (.A(_04434_), .B(_04542_), .Y(_04543_));
NOR_g _25326_ (.A(_04432_), .B(_04543_), .Y(_01030_));
NOR_g _25327_ (.A(pcpi_rs1[13]), .B(_14488_), .Y(_04544_));
XOR_g _25328_ (.A(decoded_imm[13]), .B(pcpi_rs1[13]), .Y(_04545_));
XNOR_g _25329_ (.A(_14576_), .B(_04545_), .Y(_04546_));
NAND_g _25330_ (.A(_14614_), .B(_04546_), .Y(_04547_));
NAND_g _25331_ (.A(reg_pc[13]), .B(_14617_), .Y(_04548_));
NAND_g _25332_ (.A(cpuregs[9][13]), .B(_09032_), .Y(_04549_));
NAND_g _25333_ (.A(cpuregs[13][13]), .B(_00008_[2]), .Y(_04550_));
NAND_g _25334_ (.A(_04549_), .B(_04550_), .Y(_04551_));
NAND_g _25335_ (.A(_00008_[0]), .B(_04551_), .Y(_04552_));
NAND_g _25336_ (.A(cpuregs[12][13]), .B(_00008_[2]), .Y(_04553_));
NAND_g _25337_ (.A(cpuregs[8][13]), .B(_09032_), .Y(_04554_));
NAND_g _25338_ (.A(_04553_), .B(_04554_), .Y(_04555_));
NAND_g _25339_ (.A(_09030_), .B(_04555_), .Y(_04556_));
NAND_g _25340_ (.A(_04552_), .B(_04556_), .Y(_04557_));
NAND_g _25341_ (.A(_00008_[3]), .B(_04557_), .Y(_04558_));
NAND_g _25342_ (.A(cpuregs[5][13]), .B(_00008_[2]), .Y(_04559_));
NAND_g _25343_ (.A(cpuregs[1][13]), .B(_09032_), .Y(_04560_));
AND_g _25344_ (.A(_04559_), .B(_04560_), .Y(_04561_));
NAND_g _25345_ (.A(cpuregs[4][13]), .B(_00008_[2]), .Y(_04562_));
NAND_g _25346_ (.A(cpuregs[0][13]), .B(_09032_), .Y(_04563_));
AND_g _25347_ (.A(_04562_), .B(_04563_), .Y(_04564_));
NAND_g _25348_ (.A(_00008_[0]), .B(_04561_), .Y(_04565_));
NAND_g _25349_ (.A(_09030_), .B(_04564_), .Y(_04566_));
AND_g _25350_ (.A(_04565_), .B(_04566_), .Y(_04567_));
NAND_g _25351_ (.A(_09033_), .B(_04567_), .Y(_04568_));
NAND_g _25352_ (.A(_04558_), .B(_04568_), .Y(_04569_));
AND_g _25353_ (.A(_09031_), .B(_04569_), .Y(_04570_));
NAND_g _25354_ (.A(cpuregs[7][13]), .B(_00008_[0]), .Y(_04571_));
NAND_g _25355_ (.A(cpuregs[6][13]), .B(_09030_), .Y(_04572_));
AND_g _25356_ (.A(_00008_[2]), .B(_04572_), .Y(_04573_));
NAND_g _25357_ (.A(_04571_), .B(_04573_), .Y(_04574_));
NAND_g _25358_ (.A(cpuregs[3][13]), .B(_00008_[0]), .Y(_04575_));
NAND_g _25359_ (.A(cpuregs[2][13]), .B(_09030_), .Y(_04576_));
AND_g _25360_ (.A(_09032_), .B(_04576_), .Y(_04577_));
NAND_g _25361_ (.A(_04575_), .B(_04577_), .Y(_04578_));
AND_g _25362_ (.A(_09033_), .B(_04578_), .Y(_04579_));
NAND_g _25363_ (.A(_04574_), .B(_04579_), .Y(_04580_));
NAND_g _25364_ (.A(cpuregs[15][13]), .B(_00008_[0]), .Y(_04581_));
NAND_g _25365_ (.A(cpuregs[14][13]), .B(_09030_), .Y(_04582_));
AND_g _25366_ (.A(_00008_[2]), .B(_04582_), .Y(_04583_));
NAND_g _25367_ (.A(_04581_), .B(_04583_), .Y(_04584_));
NAND_g _25368_ (.A(cpuregs[11][13]), .B(_00008_[0]), .Y(_04585_));
NAND_g _25369_ (.A(cpuregs[10][13]), .B(_09030_), .Y(_04586_));
AND_g _25370_ (.A(_09032_), .B(_04586_), .Y(_04587_));
NAND_g _25371_ (.A(_04585_), .B(_04587_), .Y(_04588_));
AND_g _25372_ (.A(_00008_[3]), .B(_04588_), .Y(_04589_));
NAND_g _25373_ (.A(_04584_), .B(_04589_), .Y(_04590_));
NAND_g _25374_ (.A(_04580_), .B(_04590_), .Y(_04591_));
NAND_g _25375_ (.A(_00008_[1]), .B(_04591_), .Y(_04592_));
NOR_g _25376_ (.A(_00008_[4]), .B(_04570_), .Y(_04593_));
NAND_g _25377_ (.A(_04592_), .B(_04593_), .Y(_04594_));
NAND_g _25378_ (.A(cpuregs[26][13]), .B(_09032_), .Y(_04595_));
NAND_g _25379_ (.A(cpuregs[30][13]), .B(_00008_[2]), .Y(_04596_));
AND_g _25380_ (.A(_09030_), .B(_04596_), .Y(_04597_));
NAND_g _25381_ (.A(_04595_), .B(_04597_), .Y(_04598_));
NAND_g _25382_ (.A(cpuregs[31][13]), .B(_00008_[2]), .Y(_04599_));
NAND_g _25383_ (.A(cpuregs[27][13]), .B(_09032_), .Y(_04600_));
AND_g _25384_ (.A(_00008_[0]), .B(_04600_), .Y(_04601_));
NAND_g _25385_ (.A(_04599_), .B(_04601_), .Y(_04602_));
NAND_g _25386_ (.A(_04598_), .B(_04602_), .Y(_04603_));
NAND_g _25387_ (.A(_00008_[3]), .B(_04603_), .Y(_04604_));
NAND_g _25388_ (.A(cpuregs[18][13]), .B(_09032_), .Y(_04605_));
NAND_g _25389_ (.A(cpuregs[22][13]), .B(_00008_[2]), .Y(_04606_));
AND_g _25390_ (.A(_09030_), .B(_04606_), .Y(_04607_));
NAND_g _25391_ (.A(_04605_), .B(_04607_), .Y(_04608_));
NAND_g _25392_ (.A(cpuregs[19][13]), .B(_09032_), .Y(_04609_));
NAND_g _25393_ (.A(cpuregs[23][13]), .B(_00008_[2]), .Y(_04610_));
AND_g _25394_ (.A(_00008_[0]), .B(_04610_), .Y(_04611_));
NAND_g _25395_ (.A(_04609_), .B(_04611_), .Y(_04612_));
NAND_g _25396_ (.A(_04608_), .B(_04612_), .Y(_04613_));
NAND_g _25397_ (.A(_09033_), .B(_04613_), .Y(_04614_));
AND_g _25398_ (.A(_04604_), .B(_04614_), .Y(_04615_));
NAND_g _25399_ (.A(cpuregs[24][13]), .B(_09032_), .Y(_04616_));
NAND_g _25400_ (.A(cpuregs[28][13]), .B(_00008_[2]), .Y(_04617_));
AND_g _25401_ (.A(_09030_), .B(_04617_), .Y(_04618_));
NAND_g _25402_ (.A(_04616_), .B(_04618_), .Y(_04619_));
NAND_g _25403_ (.A(cpuregs[29][13]), .B(_00008_[2]), .Y(_04620_));
NAND_g _25404_ (.A(cpuregs[25][13]), .B(_09032_), .Y(_04621_));
AND_g _25405_ (.A(_00008_[0]), .B(_04621_), .Y(_04622_));
NAND_g _25406_ (.A(_04620_), .B(_04622_), .Y(_04623_));
NAND_g _25407_ (.A(_04619_), .B(_04623_), .Y(_04624_));
NAND_g _25408_ (.A(_00008_[3]), .B(_04624_), .Y(_04625_));
NAND_g _25409_ (.A(cpuregs[16][13]), .B(_09032_), .Y(_04626_));
NAND_g _25410_ (.A(cpuregs[20][13]), .B(_00008_[2]), .Y(_04627_));
AND_g _25411_ (.A(_09030_), .B(_04627_), .Y(_04628_));
NAND_g _25412_ (.A(_04626_), .B(_04628_), .Y(_04629_));
NAND_g _25413_ (.A(cpuregs[17][13]), .B(_09032_), .Y(_04630_));
NAND_g _25414_ (.A(cpuregs[21][13]), .B(_00008_[2]), .Y(_04631_));
AND_g _25415_ (.A(_00008_[0]), .B(_04631_), .Y(_04632_));
NAND_g _25416_ (.A(_04630_), .B(_04632_), .Y(_04633_));
NAND_g _25417_ (.A(_04629_), .B(_04633_), .Y(_04634_));
NAND_g _25418_ (.A(_09033_), .B(_04634_), .Y(_04635_));
AND_g _25419_ (.A(_04625_), .B(_04635_), .Y(_04636_));
NAND_g _25420_ (.A(_00008_[1]), .B(_04615_), .Y(_04637_));
NAND_g _25421_ (.A(_09031_), .B(_04636_), .Y(_04638_));
AND_g _25422_ (.A(_00008_[4]), .B(_04637_), .Y(_04639_));
NAND_g _25423_ (.A(_04638_), .B(_04639_), .Y(_04640_));
AND_g _25424_ (.A(_14624_), .B(_04640_), .Y(_04641_));
NAND_g _25425_ (.A(_04594_), .B(_04641_), .Y(_04642_));
NAND_g _25426_ (.A(_04548_), .B(_04642_), .Y(_04643_));
NAND_g _25427_ (.A(_10595_), .B(_04643_), .Y(_04644_));
NAND_g _25428_ (.A(pcpi_rs1[12]), .B(_14481_), .Y(_04645_));
AND_g _25429_ (.A(_04312_), .B(_04645_), .Y(_04646_));
NAND_g _25430_ (.A(pcpi_rs1[17]), .B(_14482_), .Y(_04647_));
AND_g _25431_ (.A(_04309_), .B(_04647_), .Y(_04648_));
NAND_g _25432_ (.A(_13880_), .B(_04648_), .Y(_04649_));
NAND_g _25433_ (.A(_13879_), .B(_04646_), .Y(_04650_));
AND_g _25434_ (.A(_13883_), .B(_04649_), .Y(_04651_));
NAND_g _25435_ (.A(_04650_), .B(_04651_), .Y(_04652_));
AND_g _25436_ (.A(_14488_), .B(_04652_), .Y(_04653_));
AND_g _25437_ (.A(_04644_), .B(_04653_), .Y(_04654_));
AND_g _25438_ (.A(_04547_), .B(_04654_), .Y(_04655_));
NOR_g _25439_ (.A(_04544_), .B(_04655_), .Y(_01031_));
NOR_g _25440_ (.A(pcpi_rs1[14]), .B(_14488_), .Y(_04656_));
XOR_g _25441_ (.A(_14524_), .B(_14578_), .Y(_04657_));
NAND_g _25442_ (.A(_14614_), .B(_04657_), .Y(_04658_));
NAND_g _25443_ (.A(reg_pc[14]), .B(_14617_), .Y(_04659_));
NAND_g _25444_ (.A(_08969_), .B(_00008_[2]), .Y(_04660_));
NOR_g _25445_ (.A(cpuregs[3][14]), .B(_00008_[2]), .Y(_04661_));
NOR_g _25446_ (.A(_09030_), .B(_04661_), .Y(_04662_));
NAND_g _25447_ (.A(_04660_), .B(_04662_), .Y(_04663_));
NOR_g _25448_ (.A(cpuregs[2][14]), .B(_00008_[2]), .Y(_04664_));
AND_g _25449_ (.A(_09009_), .B(_00008_[2]), .Y(_04665_));
NOR_g _25450_ (.A(_04664_), .B(_04665_), .Y(_04666_));
NAND_g _25451_ (.A(_09030_), .B(_04666_), .Y(_04667_));
NAND_g _25452_ (.A(_04663_), .B(_04667_), .Y(_04668_));
NAND_g _25453_ (.A(_00008_[1]), .B(_04668_), .Y(_04669_));
NAND_g _25454_ (.A(_08952_), .B(_00008_[2]), .Y(_04670_));
NOR_g _25455_ (.A(cpuregs[1][14]), .B(_00008_[2]), .Y(_04671_));
NOR_g _25456_ (.A(_09030_), .B(_04671_), .Y(_04672_));
NAND_g _25457_ (.A(_04670_), .B(_04672_), .Y(_04673_));
NOR_g _25458_ (.A(cpuregs[0][14]), .B(_00008_[2]), .Y(_04674_));
AND_g _25459_ (.A(_08910_), .B(_00008_[2]), .Y(_04675_));
NOR_g _25460_ (.A(_04674_), .B(_04675_), .Y(_04676_));
NAND_g _25461_ (.A(_09030_), .B(_04676_), .Y(_04677_));
NAND_g _25462_ (.A(_04673_), .B(_04677_), .Y(_04678_));
NAND_g _25463_ (.A(_09031_), .B(_04678_), .Y(_04679_));
NAND_g _25464_ (.A(_04669_), .B(_04679_), .Y(_04680_));
NAND_g _25465_ (.A(_09033_), .B(_04680_), .Y(_04681_));
NAND_g _25466_ (.A(cpuregs[13][14]), .B(_00008_[0]), .Y(_04682_));
NAND_g _25467_ (.A(cpuregs[12][14]), .B(_09030_), .Y(_04683_));
AND_g _25468_ (.A(_00008_[2]), .B(_04683_), .Y(_04684_));
NAND_g _25469_ (.A(_04682_), .B(_04684_), .Y(_04685_));
NAND_g _25470_ (.A(cpuregs[9][14]), .B(_00008_[0]), .Y(_04686_));
NAND_g _25471_ (.A(cpuregs[8][14]), .B(_09030_), .Y(_04687_));
AND_g _25472_ (.A(_09032_), .B(_04687_), .Y(_04688_));
NAND_g _25473_ (.A(_04686_), .B(_04688_), .Y(_04689_));
AND_g _25474_ (.A(_09031_), .B(_04689_), .Y(_04690_));
NAND_g _25475_ (.A(_04685_), .B(_04690_), .Y(_04691_));
NAND_g _25476_ (.A(cpuregs[15][14]), .B(_00008_[0]), .Y(_04692_));
NAND_g _25477_ (.A(cpuregs[14][14]), .B(_09030_), .Y(_04693_));
AND_g _25478_ (.A(_00008_[2]), .B(_04693_), .Y(_04694_));
NAND_g _25479_ (.A(_04692_), .B(_04694_), .Y(_04695_));
NAND_g _25480_ (.A(cpuregs[11][14]), .B(_00008_[0]), .Y(_04696_));
NAND_g _25481_ (.A(cpuregs[10][14]), .B(_09030_), .Y(_04697_));
AND_g _25482_ (.A(_09032_), .B(_04697_), .Y(_04698_));
NAND_g _25483_ (.A(_04696_), .B(_04698_), .Y(_04699_));
AND_g _25484_ (.A(_00008_[1]), .B(_04699_), .Y(_04700_));
NAND_g _25485_ (.A(_04695_), .B(_04700_), .Y(_04701_));
NAND_g _25486_ (.A(_04691_), .B(_04701_), .Y(_04702_));
AND_g _25487_ (.A(_00008_[3]), .B(_04702_), .Y(_04703_));
NOR_g _25488_ (.A(_00008_[4]), .B(_04703_), .Y(_04704_));
NAND_g _25489_ (.A(_04681_), .B(_04704_), .Y(_04705_));
NAND_g _25490_ (.A(cpuregs[25][14]), .B(_09032_), .Y(_04706_));
NAND_g _25491_ (.A(cpuregs[29][14]), .B(_00008_[2]), .Y(_04707_));
AND_g _25492_ (.A(_09031_), .B(_04707_), .Y(_04708_));
NAND_g _25493_ (.A(_04706_), .B(_04708_), .Y(_04709_));
NAND_g _25494_ (.A(cpuregs[31][14]), .B(_00008_[2]), .Y(_04710_));
NAND_g _25495_ (.A(cpuregs[27][14]), .B(_09032_), .Y(_04711_));
AND_g _25496_ (.A(_00008_[1]), .B(_04711_), .Y(_04712_));
NAND_g _25497_ (.A(_04710_), .B(_04712_), .Y(_04713_));
NAND_g _25498_ (.A(_04709_), .B(_04713_), .Y(_04714_));
NAND_g _25499_ (.A(_00008_[0]), .B(_04714_), .Y(_04715_));
NAND_g _25500_ (.A(cpuregs[24][14]), .B(_09032_), .Y(_04716_));
NAND_g _25501_ (.A(cpuregs[28][14]), .B(_00008_[2]), .Y(_04717_));
AND_g _25502_ (.A(_09031_), .B(_04717_), .Y(_04718_));
NAND_g _25503_ (.A(_04716_), .B(_04718_), .Y(_04719_));
NAND_g _25504_ (.A(cpuregs[26][14]), .B(_09032_), .Y(_04720_));
NAND_g _25505_ (.A(cpuregs[30][14]), .B(_00008_[2]), .Y(_04721_));
AND_g _25506_ (.A(_00008_[1]), .B(_04721_), .Y(_04722_));
NAND_g _25507_ (.A(_04720_), .B(_04722_), .Y(_04723_));
NAND_g _25508_ (.A(_04719_), .B(_04723_), .Y(_04724_));
NAND_g _25509_ (.A(_09030_), .B(_04724_), .Y(_04725_));
NAND_g _25510_ (.A(_04715_), .B(_04725_), .Y(_04726_));
NAND_g _25511_ (.A(_00008_[3]), .B(_04726_), .Y(_04727_));
NAND_g _25512_ (.A(cpuregs[17][14]), .B(_09031_), .Y(_04728_));
NAND_g _25513_ (.A(cpuregs[19][14]), .B(_00008_[1]), .Y(_04729_));
AND_g _25514_ (.A(_09032_), .B(_04729_), .Y(_04730_));
NAND_g _25515_ (.A(_04728_), .B(_04730_), .Y(_04731_));
NAND_g _25516_ (.A(cpuregs[21][14]), .B(_09031_), .Y(_04732_));
NAND_g _25517_ (.A(cpuregs[23][14]), .B(_00008_[1]), .Y(_04733_));
AND_g _25518_ (.A(_00008_[2]), .B(_04733_), .Y(_04734_));
NAND_g _25519_ (.A(_04732_), .B(_04734_), .Y(_04735_));
NAND_g _25520_ (.A(_04731_), .B(_04735_), .Y(_04736_));
NAND_g _25521_ (.A(_00008_[0]), .B(_04736_), .Y(_04737_));
NAND_g _25522_ (.A(cpuregs[16][14]), .B(_09031_), .Y(_04738_));
NAND_g _25523_ (.A(cpuregs[18][14]), .B(_00008_[1]), .Y(_04739_));
AND_g _25524_ (.A(_09032_), .B(_04739_), .Y(_04740_));
NAND_g _25525_ (.A(_04738_), .B(_04740_), .Y(_04741_));
NAND_g _25526_ (.A(cpuregs[20][14]), .B(_09031_), .Y(_04742_));
NAND_g _25527_ (.A(cpuregs[22][14]), .B(_00008_[1]), .Y(_04743_));
AND_g _25528_ (.A(_00008_[2]), .B(_04743_), .Y(_04744_));
NAND_g _25529_ (.A(_04742_), .B(_04744_), .Y(_04745_));
NAND_g _25530_ (.A(_04741_), .B(_04745_), .Y(_04746_));
NAND_g _25531_ (.A(_09030_), .B(_04746_), .Y(_04747_));
NAND_g _25532_ (.A(_04737_), .B(_04747_), .Y(_04748_));
AND_g _25533_ (.A(_09033_), .B(_04748_), .Y(_04749_));
NOT_g _25534_ (.A(_04749_), .Y(_04750_));
NAND_g _25535_ (.A(_04727_), .B(_04750_), .Y(_04751_));
NAND_g _25536_ (.A(_00008_[4]), .B(_04751_), .Y(_04752_));
AND_g _25537_ (.A(_14624_), .B(_04752_), .Y(_04753_));
NAND_g _25538_ (.A(_04705_), .B(_04753_), .Y(_04754_));
NAND_g _25539_ (.A(_04659_), .B(_04754_), .Y(_04755_));
NAND_g _25540_ (.A(_10595_), .B(_04755_), .Y(_04756_));
NAND_g _25541_ (.A(pcpi_rs1[13]), .B(_14481_), .Y(_04757_));
AND_g _25542_ (.A(_04423_), .B(_04757_), .Y(_04758_));
NAND_g _25543_ (.A(_13879_), .B(_04758_), .Y(_04759_));
NAND_g _25544_ (.A(pcpi_rs1[18]), .B(_14482_), .Y(_04760_));
AND_g _25545_ (.A(_04421_), .B(_04760_), .Y(_04761_));
NAND_g _25546_ (.A(_13880_), .B(_04761_), .Y(_04762_));
AND_g _25547_ (.A(_04759_), .B(_04762_), .Y(_04763_));
NAND_g _25548_ (.A(_13883_), .B(_04763_), .Y(_04764_));
AND_g _25549_ (.A(_14488_), .B(_04756_), .Y(_04765_));
AND_g _25550_ (.A(_04764_), .B(_04765_), .Y(_04766_));
AND_g _25551_ (.A(_04658_), .B(_04766_), .Y(_04767_));
NOR_g _25552_ (.A(_04656_), .B(_04767_), .Y(_01032_));
NOR_g _25553_ (.A(pcpi_rs1[15]), .B(_14488_), .Y(_04768_));
XOR_g _25554_ (.A(decoded_imm[15]), .B(pcpi_rs1[15]), .Y(_04769_));
XNOR_g _25555_ (.A(_14580_), .B(_04769_), .Y(_04770_));
NAND_g _25556_ (.A(_14614_), .B(_04770_), .Y(_04771_));
NAND_g _25557_ (.A(reg_pc[15]), .B(_14617_), .Y(_04772_));
NAND_g _25558_ (.A(cpuregs[13][15]), .B(_00008_[2]), .Y(_04773_));
NAND_g _25559_ (.A(cpuregs[9][15]), .B(_09032_), .Y(_04774_));
NAND_g _25560_ (.A(_04773_), .B(_04774_), .Y(_04775_));
NAND_g _25561_ (.A(_00008_[0]), .B(_04775_), .Y(_04776_));
NAND_g _25562_ (.A(cpuregs[12][15]), .B(_00008_[2]), .Y(_04777_));
NAND_g _25563_ (.A(cpuregs[8][15]), .B(_09032_), .Y(_04778_));
AND_g _25564_ (.A(_04777_), .B(_04778_), .Y(_04779_));
NOR_g _25565_ (.A(_00008_[0]), .B(_04779_), .Y(_04780_));
NAND_g _25566_ (.A(_08911_), .B(_00008_[2]), .Y(_04781_));
NOR_g _25567_ (.A(cpuregs[0][15]), .B(_00008_[2]), .Y(_04782_));
NOR_g _25568_ (.A(_00008_[0]), .B(_04782_), .Y(_04783_));
NAND_g _25569_ (.A(_04781_), .B(_04783_), .Y(_04784_));
NAND_g _25570_ (.A(_08953_), .B(_00008_[2]), .Y(_04785_));
NOR_g _25571_ (.A(cpuregs[1][15]), .B(_00008_[2]), .Y(_04786_));
NOR_g _25572_ (.A(_09030_), .B(_04786_), .Y(_04787_));
NAND_g _25573_ (.A(_04785_), .B(_04787_), .Y(_04788_));
NAND_g _25574_ (.A(cpuregs[11][15]), .B(_09032_), .Y(_04789_));
NAND_g _25575_ (.A(cpuregs[15][15]), .B(_00008_[2]), .Y(_04790_));
NAND_g _25576_ (.A(_04789_), .B(_04790_), .Y(_04791_));
AND_g _25577_ (.A(_00008_[0]), .B(_04791_), .Y(_04792_));
NAND_g _25578_ (.A(cpuregs[14][15]), .B(_00008_[2]), .Y(_04793_));
NAND_g _25579_ (.A(cpuregs[10][15]), .B(_09032_), .Y(_04794_));
AND_g _25580_ (.A(_04793_), .B(_04794_), .Y(_04795_));
NOR_g _25581_ (.A(_00008_[0]), .B(_04795_), .Y(_04796_));
NOR_g _25582_ (.A(_04792_), .B(_04796_), .Y(_04797_));
NAND_g _25583_ (.A(_09010_), .B(_00008_[2]), .Y(_04798_));
NOR_g _25584_ (.A(cpuregs[2][15]), .B(_00008_[2]), .Y(_04799_));
NOR_g _25585_ (.A(_00008_[0]), .B(_04799_), .Y(_04800_));
NAND_g _25586_ (.A(_04798_), .B(_04800_), .Y(_04801_));
NAND_g _25587_ (.A(_08970_), .B(_00008_[2]), .Y(_04802_));
NOR_g _25588_ (.A(cpuregs[3][15]), .B(_00008_[2]), .Y(_04803_));
NOR_g _25589_ (.A(_09030_), .B(_04803_), .Y(_04804_));
NAND_g _25590_ (.A(_04802_), .B(_04804_), .Y(_04805_));
AND_g _25591_ (.A(_04801_), .B(_04805_), .Y(_04806_));
AND_g _25592_ (.A(_09031_), .B(_04784_), .Y(_04807_));
NAND_g _25593_ (.A(_04788_), .B(_04807_), .Y(_04808_));
NAND_g _25594_ (.A(_00008_[1]), .B(_04806_), .Y(_04809_));
AND_g _25595_ (.A(_04808_), .B(_04809_), .Y(_04810_));
NAND_g _25596_ (.A(_09033_), .B(_04810_), .Y(_04811_));
NAND_g _25597_ (.A(_00008_[1]), .B(_04797_), .Y(_04812_));
NOR_g _25598_ (.A(_00008_[1]), .B(_04780_), .Y(_04813_));
NAND_g _25599_ (.A(_04776_), .B(_04813_), .Y(_04814_));
AND_g _25600_ (.A(_00008_[3]), .B(_04814_), .Y(_04815_));
AND_g _25601_ (.A(_04812_), .B(_04815_), .Y(_04816_));
NOR_g _25602_ (.A(_00008_[4]), .B(_04816_), .Y(_04817_));
NAND_g _25603_ (.A(_04811_), .B(_04817_), .Y(_04818_));
NAND_g _25604_ (.A(_08893_), .B(_00008_[2]), .Y(_04819_));
NOR_g _25605_ (.A(cpuregs[19][15]), .B(_00008_[2]), .Y(_04820_));
NOR_g _25606_ (.A(cpuregs[18][15]), .B(_00008_[2]), .Y(_04821_));
AND_g _25607_ (.A(_08922_), .B(_00008_[2]), .Y(_04822_));
NOR_g _25608_ (.A(_04821_), .B(_04822_), .Y(_04823_));
NOR_g _25609_ (.A(_09030_), .B(_04820_), .Y(_04824_));
NAND_g _25610_ (.A(_04819_), .B(_04824_), .Y(_04825_));
NAND_g _25611_ (.A(_09030_), .B(_04823_), .Y(_04826_));
AND_g _25612_ (.A(_04825_), .B(_04826_), .Y(_04827_));
NAND_g _25613_ (.A(_00008_[1]), .B(_04827_), .Y(_04828_));
NOR_g _25614_ (.A(cpuregs[17][15]), .B(_00008_[2]), .Y(_04829_));
NAND_g _25615_ (.A(_08992_), .B(_00008_[2]), .Y(_04830_));
NOR_g _25616_ (.A(cpuregs[16][15]), .B(_00008_[2]), .Y(_04831_));
AND_g _25617_ (.A(_08848_), .B(_00008_[2]), .Y(_04832_));
NOR_g _25618_ (.A(_04831_), .B(_04832_), .Y(_04833_));
NOR_g _25619_ (.A(_09030_), .B(_04829_), .Y(_04834_));
NAND_g _25620_ (.A(_04830_), .B(_04834_), .Y(_04835_));
NAND_g _25621_ (.A(_09030_), .B(_04833_), .Y(_04836_));
AND_g _25622_ (.A(_04835_), .B(_04836_), .Y(_04837_));
NAND_g _25623_ (.A(_09031_), .B(_04837_), .Y(_04838_));
NAND_g _25624_ (.A(_04828_), .B(_04838_), .Y(_04839_));
NAND_g _25625_ (.A(_09033_), .B(_04839_), .Y(_04840_));
NAND_g _25626_ (.A(cpuregs[25][15]), .B(_09031_), .Y(_04841_));
NAND_g _25627_ (.A(cpuregs[27][15]), .B(_00008_[1]), .Y(_04842_));
AND_g _25628_ (.A(_09032_), .B(_04842_), .Y(_04843_));
NAND_g _25629_ (.A(_04841_), .B(_04843_), .Y(_04844_));
NAND_g _25630_ (.A(cpuregs[29][15]), .B(_09031_), .Y(_04845_));
NAND_g _25631_ (.A(cpuregs[31][15]), .B(_00008_[1]), .Y(_04846_));
AND_g _25632_ (.A(_00008_[2]), .B(_04846_), .Y(_04847_));
NAND_g _25633_ (.A(_04845_), .B(_04847_), .Y(_04848_));
NAND_g _25634_ (.A(_04844_), .B(_04848_), .Y(_04849_));
NAND_g _25635_ (.A(_00008_[0]), .B(_04849_), .Y(_04850_));
NAND_g _25636_ (.A(cpuregs[24][15]), .B(_09031_), .Y(_04851_));
NAND_g _25637_ (.A(cpuregs[26][15]), .B(_00008_[1]), .Y(_04852_));
AND_g _25638_ (.A(_09032_), .B(_04852_), .Y(_04853_));
NAND_g _25639_ (.A(_04851_), .B(_04853_), .Y(_04854_));
NAND_g _25640_ (.A(cpuregs[28][15]), .B(_09031_), .Y(_04855_));
NAND_g _25641_ (.A(cpuregs[30][15]), .B(_00008_[1]), .Y(_04856_));
AND_g _25642_ (.A(_00008_[2]), .B(_04856_), .Y(_04857_));
NAND_g _25643_ (.A(_04855_), .B(_04857_), .Y(_04858_));
NAND_g _25644_ (.A(_04854_), .B(_04858_), .Y(_04859_));
NAND_g _25645_ (.A(_09030_), .B(_04859_), .Y(_04860_));
NAND_g _25646_ (.A(_04850_), .B(_04860_), .Y(_04861_));
NAND_g _25647_ (.A(_00008_[3]), .B(_04861_), .Y(_04862_));
NAND_g _25648_ (.A(_04840_), .B(_04862_), .Y(_04863_));
NAND_g _25649_ (.A(_00008_[4]), .B(_04863_), .Y(_04864_));
AND_g _25650_ (.A(_14624_), .B(_04818_), .Y(_04865_));
NAND_g _25651_ (.A(_04864_), .B(_04865_), .Y(_04866_));
NAND_g _25652_ (.A(_04772_), .B(_04866_), .Y(_04867_));
NAND_g _25653_ (.A(_10595_), .B(_04867_), .Y(_04868_));
NAND_g _25654_ (.A(pcpi_rs1[14]), .B(_14481_), .Y(_04869_));
AND_g _25655_ (.A(_04536_), .B(_04869_), .Y(_04870_));
NAND_g _25656_ (.A(pcpi_rs1[19]), .B(_14482_), .Y(_04871_));
AND_g _25657_ (.A(_04533_), .B(_04871_), .Y(_04872_));
NAND_g _25658_ (.A(_13880_), .B(_04872_), .Y(_04873_));
NAND_g _25659_ (.A(_13879_), .B(_04870_), .Y(_04874_));
AND_g _25660_ (.A(_13883_), .B(_04873_), .Y(_04875_));
NAND_g _25661_ (.A(_04874_), .B(_04875_), .Y(_04876_));
AND_g _25662_ (.A(_14488_), .B(_04876_), .Y(_04877_));
AND_g _25663_ (.A(_04868_), .B(_04877_), .Y(_04878_));
AND_g _25664_ (.A(_04771_), .B(_04878_), .Y(_04879_));
NOR_g _25665_ (.A(_04768_), .B(_04879_), .Y(_01033_));
NOR_g _25666_ (.A(pcpi_rs1[16]), .B(_14488_), .Y(_04880_));
NAND_g _25667_ (.A(reg_pc[16]), .B(_14617_), .Y(_04881_));
NAND_g _25668_ (.A(cpuregs[12][16]), .B(_00008_[2]), .Y(_04882_));
NAND_g _25669_ (.A(cpuregs[8][16]), .B(_09032_), .Y(_04883_));
NAND_g _25670_ (.A(_04882_), .B(_04883_), .Y(_04884_));
NAND_g _25671_ (.A(_09030_), .B(_04884_), .Y(_04885_));
NAND_g _25672_ (.A(cpuregs[13][16]), .B(_00008_[2]), .Y(_04886_));
NAND_g _25673_ (.A(cpuregs[9][16]), .B(_09032_), .Y(_04887_));
NAND_g _25674_ (.A(_04886_), .B(_04887_), .Y(_04888_));
NAND_g _25675_ (.A(_00008_[0]), .B(_04888_), .Y(_04889_));
NAND_g _25676_ (.A(_04885_), .B(_04889_), .Y(_04890_));
NAND_g _25677_ (.A(_00008_[3]), .B(_04890_), .Y(_04891_));
NAND_g _25678_ (.A(cpuregs[5][16]), .B(_00008_[2]), .Y(_04892_));
NAND_g _25679_ (.A(cpuregs[1][16]), .B(_09032_), .Y(_04893_));
NAND_g _25680_ (.A(_04892_), .B(_04893_), .Y(_04894_));
NAND_g _25681_ (.A(_00008_[0]), .B(_04894_), .Y(_04895_));
NAND_g _25682_ (.A(cpuregs[4][16]), .B(_00008_[2]), .Y(_04896_));
NAND_g _25683_ (.A(cpuregs[0][16]), .B(_09032_), .Y(_04897_));
NAND_g _25684_ (.A(_04896_), .B(_04897_), .Y(_04898_));
NAND_g _25685_ (.A(_09030_), .B(_04898_), .Y(_04899_));
NAND_g _25686_ (.A(_04895_), .B(_04899_), .Y(_04900_));
NAND_g _25687_ (.A(_09033_), .B(_04900_), .Y(_04901_));
NAND_g _25688_ (.A(_04891_), .B(_04901_), .Y(_04902_));
AND_g _25689_ (.A(_09031_), .B(_04902_), .Y(_04903_));
NAND_g _25690_ (.A(cpuregs[11][16]), .B(_09032_), .Y(_04904_));
NAND_g _25691_ (.A(cpuregs[15][16]), .B(_00008_[2]), .Y(_04905_));
NAND_g _25692_ (.A(_04904_), .B(_04905_), .Y(_04906_));
NAND_g _25693_ (.A(_00008_[0]), .B(_04906_), .Y(_04907_));
NAND_g _25694_ (.A(cpuregs[14][16]), .B(_00008_[2]), .Y(_04908_));
NAND_g _25695_ (.A(cpuregs[10][16]), .B(_09032_), .Y(_04909_));
NAND_g _25696_ (.A(_04908_), .B(_04909_), .Y(_04910_));
NAND_g _25697_ (.A(_09030_), .B(_04910_), .Y(_04911_));
NAND_g _25698_ (.A(_04907_), .B(_04911_), .Y(_04912_));
NAND_g _25699_ (.A(_00008_[3]), .B(_04912_), .Y(_04913_));
NAND_g _25700_ (.A(cpuregs[7][16]), .B(_00008_[2]), .Y(_04914_));
NAND_g _25701_ (.A(cpuregs[3][16]), .B(_09032_), .Y(_04915_));
AND_g _25702_ (.A(_04914_), .B(_04915_), .Y(_04916_));
NAND_g _25703_ (.A(cpuregs[6][16]), .B(_00008_[2]), .Y(_04917_));
NAND_g _25704_ (.A(cpuregs[2][16]), .B(_09032_), .Y(_04918_));
AND_g _25705_ (.A(_04917_), .B(_04918_), .Y(_04919_));
NAND_g _25706_ (.A(_00008_[0]), .B(_04916_), .Y(_04920_));
NAND_g _25707_ (.A(_09030_), .B(_04919_), .Y(_04921_));
AND_g _25708_ (.A(_04920_), .B(_04921_), .Y(_04922_));
NAND_g _25709_ (.A(_09033_), .B(_04922_), .Y(_04923_));
NAND_g _25710_ (.A(_04913_), .B(_04923_), .Y(_04924_));
NAND_g _25711_ (.A(_00008_[1]), .B(_04924_), .Y(_04925_));
NOR_g _25712_ (.A(_00008_[4]), .B(_04903_), .Y(_04926_));
NAND_g _25713_ (.A(_04925_), .B(_04926_), .Y(_04927_));
NAND_g _25714_ (.A(cpuregs[25][16]), .B(_09032_), .Y(_04928_));
NAND_g _25715_ (.A(cpuregs[29][16]), .B(_00008_[2]), .Y(_04929_));
AND_g _25716_ (.A(_09031_), .B(_04929_), .Y(_04930_));
NAND_g _25717_ (.A(_04928_), .B(_04930_), .Y(_04931_));
NAND_g _25718_ (.A(cpuregs[31][16]), .B(_00008_[2]), .Y(_04932_));
NAND_g _25719_ (.A(cpuregs[27][16]), .B(_09032_), .Y(_04933_));
AND_g _25720_ (.A(_00008_[1]), .B(_04933_), .Y(_04934_));
NAND_g _25721_ (.A(_04932_), .B(_04934_), .Y(_04935_));
NAND_g _25722_ (.A(_04931_), .B(_04935_), .Y(_04936_));
NAND_g _25723_ (.A(_00008_[0]), .B(_04936_), .Y(_04937_));
NAND_g _25724_ (.A(cpuregs[24][16]), .B(_09032_), .Y(_04938_));
NAND_g _25725_ (.A(cpuregs[28][16]), .B(_00008_[2]), .Y(_04939_));
AND_g _25726_ (.A(_09031_), .B(_04939_), .Y(_04940_));
NAND_g _25727_ (.A(_04938_), .B(_04940_), .Y(_04941_));
NAND_g _25728_ (.A(cpuregs[26][16]), .B(_09032_), .Y(_04942_));
NAND_g _25729_ (.A(cpuregs[30][16]), .B(_00008_[2]), .Y(_04943_));
AND_g _25730_ (.A(_00008_[1]), .B(_04943_), .Y(_04944_));
NAND_g _25731_ (.A(_04942_), .B(_04944_), .Y(_04945_));
NAND_g _25732_ (.A(_04941_), .B(_04945_), .Y(_04946_));
NAND_g _25733_ (.A(_09030_), .B(_04946_), .Y(_04947_));
NAND_g _25734_ (.A(_04937_), .B(_04947_), .Y(_04948_));
NAND_g _25735_ (.A(_00008_[3]), .B(_04948_), .Y(_04949_));
NAND_g _25736_ (.A(cpuregs[17][16]), .B(_09031_), .Y(_04950_));
NAND_g _25737_ (.A(cpuregs[19][16]), .B(_00008_[1]), .Y(_04951_));
AND_g _25738_ (.A(_09032_), .B(_04951_), .Y(_04952_));
NAND_g _25739_ (.A(_04950_), .B(_04952_), .Y(_04953_));
NAND_g _25740_ (.A(cpuregs[21][16]), .B(_09031_), .Y(_04954_));
NAND_g _25741_ (.A(cpuregs[23][16]), .B(_00008_[1]), .Y(_04955_));
AND_g _25742_ (.A(_00008_[2]), .B(_04955_), .Y(_04956_));
NAND_g _25743_ (.A(_04954_), .B(_04956_), .Y(_04957_));
NAND_g _25744_ (.A(_04953_), .B(_04957_), .Y(_04958_));
NAND_g _25745_ (.A(_00008_[0]), .B(_04958_), .Y(_04959_));
NAND_g _25746_ (.A(cpuregs[16][16]), .B(_09031_), .Y(_04960_));
NAND_g _25747_ (.A(cpuregs[18][16]), .B(_00008_[1]), .Y(_04961_));
AND_g _25748_ (.A(_09032_), .B(_04961_), .Y(_04962_));
NAND_g _25749_ (.A(_04960_), .B(_04962_), .Y(_04963_));
NAND_g _25750_ (.A(cpuregs[20][16]), .B(_09031_), .Y(_04964_));
NAND_g _25751_ (.A(cpuregs[22][16]), .B(_00008_[1]), .Y(_04965_));
AND_g _25752_ (.A(_00008_[2]), .B(_04965_), .Y(_04966_));
NAND_g _25753_ (.A(_04964_), .B(_04966_), .Y(_04967_));
NAND_g _25754_ (.A(_04963_), .B(_04967_), .Y(_04968_));
NAND_g _25755_ (.A(_09030_), .B(_04968_), .Y(_04969_));
NAND_g _25756_ (.A(_04959_), .B(_04969_), .Y(_04970_));
AND_g _25757_ (.A(_09033_), .B(_04970_), .Y(_04971_));
NOT_g _25758_ (.A(_04971_), .Y(_04972_));
NAND_g _25759_ (.A(_04949_), .B(_04972_), .Y(_04973_));
NAND_g _25760_ (.A(_00008_[4]), .B(_04973_), .Y(_04974_));
AND_g _25761_ (.A(_14624_), .B(_04974_), .Y(_04975_));
NAND_g _25762_ (.A(_04927_), .B(_04975_), .Y(_04976_));
NAND_g _25763_ (.A(_04881_), .B(_04976_), .Y(_04977_));
NAND_g _25764_ (.A(_10595_), .B(_04977_), .Y(_04978_));
NAND_g _25765_ (.A(pcpi_rs1[15]), .B(_14481_), .Y(_04979_));
AND_g _25766_ (.A(_04647_), .B(_04979_), .Y(_04980_));
NAND_g _25767_ (.A(pcpi_rs1[20]), .B(_14482_), .Y(_04981_));
AND_g _25768_ (.A(_04645_), .B(_04981_), .Y(_04982_));
NAND_g _25769_ (.A(_13879_), .B(_04980_), .Y(_04983_));
NAND_g _25770_ (.A(_13880_), .B(_04982_), .Y(_04984_));
AND_g _25771_ (.A(_13883_), .B(_04983_), .Y(_04985_));
NAND_g _25772_ (.A(_04984_), .B(_04985_), .Y(_04986_));
AND_g _25773_ (.A(_14488_), .B(_04986_), .Y(_04987_));
AND_g _25774_ (.A(_04978_), .B(_04987_), .Y(_04988_));
XOR_g _25775_ (.A(_14520_), .B(_14582_), .Y(_04989_));
NAND_g _25776_ (.A(_14614_), .B(_04989_), .Y(_04990_));
AND_g _25777_ (.A(_04988_), .B(_04990_), .Y(_04991_));
NOR_g _25778_ (.A(_04880_), .B(_04991_), .Y(_01034_));
NOR_g _25779_ (.A(pcpi_rs1[17]), .B(_14488_), .Y(_04992_));
NAND_g _25780_ (.A(reg_pc[17]), .B(_14617_), .Y(_04993_));
NAND_g _25781_ (.A(cpuregs[7][17]), .B(_00008_[2]), .Y(_04994_));
NAND_g _25782_ (.A(cpuregs[3][17]), .B(_09032_), .Y(_04995_));
NAND_g _25783_ (.A(_04994_), .B(_04995_), .Y(_04996_));
AND_g _25784_ (.A(_00008_[0]), .B(_04996_), .Y(_04997_));
NAND_g _25785_ (.A(cpuregs[6][17]), .B(_00008_[2]), .Y(_04998_));
NAND_g _25786_ (.A(cpuregs[2][17]), .B(_09032_), .Y(_04999_));
AND_g _25787_ (.A(_04998_), .B(_04999_), .Y(_05000_));
NOR_g _25788_ (.A(_00008_[0]), .B(_05000_), .Y(_05001_));
NOR_g _25789_ (.A(_04997_), .B(_05001_), .Y(_05002_));
NAND_g _25790_ (.A(cpuregs[5][17]), .B(_00008_[2]), .Y(_05003_));
NAND_g _25791_ (.A(cpuregs[1][17]), .B(_09032_), .Y(_05004_));
NAND_g _25792_ (.A(_05003_), .B(_05004_), .Y(_05005_));
NAND_g _25793_ (.A(_00008_[0]), .B(_05005_), .Y(_05006_));
NAND_g _25794_ (.A(cpuregs[4][17]), .B(_00008_[2]), .Y(_05007_));
NAND_g _25795_ (.A(cpuregs[0][17]), .B(_09032_), .Y(_05008_));
AND_g _25796_ (.A(_05007_), .B(_05008_), .Y(_05009_));
NOR_g _25797_ (.A(_00008_[0]), .B(_05009_), .Y(_05010_));
NAND_g _25798_ (.A(_00008_[1]), .B(_05002_), .Y(_05011_));
NOR_g _25799_ (.A(_00008_[1]), .B(_05010_), .Y(_05012_));
NAND_g _25800_ (.A(_05006_), .B(_05012_), .Y(_05013_));
AND_g _25801_ (.A(_09033_), .B(_05013_), .Y(_05014_));
NAND_g _25802_ (.A(_05011_), .B(_05014_), .Y(_05015_));
NAND_g _25803_ (.A(cpuregs[13][17]), .B(_00008_[0]), .Y(_05016_));
NAND_g _25804_ (.A(cpuregs[12][17]), .B(_09030_), .Y(_05017_));
AND_g _25805_ (.A(_00008_[2]), .B(_05017_), .Y(_05018_));
NAND_g _25806_ (.A(_05016_), .B(_05018_), .Y(_05019_));
NAND_g _25807_ (.A(cpuregs[9][17]), .B(_00008_[0]), .Y(_05020_));
NAND_g _25808_ (.A(cpuregs[8][17]), .B(_09030_), .Y(_05021_));
AND_g _25809_ (.A(_09032_), .B(_05021_), .Y(_05022_));
NAND_g _25810_ (.A(_05020_), .B(_05022_), .Y(_05023_));
AND_g _25811_ (.A(_09031_), .B(_05023_), .Y(_05024_));
NAND_g _25812_ (.A(_05019_), .B(_05024_), .Y(_05025_));
NAND_g _25813_ (.A(cpuregs[15][17]), .B(_00008_[0]), .Y(_05026_));
NAND_g _25814_ (.A(cpuregs[14][17]), .B(_09030_), .Y(_05027_));
AND_g _25815_ (.A(_00008_[2]), .B(_05027_), .Y(_05028_));
NAND_g _25816_ (.A(_05026_), .B(_05028_), .Y(_05029_));
NAND_g _25817_ (.A(cpuregs[11][17]), .B(_00008_[0]), .Y(_05030_));
NAND_g _25818_ (.A(cpuregs[10][17]), .B(_09030_), .Y(_05031_));
AND_g _25819_ (.A(_09032_), .B(_05031_), .Y(_05032_));
NAND_g _25820_ (.A(_05030_), .B(_05032_), .Y(_05033_));
AND_g _25821_ (.A(_00008_[1]), .B(_05033_), .Y(_05034_));
NAND_g _25822_ (.A(_05029_), .B(_05034_), .Y(_05035_));
NAND_g _25823_ (.A(_05025_), .B(_05035_), .Y(_05036_));
AND_g _25824_ (.A(_00008_[3]), .B(_05036_), .Y(_05037_));
NOR_g _25825_ (.A(_00008_[4]), .B(_05037_), .Y(_05038_));
NAND_g _25826_ (.A(_05015_), .B(_05038_), .Y(_05039_));
NAND_g _25827_ (.A(cpuregs[25][17]), .B(_09032_), .Y(_05040_));
NAND_g _25828_ (.A(cpuregs[29][17]), .B(_00008_[2]), .Y(_05041_));
AND_g _25829_ (.A(_09031_), .B(_05041_), .Y(_05042_));
NAND_g _25830_ (.A(_05040_), .B(_05042_), .Y(_05043_));
NAND_g _25831_ (.A(cpuregs[31][17]), .B(_00008_[2]), .Y(_05044_));
NAND_g _25832_ (.A(cpuregs[27][17]), .B(_09032_), .Y(_05045_));
AND_g _25833_ (.A(_00008_[1]), .B(_05045_), .Y(_05046_));
NAND_g _25834_ (.A(_05044_), .B(_05046_), .Y(_05047_));
NAND_g _25835_ (.A(_05043_), .B(_05047_), .Y(_05048_));
NAND_g _25836_ (.A(_00008_[0]), .B(_05048_), .Y(_05049_));
NAND_g _25837_ (.A(cpuregs[24][17]), .B(_09032_), .Y(_05050_));
NAND_g _25838_ (.A(cpuregs[28][17]), .B(_00008_[2]), .Y(_05051_));
AND_g _25839_ (.A(_09031_), .B(_05051_), .Y(_05052_));
NAND_g _25840_ (.A(_05050_), .B(_05052_), .Y(_05053_));
NAND_g _25841_ (.A(cpuregs[26][17]), .B(_09032_), .Y(_05054_));
NAND_g _25842_ (.A(cpuregs[30][17]), .B(_00008_[2]), .Y(_05055_));
AND_g _25843_ (.A(_00008_[1]), .B(_05055_), .Y(_05056_));
NAND_g _25844_ (.A(_05054_), .B(_05056_), .Y(_05057_));
NAND_g _25845_ (.A(_05053_), .B(_05057_), .Y(_05058_));
NAND_g _25846_ (.A(_09030_), .B(_05058_), .Y(_05059_));
NAND_g _25847_ (.A(_05049_), .B(_05059_), .Y(_05060_));
NAND_g _25848_ (.A(_00008_[3]), .B(_05060_), .Y(_05061_));
NAND_g _25849_ (.A(cpuregs[17][17]), .B(_09031_), .Y(_05062_));
NAND_g _25850_ (.A(cpuregs[19][17]), .B(_00008_[1]), .Y(_05063_));
AND_g _25851_ (.A(_09032_), .B(_05063_), .Y(_05064_));
NAND_g _25852_ (.A(_05062_), .B(_05064_), .Y(_05065_));
NAND_g _25853_ (.A(cpuregs[21][17]), .B(_09031_), .Y(_05066_));
NAND_g _25854_ (.A(cpuregs[23][17]), .B(_00008_[1]), .Y(_05067_));
AND_g _25855_ (.A(_00008_[2]), .B(_05067_), .Y(_05068_));
NAND_g _25856_ (.A(_05066_), .B(_05068_), .Y(_05069_));
NAND_g _25857_ (.A(_05065_), .B(_05069_), .Y(_05070_));
NAND_g _25858_ (.A(_00008_[0]), .B(_05070_), .Y(_05071_));
NAND_g _25859_ (.A(cpuregs[16][17]), .B(_09031_), .Y(_05072_));
NAND_g _25860_ (.A(cpuregs[18][17]), .B(_00008_[1]), .Y(_05073_));
AND_g _25861_ (.A(_09032_), .B(_05073_), .Y(_05074_));
NAND_g _25862_ (.A(_05072_), .B(_05074_), .Y(_05075_));
NAND_g _25863_ (.A(cpuregs[20][17]), .B(_09031_), .Y(_05076_));
NAND_g _25864_ (.A(cpuregs[22][17]), .B(_00008_[1]), .Y(_05077_));
AND_g _25865_ (.A(_00008_[2]), .B(_05077_), .Y(_05078_));
NAND_g _25866_ (.A(_05076_), .B(_05078_), .Y(_05079_));
NAND_g _25867_ (.A(_05075_), .B(_05079_), .Y(_05080_));
NAND_g _25868_ (.A(_09030_), .B(_05080_), .Y(_05081_));
NAND_g _25869_ (.A(_05071_), .B(_05081_), .Y(_05082_));
AND_g _25870_ (.A(_09033_), .B(_05082_), .Y(_05083_));
NOT_g _25871_ (.A(_05083_), .Y(_05084_));
NAND_g _25872_ (.A(_05061_), .B(_05084_), .Y(_05085_));
NAND_g _25873_ (.A(_00008_[4]), .B(_05085_), .Y(_05086_));
AND_g _25874_ (.A(_14624_), .B(_05086_), .Y(_05087_));
NAND_g _25875_ (.A(_05039_), .B(_05087_), .Y(_05088_));
NAND_g _25876_ (.A(_04993_), .B(_05088_), .Y(_05089_));
NAND_g _25877_ (.A(_10595_), .B(_05089_), .Y(_05090_));
NAND_g _25878_ (.A(pcpi_rs1[16]), .B(_14481_), .Y(_05091_));
AND_g _25879_ (.A(_04760_), .B(_05091_), .Y(_05092_));
NAND_g _25880_ (.A(pcpi_rs1[21]), .B(_14482_), .Y(_05093_));
AND_g _25881_ (.A(_04757_), .B(_05093_), .Y(_05094_));
NAND_g _25882_ (.A(_13880_), .B(_05094_), .Y(_05095_));
NAND_g _25883_ (.A(_13879_), .B(_05092_), .Y(_05096_));
AND_g _25884_ (.A(_13883_), .B(_05095_), .Y(_05097_));
NAND_g _25885_ (.A(_05096_), .B(_05097_), .Y(_05098_));
AND_g _25886_ (.A(_14488_), .B(_05098_), .Y(_05099_));
AND_g _25887_ (.A(_05090_), .B(_05099_), .Y(_05100_));
XOR_g _25888_ (.A(decoded_imm[17]), .B(pcpi_rs1[17]), .Y(_05101_));
XNOR_g _25889_ (.A(_14584_), .B(_05101_), .Y(_05102_));
NAND_g _25890_ (.A(_14614_), .B(_05102_), .Y(_05103_));
AND_g _25891_ (.A(_05100_), .B(_05103_), .Y(_05104_));
NOR_g _25892_ (.A(_04992_), .B(_05104_), .Y(_01035_));
NOR_g _25893_ (.A(pcpi_rs1[18]), .B(_14488_), .Y(_05105_));
XOR_g _25894_ (.A(_14516_), .B(_14586_), .Y(_05106_));
NAND_g _25895_ (.A(_14614_), .B(_05106_), .Y(_05107_));
NAND_g _25896_ (.A(reg_pc[18]), .B(_14617_), .Y(_05108_));
NAND_g _25897_ (.A(cpuregs[13][18]), .B(_00008_[2]), .Y(_05109_));
NAND_g _25898_ (.A(cpuregs[9][18]), .B(_09032_), .Y(_05110_));
NAND_g _25899_ (.A(_05109_), .B(_05110_), .Y(_05111_));
NAND_g _25900_ (.A(_00008_[0]), .B(_05111_), .Y(_05112_));
NAND_g _25901_ (.A(cpuregs[12][18]), .B(_00008_[2]), .Y(_05113_));
NAND_g _25902_ (.A(cpuregs[8][18]), .B(_09032_), .Y(_05114_));
AND_g _25903_ (.A(_05113_), .B(_05114_), .Y(_05115_));
NOR_g _25904_ (.A(_00008_[0]), .B(_05115_), .Y(_05116_));
NAND_g _25905_ (.A(_08913_), .B(_00008_[2]), .Y(_05117_));
NOR_g _25906_ (.A(cpuregs[0][18]), .B(_00008_[2]), .Y(_05118_));
NOR_g _25907_ (.A(_00008_[0]), .B(_05118_), .Y(_05119_));
NAND_g _25908_ (.A(_05117_), .B(_05119_), .Y(_05120_));
NAND_g _25909_ (.A(_08955_), .B(_00008_[2]), .Y(_05121_));
NOR_g _25910_ (.A(cpuregs[1][18]), .B(_00008_[2]), .Y(_05122_));
NOR_g _25911_ (.A(_09030_), .B(_05122_), .Y(_05123_));
NAND_g _25912_ (.A(_05121_), .B(_05123_), .Y(_05124_));
NAND_g _25913_ (.A(cpuregs[11][18]), .B(_09032_), .Y(_05125_));
NAND_g _25914_ (.A(cpuregs[15][18]), .B(_00008_[2]), .Y(_05126_));
NAND_g _25915_ (.A(_05125_), .B(_05126_), .Y(_05127_));
AND_g _25916_ (.A(_00008_[0]), .B(_05127_), .Y(_05128_));
NAND_g _25917_ (.A(cpuregs[14][18]), .B(_00008_[2]), .Y(_05129_));
NAND_g _25918_ (.A(cpuregs[10][18]), .B(_09032_), .Y(_05130_));
AND_g _25919_ (.A(_05129_), .B(_05130_), .Y(_05131_));
NOR_g _25920_ (.A(_00008_[0]), .B(_05131_), .Y(_05132_));
NOR_g _25921_ (.A(_05128_), .B(_05132_), .Y(_05133_));
NAND_g _25922_ (.A(_09012_), .B(_00008_[2]), .Y(_05134_));
NOR_g _25923_ (.A(cpuregs[2][18]), .B(_00008_[2]), .Y(_05135_));
NOR_g _25924_ (.A(_00008_[0]), .B(_05135_), .Y(_05136_));
NAND_g _25925_ (.A(_05134_), .B(_05136_), .Y(_05137_));
NAND_g _25926_ (.A(_08972_), .B(_00008_[2]), .Y(_05138_));
NOR_g _25927_ (.A(cpuregs[3][18]), .B(_00008_[2]), .Y(_05139_));
NOR_g _25928_ (.A(_09030_), .B(_05139_), .Y(_05140_));
NAND_g _25929_ (.A(_05138_), .B(_05140_), .Y(_05141_));
AND_g _25930_ (.A(_05137_), .B(_05141_), .Y(_05142_));
NAND_g _25931_ (.A(_00008_[1]), .B(_05142_), .Y(_05143_));
AND_g _25932_ (.A(_09031_), .B(_05120_), .Y(_05144_));
NAND_g _25933_ (.A(_05124_), .B(_05144_), .Y(_05145_));
AND_g _25934_ (.A(_05143_), .B(_05145_), .Y(_05146_));
NAND_g _25935_ (.A(_09033_), .B(_05146_), .Y(_05147_));
NAND_g _25936_ (.A(_00008_[1]), .B(_05133_), .Y(_05148_));
NOR_g _25937_ (.A(_00008_[1]), .B(_05116_), .Y(_05149_));
NAND_g _25938_ (.A(_05112_), .B(_05149_), .Y(_05150_));
AND_g _25939_ (.A(_00008_[3]), .B(_05150_), .Y(_05151_));
AND_g _25940_ (.A(_05148_), .B(_05151_), .Y(_05152_));
NOR_g _25941_ (.A(_00008_[4]), .B(_05152_), .Y(_05153_));
NAND_g _25942_ (.A(_05147_), .B(_05153_), .Y(_05154_));
NAND_g _25943_ (.A(cpuregs[26][18]), .B(_09032_), .Y(_05155_));
NAND_g _25944_ (.A(cpuregs[30][18]), .B(_00008_[2]), .Y(_05156_));
AND_g _25945_ (.A(_09030_), .B(_05156_), .Y(_05157_));
NAND_g _25946_ (.A(_05155_), .B(_05157_), .Y(_05158_));
NAND_g _25947_ (.A(cpuregs[31][18]), .B(_00008_[2]), .Y(_05159_));
NAND_g _25948_ (.A(cpuregs[27][18]), .B(_09032_), .Y(_05160_));
AND_g _25949_ (.A(_00008_[0]), .B(_05160_), .Y(_05161_));
NAND_g _25950_ (.A(_05159_), .B(_05161_), .Y(_05162_));
NAND_g _25951_ (.A(_05158_), .B(_05162_), .Y(_05163_));
NAND_g _25952_ (.A(_00008_[3]), .B(_05163_), .Y(_05164_));
NAND_g _25953_ (.A(cpuregs[18][18]), .B(_09032_), .Y(_05165_));
NAND_g _25954_ (.A(cpuregs[22][18]), .B(_00008_[2]), .Y(_05166_));
AND_g _25955_ (.A(_09030_), .B(_05166_), .Y(_05167_));
NAND_g _25956_ (.A(_05165_), .B(_05167_), .Y(_05168_));
NAND_g _25957_ (.A(cpuregs[19][18]), .B(_09032_), .Y(_05169_));
NAND_g _25958_ (.A(cpuregs[23][18]), .B(_00008_[2]), .Y(_05170_));
AND_g _25959_ (.A(_00008_[0]), .B(_05170_), .Y(_05171_));
NAND_g _25960_ (.A(_05169_), .B(_05171_), .Y(_05172_));
NAND_g _25961_ (.A(_05168_), .B(_05172_), .Y(_05173_));
NAND_g _25962_ (.A(_09033_), .B(_05173_), .Y(_05174_));
NOR_g _25963_ (.A(cpuregs[25][18]), .B(_00008_[2]), .Y(_05175_));
NAND_g _25964_ (.A(_08878_), .B(_00008_[2]), .Y(_05176_));
NOR_g _25965_ (.A(cpuregs[24][18]), .B(_00008_[2]), .Y(_05177_));
NOR_g _25966_ (.A(cpuregs[28][18]), .B(_09032_), .Y(_05178_));
NOR_g _25967_ (.A(_05177_), .B(_05178_), .Y(_05179_));
NAND_g _25968_ (.A(_00008_[0]), .B(_05176_), .Y(_05180_));
NOR_g _25969_ (.A(_05175_), .B(_05180_), .Y(_05181_));
AND_g _25970_ (.A(_09030_), .B(_05179_), .Y(_05182_));
NOR_g _25971_ (.A(_05181_), .B(_05182_), .Y(_05183_));
NAND_g _25972_ (.A(_00008_[3]), .B(_05183_), .Y(_05184_));
NAND_g _25973_ (.A(cpuregs[20][18]), .B(_00008_[2]), .Y(_05185_));
NAND_g _25974_ (.A(cpuregs[16][18]), .B(_09032_), .Y(_05186_));
AND_g _25975_ (.A(_05185_), .B(_05186_), .Y(_05187_));
NAND_g _25976_ (.A(_09030_), .B(_05187_), .Y(_05188_));
NAND_g _25977_ (.A(cpuregs[21][18]), .B(_00008_[2]), .Y(_05189_));
NAND_g _25978_ (.A(cpuregs[17][18]), .B(_09032_), .Y(_05190_));
AND_g _25979_ (.A(_00008_[0]), .B(_05190_), .Y(_05191_));
NAND_g _25980_ (.A(_05189_), .B(_05191_), .Y(_05192_));
NAND_g _25981_ (.A(_05188_), .B(_05192_), .Y(_05193_));
NAND_g _25982_ (.A(_09033_), .B(_05193_), .Y(_05194_));
AND_g _25983_ (.A(_05184_), .B(_05194_), .Y(_05195_));
NAND_g _25984_ (.A(_09031_), .B(_05195_), .Y(_05196_));
AND_g _25985_ (.A(_00008_[1]), .B(_05174_), .Y(_05197_));
NAND_g _25986_ (.A(_05164_), .B(_05197_), .Y(_05198_));
AND_g _25987_ (.A(_00008_[4]), .B(_05198_), .Y(_05199_));
NAND_g _25988_ (.A(_05196_), .B(_05199_), .Y(_05200_));
AND_g _25989_ (.A(_14624_), .B(_05154_), .Y(_05201_));
NAND_g _25990_ (.A(_05200_), .B(_05201_), .Y(_05202_));
NAND_g _25991_ (.A(_05108_), .B(_05202_), .Y(_05203_));
NAND_g _25992_ (.A(_10595_), .B(_05203_), .Y(_05204_));
NAND_g _25993_ (.A(pcpi_rs1[17]), .B(_14481_), .Y(_05205_));
AND_g _25994_ (.A(_04871_), .B(_05205_), .Y(_05206_));
NAND_g _25995_ (.A(pcpi_rs1[22]), .B(_14482_), .Y(_05207_));
AND_g _25996_ (.A(_04869_), .B(_05207_), .Y(_05208_));
NAND_g _25997_ (.A(_13880_), .B(_05208_), .Y(_05209_));
NAND_g _25998_ (.A(_13879_), .B(_05206_), .Y(_05210_));
AND_g _25999_ (.A(_13883_), .B(_05209_), .Y(_05211_));
NAND_g _26000_ (.A(_05210_), .B(_05211_), .Y(_05212_));
AND_g _26001_ (.A(_14488_), .B(_05212_), .Y(_05213_));
AND_g _26002_ (.A(_05204_), .B(_05213_), .Y(_05214_));
AND_g _26003_ (.A(_05107_), .B(_05214_), .Y(_05215_));
NOR_g _26004_ (.A(_05105_), .B(_05215_), .Y(_01036_));
NOR_g _26005_ (.A(pcpi_rs1[19]), .B(_14488_), .Y(_05216_));
XNOR_g _26006_ (.A(decoded_imm[19]), .B(pcpi_rs1[19]), .Y(_05217_));
NOR_g _26007_ (.A(_14588_), .B(_05217_), .Y(_05218_));
NAND_g _26008_ (.A(_14588_), .B(_05217_), .Y(_05219_));
NAND_g _26009_ (.A(_14614_), .B(_05219_), .Y(_05220_));
NOR_g _26010_ (.A(_05218_), .B(_05220_), .Y(_05221_));
NAND_g _26011_ (.A(reg_pc[19]), .B(_14617_), .Y(_05222_));
NAND_g _26012_ (.A(_08930_), .B(_00008_[2]), .Y(_05223_));
NOR_g _26013_ (.A(cpuregs[9][19]), .B(_00008_[2]), .Y(_05224_));
NOR_g _26014_ (.A(_09030_), .B(_05224_), .Y(_05225_));
AND_g _26015_ (.A(_05223_), .B(_05225_), .Y(_05226_));
NAND_g _26016_ (.A(cpuregs[12][19]), .B(_00008_[2]), .Y(_05227_));
NAND_g _26017_ (.A(cpuregs[8][19]), .B(_09032_), .Y(_05228_));
AND_g _26018_ (.A(_05227_), .B(_05228_), .Y(_05229_));
NOR_g _26019_ (.A(_00008_[0]), .B(_05229_), .Y(_05230_));
NOR_g _26020_ (.A(_05226_), .B(_05230_), .Y(_05231_));
NAND_g _26021_ (.A(_08914_), .B(_00008_[2]), .Y(_05232_));
NOR_g _26022_ (.A(cpuregs[0][19]), .B(_00008_[2]), .Y(_05233_));
NOR_g _26023_ (.A(_00008_[0]), .B(_05233_), .Y(_05234_));
NAND_g _26024_ (.A(_05232_), .B(_05234_), .Y(_05235_));
NAND_g _26025_ (.A(_08956_), .B(_00008_[2]), .Y(_05236_));
NOR_g _26026_ (.A(cpuregs[1][19]), .B(_00008_[2]), .Y(_05237_));
NOR_g _26027_ (.A(_09030_), .B(_05237_), .Y(_05238_));
NAND_g _26028_ (.A(_05236_), .B(_05238_), .Y(_05239_));
NAND_g _26029_ (.A(_08809_), .B(_00008_[2]), .Y(_05240_));
NOR_g _26030_ (.A(cpuregs[11][19]), .B(_00008_[2]), .Y(_05241_));
NOR_g _26031_ (.A(_09030_), .B(_05241_), .Y(_05242_));
NAND_g _26032_ (.A(_05240_), .B(_05242_), .Y(_05243_));
NOR_g _26033_ (.A(cpuregs[10][19]), .B(_00008_[2]), .Y(_05244_));
AND_g _26034_ (.A(_08939_), .B(_00008_[2]), .Y(_05245_));
NOR_g _26035_ (.A(_05244_), .B(_05245_), .Y(_05246_));
NAND_g _26036_ (.A(_09030_), .B(_05246_), .Y(_05247_));
AND_g _26037_ (.A(_05243_), .B(_05247_), .Y(_05248_));
NAND_g _26038_ (.A(_09013_), .B(_00008_[2]), .Y(_05249_));
NOR_g _26039_ (.A(cpuregs[2][19]), .B(_00008_[2]), .Y(_05250_));
NOR_g _26040_ (.A(_00008_[0]), .B(_05250_), .Y(_05251_));
NAND_g _26041_ (.A(_05249_), .B(_05251_), .Y(_05252_));
NAND_g _26042_ (.A(_08973_), .B(_00008_[2]), .Y(_05253_));
NOR_g _26043_ (.A(cpuregs[3][19]), .B(_00008_[2]), .Y(_05254_));
NOR_g _26044_ (.A(_09030_), .B(_05254_), .Y(_05255_));
NAND_g _26045_ (.A(_05253_), .B(_05255_), .Y(_05256_));
AND_g _26046_ (.A(_05252_), .B(_05256_), .Y(_05257_));
AND_g _26047_ (.A(_09031_), .B(_05235_), .Y(_05258_));
NAND_g _26048_ (.A(_05239_), .B(_05258_), .Y(_05259_));
NAND_g _26049_ (.A(_00008_[1]), .B(_05257_), .Y(_05260_));
AND_g _26050_ (.A(_05259_), .B(_05260_), .Y(_05261_));
NAND_g _26051_ (.A(_09033_), .B(_05261_), .Y(_05262_));
NAND_g _26052_ (.A(_00008_[1]), .B(_05248_), .Y(_05263_));
NAND_g _26053_ (.A(_09031_), .B(_05231_), .Y(_05264_));
AND_g _26054_ (.A(_00008_[3]), .B(_05264_), .Y(_05265_));
AND_g _26055_ (.A(_05263_), .B(_05265_), .Y(_05266_));
NOR_g _26056_ (.A(_00008_[4]), .B(_05266_), .Y(_05267_));
NAND_g _26057_ (.A(_05262_), .B(_05267_), .Y(_05268_));
NAND_g _26058_ (.A(_08895_), .B(_00008_[2]), .Y(_05269_));
NOR_g _26059_ (.A(cpuregs[19][19]), .B(_00008_[2]), .Y(_05270_));
NOR_g _26060_ (.A(cpuregs[18][19]), .B(_00008_[2]), .Y(_05271_));
NOR_g _26061_ (.A(cpuregs[22][19]), .B(_09032_), .Y(_05272_));
NOR_g _26062_ (.A(_05271_), .B(_05272_), .Y(_05273_));
NOR_g _26063_ (.A(_09030_), .B(_05270_), .Y(_05274_));
NAND_g _26064_ (.A(_05269_), .B(_05274_), .Y(_05275_));
NAND_g _26065_ (.A(_09030_), .B(_05273_), .Y(_05276_));
AND_g _26066_ (.A(_05275_), .B(_05276_), .Y(_05277_));
NAND_g _26067_ (.A(_00008_[1]), .B(_05277_), .Y(_05278_));
NOR_g _26068_ (.A(cpuregs[17][19]), .B(_00008_[2]), .Y(_05279_));
NAND_g _26069_ (.A(_08994_), .B(_00008_[2]), .Y(_05280_));
NOR_g _26070_ (.A(cpuregs[16][19]), .B(_00008_[2]), .Y(_05281_));
NOR_g _26071_ (.A(cpuregs[20][19]), .B(_09032_), .Y(_05282_));
NOR_g _26072_ (.A(_05281_), .B(_05282_), .Y(_05283_));
NOR_g _26073_ (.A(_09030_), .B(_05279_), .Y(_05284_));
NAND_g _26074_ (.A(_05280_), .B(_05284_), .Y(_05285_));
NAND_g _26075_ (.A(_09030_), .B(_05283_), .Y(_05286_));
AND_g _26076_ (.A(_05285_), .B(_05286_), .Y(_05287_));
NAND_g _26077_ (.A(_09031_), .B(_05287_), .Y(_05288_));
NAND_g _26078_ (.A(_05278_), .B(_05288_), .Y(_05289_));
NAND_g _26079_ (.A(_09033_), .B(_05289_), .Y(_05290_));
NAND_g _26080_ (.A(cpuregs[25][19]), .B(_09031_), .Y(_05291_));
NAND_g _26081_ (.A(cpuregs[27][19]), .B(_00008_[1]), .Y(_05292_));
AND_g _26082_ (.A(_09032_), .B(_05292_), .Y(_05293_));
NAND_g _26083_ (.A(_05291_), .B(_05293_), .Y(_05294_));
NAND_g _26084_ (.A(cpuregs[29][19]), .B(_09031_), .Y(_05295_));
NAND_g _26085_ (.A(cpuregs[31][19]), .B(_00008_[1]), .Y(_05296_));
AND_g _26086_ (.A(_00008_[2]), .B(_05296_), .Y(_05297_));
NAND_g _26087_ (.A(_05295_), .B(_05297_), .Y(_05298_));
NAND_g _26088_ (.A(_05294_), .B(_05298_), .Y(_05299_));
NAND_g _26089_ (.A(_00008_[0]), .B(_05299_), .Y(_05300_));
NAND_g _26090_ (.A(cpuregs[24][19]), .B(_09031_), .Y(_05301_));
NAND_g _26091_ (.A(cpuregs[26][19]), .B(_00008_[1]), .Y(_05302_));
AND_g _26092_ (.A(_09032_), .B(_05302_), .Y(_05303_));
NAND_g _26093_ (.A(_05301_), .B(_05303_), .Y(_05304_));
NAND_g _26094_ (.A(cpuregs[28][19]), .B(_09031_), .Y(_05305_));
NAND_g _26095_ (.A(cpuregs[30][19]), .B(_00008_[1]), .Y(_05306_));
AND_g _26096_ (.A(_00008_[2]), .B(_05306_), .Y(_05307_));
NAND_g _26097_ (.A(_05305_), .B(_05307_), .Y(_05308_));
NAND_g _26098_ (.A(_05304_), .B(_05308_), .Y(_05309_));
NAND_g _26099_ (.A(_09030_), .B(_05309_), .Y(_05310_));
NAND_g _26100_ (.A(_05300_), .B(_05310_), .Y(_05311_));
NAND_g _26101_ (.A(_00008_[3]), .B(_05311_), .Y(_05312_));
NAND_g _26102_ (.A(_05290_), .B(_05312_), .Y(_05313_));
NAND_g _26103_ (.A(_00008_[4]), .B(_05313_), .Y(_05314_));
AND_g _26104_ (.A(_14624_), .B(_05268_), .Y(_05315_));
NAND_g _26105_ (.A(_05314_), .B(_05315_), .Y(_05316_));
NAND_g _26106_ (.A(_05222_), .B(_05316_), .Y(_05317_));
NAND_g _26107_ (.A(_10595_), .B(_05317_), .Y(_05318_));
NAND_g _26108_ (.A(pcpi_rs1[18]), .B(_14481_), .Y(_05319_));
AND_g _26109_ (.A(_04981_), .B(_05319_), .Y(_05320_));
NAND_g _26110_ (.A(pcpi_rs1[23]), .B(_14482_), .Y(_05321_));
AND_g _26111_ (.A(_04979_), .B(_05321_), .Y(_05322_));
NAND_g _26112_ (.A(_13880_), .B(_05322_), .Y(_05323_));
NAND_g _26113_ (.A(_13879_), .B(_05320_), .Y(_05324_));
AND_g _26114_ (.A(_13883_), .B(_05323_), .Y(_05325_));
NAND_g _26115_ (.A(_05324_), .B(_05325_), .Y(_05326_));
AND_g _26116_ (.A(_14488_), .B(_05326_), .Y(_05327_));
NAND_g _26117_ (.A(_05318_), .B(_05327_), .Y(_05328_));
NOR_g _26118_ (.A(_05221_), .B(_05328_), .Y(_05329_));
NOR_g _26119_ (.A(_05216_), .B(_05329_), .Y(_01037_));
NOR_g _26120_ (.A(pcpi_rs1[20]), .B(_14488_), .Y(_05330_));
XOR_g _26121_ (.A(_14512_), .B(_14590_), .Y(_05331_));
NAND_g _26122_ (.A(_14614_), .B(_05331_), .Y(_05332_));
NAND_g _26123_ (.A(reg_pc[20]), .B(_14617_), .Y(_05333_));
NAND_g _26124_ (.A(_08931_), .B(_00008_[2]), .Y(_05334_));
NOR_g _26125_ (.A(cpuregs[9][20]), .B(_00008_[2]), .Y(_05335_));
NOR_g _26126_ (.A(_09030_), .B(_05335_), .Y(_05336_));
AND_g _26127_ (.A(_05334_), .B(_05336_), .Y(_05337_));
NAND_g _26128_ (.A(cpuregs[12][20]), .B(_00008_[2]), .Y(_05338_));
NAND_g _26129_ (.A(cpuregs[8][20]), .B(_09032_), .Y(_05339_));
AND_g _26130_ (.A(_05338_), .B(_05339_), .Y(_05340_));
NOR_g _26131_ (.A(_00008_[0]), .B(_05340_), .Y(_05341_));
NOR_g _26132_ (.A(_05337_), .B(_05341_), .Y(_05342_));
NAND_g _26133_ (.A(_08915_), .B(_00008_[2]), .Y(_05343_));
NOR_g _26134_ (.A(cpuregs[0][20]), .B(_00008_[2]), .Y(_05344_));
NOR_g _26135_ (.A(_00008_[0]), .B(_05344_), .Y(_05345_));
NAND_g _26136_ (.A(_05343_), .B(_05345_), .Y(_05346_));
NAND_g _26137_ (.A(_08957_), .B(_00008_[2]), .Y(_05347_));
NOR_g _26138_ (.A(cpuregs[1][20]), .B(_00008_[2]), .Y(_05348_));
NOR_g _26139_ (.A(_09030_), .B(_05348_), .Y(_05349_));
NAND_g _26140_ (.A(_05347_), .B(_05349_), .Y(_05350_));
NAND_g _26141_ (.A(_08810_), .B(_00008_[2]), .Y(_05351_));
NOR_g _26142_ (.A(cpuregs[11][20]), .B(_00008_[2]), .Y(_05352_));
NOR_g _26143_ (.A(_09030_), .B(_05352_), .Y(_05353_));
NAND_g _26144_ (.A(_05351_), .B(_05353_), .Y(_05354_));
NOR_g _26145_ (.A(cpuregs[10][20]), .B(_00008_[2]), .Y(_05355_));
AND_g _26146_ (.A(_08940_), .B(_00008_[2]), .Y(_05356_));
NOR_g _26147_ (.A(_05355_), .B(_05356_), .Y(_05357_));
NAND_g _26148_ (.A(_09030_), .B(_05357_), .Y(_05358_));
AND_g _26149_ (.A(_05354_), .B(_05358_), .Y(_05359_));
NAND_g _26150_ (.A(_09014_), .B(_00008_[2]), .Y(_05360_));
NOR_g _26151_ (.A(cpuregs[2][20]), .B(_00008_[2]), .Y(_05361_));
NOR_g _26152_ (.A(_00008_[0]), .B(_05361_), .Y(_05362_));
NAND_g _26153_ (.A(_05360_), .B(_05362_), .Y(_05363_));
NAND_g _26154_ (.A(_08974_), .B(_00008_[2]), .Y(_05364_));
NOR_g _26155_ (.A(cpuregs[3][20]), .B(_00008_[2]), .Y(_05365_));
NOR_g _26156_ (.A(_09030_), .B(_05365_), .Y(_05366_));
NAND_g _26157_ (.A(_05364_), .B(_05366_), .Y(_05367_));
AND_g _26158_ (.A(_05363_), .B(_05367_), .Y(_05368_));
AND_g _26159_ (.A(_09031_), .B(_05346_), .Y(_05369_));
NAND_g _26160_ (.A(_05350_), .B(_05369_), .Y(_05370_));
NAND_g _26161_ (.A(_00008_[1]), .B(_05368_), .Y(_05371_));
AND_g _26162_ (.A(_05370_), .B(_05371_), .Y(_05372_));
NAND_g _26163_ (.A(_09033_), .B(_05372_), .Y(_05373_));
NAND_g _26164_ (.A(_00008_[1]), .B(_05359_), .Y(_05374_));
NAND_g _26165_ (.A(_09031_), .B(_05342_), .Y(_05375_));
AND_g _26166_ (.A(_00008_[3]), .B(_05375_), .Y(_05376_));
AND_g _26167_ (.A(_05374_), .B(_05376_), .Y(_05377_));
NOR_g _26168_ (.A(_00008_[4]), .B(_05377_), .Y(_05378_));
NAND_g _26169_ (.A(_05373_), .B(_05378_), .Y(_05379_));
NAND_g _26170_ (.A(_08896_), .B(_00008_[2]), .Y(_05380_));
NOR_g _26171_ (.A(cpuregs[19][20]), .B(_00008_[2]), .Y(_05381_));
NOR_g _26172_ (.A(cpuregs[18][20]), .B(_00008_[2]), .Y(_05382_));
NOR_g _26173_ (.A(cpuregs[22][20]), .B(_09032_), .Y(_05383_));
NOR_g _26174_ (.A(_05382_), .B(_05383_), .Y(_05384_));
NOR_g _26175_ (.A(_09030_), .B(_05381_), .Y(_05385_));
NAND_g _26176_ (.A(_05380_), .B(_05385_), .Y(_05386_));
NAND_g _26177_ (.A(_09030_), .B(_05384_), .Y(_05387_));
AND_g _26178_ (.A(_05386_), .B(_05387_), .Y(_05388_));
NAND_g _26179_ (.A(_00008_[1]), .B(_05388_), .Y(_05389_));
NOR_g _26180_ (.A(cpuregs[17][20]), .B(_00008_[2]), .Y(_05390_));
NAND_g _26181_ (.A(_08995_), .B(_00008_[2]), .Y(_05391_));
NOR_g _26182_ (.A(cpuregs[16][20]), .B(_00008_[2]), .Y(_05392_));
NOR_g _26183_ (.A(cpuregs[20][20]), .B(_09032_), .Y(_05393_));
NOR_g _26184_ (.A(_05392_), .B(_05393_), .Y(_05394_));
NOR_g _26185_ (.A(_09030_), .B(_05390_), .Y(_05395_));
NAND_g _26186_ (.A(_05391_), .B(_05395_), .Y(_05396_));
NAND_g _26187_ (.A(_09030_), .B(_05394_), .Y(_05397_));
AND_g _26188_ (.A(_05396_), .B(_05397_), .Y(_05398_));
NAND_g _26189_ (.A(_09031_), .B(_05398_), .Y(_05399_));
NAND_g _26190_ (.A(_05389_), .B(_05399_), .Y(_05400_));
NAND_g _26191_ (.A(_09033_), .B(_05400_), .Y(_05401_));
NAND_g _26192_ (.A(cpuregs[25][20]), .B(_09031_), .Y(_05402_));
NAND_g _26193_ (.A(cpuregs[27][20]), .B(_00008_[1]), .Y(_05403_));
AND_g _26194_ (.A(_09032_), .B(_05403_), .Y(_05404_));
NAND_g _26195_ (.A(_05402_), .B(_05404_), .Y(_05405_));
NAND_g _26196_ (.A(cpuregs[29][20]), .B(_09031_), .Y(_05406_));
NAND_g _26197_ (.A(cpuregs[31][20]), .B(_00008_[1]), .Y(_05407_));
AND_g _26198_ (.A(_00008_[2]), .B(_05407_), .Y(_05408_));
NAND_g _26199_ (.A(_05406_), .B(_05408_), .Y(_05409_));
NAND_g _26200_ (.A(_05405_), .B(_05409_), .Y(_05410_));
NAND_g _26201_ (.A(_00008_[0]), .B(_05410_), .Y(_05411_));
NAND_g _26202_ (.A(cpuregs[24][20]), .B(_09031_), .Y(_05412_));
NAND_g _26203_ (.A(cpuregs[26][20]), .B(_00008_[1]), .Y(_05413_));
AND_g _26204_ (.A(_09032_), .B(_05413_), .Y(_05414_));
NAND_g _26205_ (.A(_05412_), .B(_05414_), .Y(_05415_));
NAND_g _26206_ (.A(cpuregs[28][20]), .B(_09031_), .Y(_05416_));
NAND_g _26207_ (.A(cpuregs[30][20]), .B(_00008_[1]), .Y(_05417_));
AND_g _26208_ (.A(_00008_[2]), .B(_05417_), .Y(_05418_));
NAND_g _26209_ (.A(_05416_), .B(_05418_), .Y(_05419_));
NAND_g _26210_ (.A(_05415_), .B(_05419_), .Y(_05420_));
NAND_g _26211_ (.A(_09030_), .B(_05420_), .Y(_05421_));
NAND_g _26212_ (.A(_05411_), .B(_05421_), .Y(_05422_));
NAND_g _26213_ (.A(_00008_[3]), .B(_05422_), .Y(_05423_));
NAND_g _26214_ (.A(_05401_), .B(_05423_), .Y(_05424_));
NAND_g _26215_ (.A(_00008_[4]), .B(_05424_), .Y(_05425_));
AND_g _26216_ (.A(_14624_), .B(_05379_), .Y(_05426_));
NAND_g _26217_ (.A(_05425_), .B(_05426_), .Y(_05427_));
NAND_g _26218_ (.A(_05333_), .B(_05427_), .Y(_05428_));
NAND_g _26219_ (.A(_10595_), .B(_05428_), .Y(_05429_));
NAND_g _26220_ (.A(pcpi_rs1[19]), .B(_14481_), .Y(_05430_));
AND_g _26221_ (.A(_05093_), .B(_05430_), .Y(_05431_));
NAND_g _26222_ (.A(_13879_), .B(_05431_), .Y(_05432_));
NAND_g _26223_ (.A(pcpi_rs1[24]), .B(_14482_), .Y(_05433_));
AND_g _26224_ (.A(_05091_), .B(_05433_), .Y(_05434_));
NAND_g _26225_ (.A(_13880_), .B(_05434_), .Y(_05435_));
AND_g _26226_ (.A(_05432_), .B(_05435_), .Y(_05436_));
NAND_g _26227_ (.A(_13883_), .B(_05436_), .Y(_05437_));
AND_g _26228_ (.A(_14488_), .B(_05429_), .Y(_05438_));
AND_g _26229_ (.A(_05437_), .B(_05438_), .Y(_05439_));
AND_g _26230_ (.A(_05332_), .B(_05439_), .Y(_05440_));
NOR_g _26231_ (.A(_05330_), .B(_05440_), .Y(_01038_));
NOR_g _26232_ (.A(pcpi_rs1[21]), .B(_14488_), .Y(_05441_));
XOR_g _26233_ (.A(decoded_imm[21]), .B(pcpi_rs1[21]), .Y(_05442_));
XNOR_g _26234_ (.A(_14592_), .B(_05442_), .Y(_05443_));
NAND_g _26235_ (.A(_14614_), .B(_05443_), .Y(_05444_));
NAND_g _26236_ (.A(reg_pc[21]), .B(_14617_), .Y(_05445_));
NAND_g _26237_ (.A(cpuregs[13][21]), .B(_00008_[2]), .Y(_05446_));
NAND_g _26238_ (.A(cpuregs[9][21]), .B(_09032_), .Y(_05447_));
NAND_g _26239_ (.A(_05446_), .B(_05447_), .Y(_05448_));
NAND_g _26240_ (.A(_00008_[0]), .B(_05448_), .Y(_05449_));
NAND_g _26241_ (.A(cpuregs[12][21]), .B(_00008_[2]), .Y(_05450_));
NAND_g _26242_ (.A(cpuregs[8][21]), .B(_09032_), .Y(_05451_));
AND_g _26243_ (.A(_05450_), .B(_05451_), .Y(_05452_));
NOR_g _26244_ (.A(_00008_[0]), .B(_05452_), .Y(_05453_));
NAND_g _26245_ (.A(_08916_), .B(_00008_[2]), .Y(_05454_));
NOR_g _26246_ (.A(cpuregs[0][21]), .B(_00008_[2]), .Y(_05455_));
NOR_g _26247_ (.A(_00008_[0]), .B(_05455_), .Y(_05456_));
NAND_g _26248_ (.A(_05454_), .B(_05456_), .Y(_05457_));
NAND_g _26249_ (.A(_08958_), .B(_00008_[2]), .Y(_05458_));
NOR_g _26250_ (.A(cpuregs[1][21]), .B(_00008_[2]), .Y(_05459_));
NOR_g _26251_ (.A(_09030_), .B(_05459_), .Y(_05460_));
NAND_g _26252_ (.A(_05458_), .B(_05460_), .Y(_05461_));
NAND_g _26253_ (.A(cpuregs[11][21]), .B(_09032_), .Y(_05462_));
NAND_g _26254_ (.A(cpuregs[15][21]), .B(_00008_[2]), .Y(_05463_));
NAND_g _26255_ (.A(_05462_), .B(_05463_), .Y(_05464_));
AND_g _26256_ (.A(_00008_[0]), .B(_05464_), .Y(_05465_));
NAND_g _26257_ (.A(cpuregs[14][21]), .B(_00008_[2]), .Y(_05466_));
NAND_g _26258_ (.A(cpuregs[10][21]), .B(_09032_), .Y(_05467_));
AND_g _26259_ (.A(_05466_), .B(_05467_), .Y(_05468_));
NOR_g _26260_ (.A(_00008_[0]), .B(_05468_), .Y(_05469_));
NOR_g _26261_ (.A(_05465_), .B(_05469_), .Y(_05470_));
NAND_g _26262_ (.A(_09015_), .B(_00008_[2]), .Y(_05471_));
NOR_g _26263_ (.A(cpuregs[2][21]), .B(_00008_[2]), .Y(_05472_));
NOR_g _26264_ (.A(_00008_[0]), .B(_05472_), .Y(_05473_));
NAND_g _26265_ (.A(_05471_), .B(_05473_), .Y(_05474_));
NAND_g _26266_ (.A(_08975_), .B(_00008_[2]), .Y(_05475_));
NOR_g _26267_ (.A(cpuregs[3][21]), .B(_00008_[2]), .Y(_05476_));
NOR_g _26268_ (.A(_09030_), .B(_05476_), .Y(_05477_));
NAND_g _26269_ (.A(_05475_), .B(_05477_), .Y(_05478_));
AND_g _26270_ (.A(_05474_), .B(_05478_), .Y(_05479_));
AND_g _26271_ (.A(_09031_), .B(_05457_), .Y(_05480_));
NAND_g _26272_ (.A(_05461_), .B(_05480_), .Y(_05481_));
NAND_g _26273_ (.A(_00008_[1]), .B(_05479_), .Y(_05482_));
AND_g _26274_ (.A(_05481_), .B(_05482_), .Y(_05483_));
NAND_g _26275_ (.A(_09033_), .B(_05483_), .Y(_05484_));
NAND_g _26276_ (.A(_00008_[1]), .B(_05470_), .Y(_05485_));
NOR_g _26277_ (.A(_00008_[1]), .B(_05453_), .Y(_05486_));
NAND_g _26278_ (.A(_05449_), .B(_05486_), .Y(_05487_));
AND_g _26279_ (.A(_00008_[3]), .B(_05487_), .Y(_05488_));
AND_g _26280_ (.A(_05485_), .B(_05488_), .Y(_05489_));
NOR_g _26281_ (.A(_00008_[4]), .B(_05489_), .Y(_05490_));
NAND_g _26282_ (.A(_05484_), .B(_05490_), .Y(_05491_));
NAND_g _26283_ (.A(_08897_), .B(_00008_[2]), .Y(_05492_));
NOR_g _26284_ (.A(cpuregs[19][21]), .B(_00008_[2]), .Y(_05493_));
NOR_g _26285_ (.A(cpuregs[18][21]), .B(_00008_[2]), .Y(_05494_));
NOR_g _26286_ (.A(cpuregs[22][21]), .B(_09032_), .Y(_05495_));
NOR_g _26287_ (.A(_05494_), .B(_05495_), .Y(_05496_));
NOR_g _26288_ (.A(_09030_), .B(_05493_), .Y(_05497_));
NAND_g _26289_ (.A(_05492_), .B(_05497_), .Y(_05498_));
NAND_g _26290_ (.A(_09030_), .B(_05496_), .Y(_05499_));
AND_g _26291_ (.A(_05498_), .B(_05499_), .Y(_05500_));
NAND_g _26292_ (.A(_00008_[1]), .B(_05500_), .Y(_05501_));
NOR_g _26293_ (.A(cpuregs[17][21]), .B(_00008_[2]), .Y(_05502_));
NAND_g _26294_ (.A(_08996_), .B(_00008_[2]), .Y(_05503_));
NOR_g _26295_ (.A(cpuregs[16][21]), .B(_00008_[2]), .Y(_05504_));
NOR_g _26296_ (.A(cpuregs[20][21]), .B(_09032_), .Y(_05505_));
NOR_g _26297_ (.A(_05504_), .B(_05505_), .Y(_05506_));
NOR_g _26298_ (.A(_09030_), .B(_05502_), .Y(_05507_));
NAND_g _26299_ (.A(_05503_), .B(_05507_), .Y(_05508_));
NAND_g _26300_ (.A(_09030_), .B(_05506_), .Y(_05509_));
AND_g _26301_ (.A(_05508_), .B(_05509_), .Y(_05510_));
NAND_g _26302_ (.A(_09031_), .B(_05510_), .Y(_05511_));
NAND_g _26303_ (.A(_05501_), .B(_05511_), .Y(_05512_));
NAND_g _26304_ (.A(_09033_), .B(_05512_), .Y(_05513_));
NAND_g _26305_ (.A(cpuregs[25][21]), .B(_09031_), .Y(_05514_));
NAND_g _26306_ (.A(cpuregs[27][21]), .B(_00008_[1]), .Y(_05515_));
AND_g _26307_ (.A(_09032_), .B(_05515_), .Y(_05516_));
NAND_g _26308_ (.A(_05514_), .B(_05516_), .Y(_05517_));
NAND_g _26309_ (.A(cpuregs[29][21]), .B(_09031_), .Y(_05518_));
NAND_g _26310_ (.A(cpuregs[31][21]), .B(_00008_[1]), .Y(_05519_));
AND_g _26311_ (.A(_00008_[2]), .B(_05519_), .Y(_05520_));
NAND_g _26312_ (.A(_05518_), .B(_05520_), .Y(_05521_));
NAND_g _26313_ (.A(_05517_), .B(_05521_), .Y(_05522_));
NAND_g _26314_ (.A(_00008_[0]), .B(_05522_), .Y(_05523_));
NAND_g _26315_ (.A(cpuregs[24][21]), .B(_09031_), .Y(_05524_));
NAND_g _26316_ (.A(cpuregs[26][21]), .B(_00008_[1]), .Y(_05525_));
AND_g _26317_ (.A(_09032_), .B(_05525_), .Y(_05526_));
NAND_g _26318_ (.A(_05524_), .B(_05526_), .Y(_05527_));
NAND_g _26319_ (.A(cpuregs[28][21]), .B(_09031_), .Y(_05528_));
NAND_g _26320_ (.A(cpuregs[30][21]), .B(_00008_[1]), .Y(_05529_));
AND_g _26321_ (.A(_00008_[2]), .B(_05529_), .Y(_05530_));
NAND_g _26322_ (.A(_05528_), .B(_05530_), .Y(_05531_));
NAND_g _26323_ (.A(_05527_), .B(_05531_), .Y(_05532_));
NAND_g _26324_ (.A(_09030_), .B(_05532_), .Y(_05533_));
NAND_g _26325_ (.A(_05523_), .B(_05533_), .Y(_05534_));
NAND_g _26326_ (.A(_00008_[3]), .B(_05534_), .Y(_05535_));
NAND_g _26327_ (.A(_05513_), .B(_05535_), .Y(_05536_));
NAND_g _26328_ (.A(_00008_[4]), .B(_05536_), .Y(_05537_));
AND_g _26329_ (.A(_14624_), .B(_05491_), .Y(_05538_));
NAND_g _26330_ (.A(_05537_), .B(_05538_), .Y(_05539_));
NAND_g _26331_ (.A(_05445_), .B(_05539_), .Y(_05540_));
NAND_g _26332_ (.A(_10595_), .B(_05540_), .Y(_05541_));
NAND_g _26333_ (.A(pcpi_rs1[20]), .B(_14481_), .Y(_05542_));
AND_g _26334_ (.A(_05207_), .B(_05542_), .Y(_05543_));
NAND_g _26335_ (.A(pcpi_rs1[25]), .B(_14482_), .Y(_05544_));
AND_g _26336_ (.A(_05205_), .B(_05544_), .Y(_05545_));
NAND_g _26337_ (.A(_13880_), .B(_05545_), .Y(_05546_));
NAND_g _26338_ (.A(_13879_), .B(_05543_), .Y(_05547_));
AND_g _26339_ (.A(_13883_), .B(_05546_), .Y(_05548_));
NAND_g _26340_ (.A(_05547_), .B(_05548_), .Y(_05549_));
AND_g _26341_ (.A(_14488_), .B(_05549_), .Y(_05550_));
AND_g _26342_ (.A(_05541_), .B(_05550_), .Y(_05551_));
AND_g _26343_ (.A(_05444_), .B(_05551_), .Y(_05552_));
NOR_g _26344_ (.A(_05441_), .B(_05552_), .Y(_01039_));
NOR_g _26345_ (.A(pcpi_rs1[22]), .B(_14488_), .Y(_05553_));
NAND_g _26346_ (.A(reg_pc[22]), .B(_14617_), .Y(_05554_));
NAND_g _26347_ (.A(_08976_), .B(_00008_[2]), .Y(_05555_));
NOR_g _26348_ (.A(cpuregs[3][22]), .B(_00008_[2]), .Y(_05556_));
NOR_g _26349_ (.A(_09030_), .B(_05556_), .Y(_05557_));
AND_g _26350_ (.A(_05555_), .B(_05557_), .Y(_05558_));
NAND_g _26351_ (.A(cpuregs[6][22]), .B(_00008_[2]), .Y(_05559_));
NAND_g _26352_ (.A(cpuregs[2][22]), .B(_09032_), .Y(_05560_));
AND_g _26353_ (.A(_05559_), .B(_05560_), .Y(_05561_));
NOR_g _26354_ (.A(_00008_[0]), .B(_05561_), .Y(_05562_));
NOR_g _26355_ (.A(_05558_), .B(_05562_), .Y(_05563_));
NAND_g _26356_ (.A(cpuregs[5][22]), .B(_00008_[2]), .Y(_05564_));
NAND_g _26357_ (.A(cpuregs[1][22]), .B(_09032_), .Y(_05565_));
NAND_g _26358_ (.A(_05564_), .B(_05565_), .Y(_05566_));
NAND_g _26359_ (.A(_00008_[0]), .B(_05566_), .Y(_05567_));
NAND_g _26360_ (.A(cpuregs[4][22]), .B(_00008_[2]), .Y(_05568_));
NAND_g _26361_ (.A(cpuregs[0][22]), .B(_09032_), .Y(_05569_));
AND_g _26362_ (.A(_05568_), .B(_05569_), .Y(_05570_));
NOR_g _26363_ (.A(_00008_[0]), .B(_05570_), .Y(_05571_));
NAND_g _26364_ (.A(_00008_[1]), .B(_05563_), .Y(_05572_));
NOR_g _26365_ (.A(_00008_[1]), .B(_05571_), .Y(_05573_));
NAND_g _26366_ (.A(_05567_), .B(_05573_), .Y(_05574_));
AND_g _26367_ (.A(_05572_), .B(_05574_), .Y(_05575_));
NAND_g _26368_ (.A(_09033_), .B(_05575_), .Y(_05576_));
NAND_g _26369_ (.A(cpuregs[13][22]), .B(_00008_[0]), .Y(_05577_));
NAND_g _26370_ (.A(cpuregs[12][22]), .B(_09030_), .Y(_05578_));
AND_g _26371_ (.A(_00008_[2]), .B(_05578_), .Y(_05579_));
NAND_g _26372_ (.A(_05577_), .B(_05579_), .Y(_05580_));
NAND_g _26373_ (.A(cpuregs[9][22]), .B(_00008_[0]), .Y(_05581_));
NAND_g _26374_ (.A(cpuregs[8][22]), .B(_09030_), .Y(_05582_));
AND_g _26375_ (.A(_09032_), .B(_05582_), .Y(_05583_));
NAND_g _26376_ (.A(_05581_), .B(_05583_), .Y(_05584_));
AND_g _26377_ (.A(_09031_), .B(_05584_), .Y(_05585_));
NAND_g _26378_ (.A(_05580_), .B(_05585_), .Y(_05586_));
NAND_g _26379_ (.A(cpuregs[15][22]), .B(_00008_[0]), .Y(_05587_));
NAND_g _26380_ (.A(cpuregs[14][22]), .B(_09030_), .Y(_05588_));
AND_g _26381_ (.A(_00008_[2]), .B(_05588_), .Y(_05589_));
NAND_g _26382_ (.A(_05587_), .B(_05589_), .Y(_05590_));
NAND_g _26383_ (.A(cpuregs[11][22]), .B(_00008_[0]), .Y(_05591_));
NAND_g _26384_ (.A(cpuregs[10][22]), .B(_09030_), .Y(_05592_));
AND_g _26385_ (.A(_09032_), .B(_05592_), .Y(_05593_));
NAND_g _26386_ (.A(_05591_), .B(_05593_), .Y(_05594_));
AND_g _26387_ (.A(_00008_[1]), .B(_05594_), .Y(_05595_));
NAND_g _26388_ (.A(_05590_), .B(_05595_), .Y(_05596_));
NAND_g _26389_ (.A(_05586_), .B(_05596_), .Y(_05597_));
AND_g _26390_ (.A(_00008_[3]), .B(_05597_), .Y(_05598_));
NOR_g _26391_ (.A(_00008_[4]), .B(_05598_), .Y(_05599_));
NAND_g _26392_ (.A(_05576_), .B(_05599_), .Y(_05600_));
NAND_g _26393_ (.A(cpuregs[26][22]), .B(_09032_), .Y(_05601_));
NAND_g _26394_ (.A(cpuregs[30][22]), .B(_00008_[2]), .Y(_05602_));
AND_g _26395_ (.A(_09030_), .B(_05602_), .Y(_05603_));
NAND_g _26396_ (.A(_05601_), .B(_05603_), .Y(_05604_));
NAND_g _26397_ (.A(cpuregs[31][22]), .B(_00008_[2]), .Y(_05605_));
NAND_g _26398_ (.A(cpuregs[27][22]), .B(_09032_), .Y(_05606_));
AND_g _26399_ (.A(_00008_[0]), .B(_05606_), .Y(_05607_));
NAND_g _26400_ (.A(_05605_), .B(_05607_), .Y(_05608_));
NAND_g _26401_ (.A(_05604_), .B(_05608_), .Y(_05609_));
NAND_g _26402_ (.A(_00008_[3]), .B(_05609_), .Y(_05610_));
NAND_g _26403_ (.A(cpuregs[18][22]), .B(_09032_), .Y(_05611_));
NAND_g _26404_ (.A(cpuregs[22][22]), .B(_00008_[2]), .Y(_05612_));
AND_g _26405_ (.A(_09030_), .B(_05612_), .Y(_05613_));
NAND_g _26406_ (.A(_05611_), .B(_05613_), .Y(_05614_));
NAND_g _26407_ (.A(cpuregs[19][22]), .B(_09032_), .Y(_05615_));
NAND_g _26408_ (.A(cpuregs[23][22]), .B(_00008_[2]), .Y(_05616_));
AND_g _26409_ (.A(_00008_[0]), .B(_05616_), .Y(_05617_));
NAND_g _26410_ (.A(_05615_), .B(_05617_), .Y(_05618_));
NAND_g _26411_ (.A(_05614_), .B(_05618_), .Y(_05619_));
NAND_g _26412_ (.A(_09033_), .B(_05619_), .Y(_05620_));
AND_g _26413_ (.A(_05610_), .B(_05620_), .Y(_05621_));
NAND_g _26414_ (.A(cpuregs[24][22]), .B(_09032_), .Y(_05622_));
NAND_g _26415_ (.A(cpuregs[28][22]), .B(_00008_[2]), .Y(_05623_));
AND_g _26416_ (.A(_09030_), .B(_05623_), .Y(_05624_));
NAND_g _26417_ (.A(_05622_), .B(_05624_), .Y(_05625_));
NAND_g _26418_ (.A(cpuregs[29][22]), .B(_00008_[2]), .Y(_05626_));
NAND_g _26419_ (.A(cpuregs[25][22]), .B(_09032_), .Y(_05627_));
AND_g _26420_ (.A(_00008_[0]), .B(_05627_), .Y(_05628_));
NAND_g _26421_ (.A(_05626_), .B(_05628_), .Y(_05629_));
NAND_g _26422_ (.A(_05625_), .B(_05629_), .Y(_05630_));
NAND_g _26423_ (.A(_00008_[3]), .B(_05630_), .Y(_05631_));
NAND_g _26424_ (.A(cpuregs[16][22]), .B(_09032_), .Y(_05632_));
NAND_g _26425_ (.A(cpuregs[20][22]), .B(_00008_[2]), .Y(_05633_));
AND_g _26426_ (.A(_09030_), .B(_05633_), .Y(_05634_));
NAND_g _26427_ (.A(_05632_), .B(_05634_), .Y(_05635_));
NAND_g _26428_ (.A(cpuregs[17][22]), .B(_09032_), .Y(_05636_));
NAND_g _26429_ (.A(cpuregs[21][22]), .B(_00008_[2]), .Y(_05637_));
AND_g _26430_ (.A(_00008_[0]), .B(_05637_), .Y(_05638_));
NAND_g _26431_ (.A(_05636_), .B(_05638_), .Y(_05639_));
NAND_g _26432_ (.A(_05635_), .B(_05639_), .Y(_05640_));
NAND_g _26433_ (.A(_09033_), .B(_05640_), .Y(_05641_));
AND_g _26434_ (.A(_05631_), .B(_05641_), .Y(_05642_));
NAND_g _26435_ (.A(_00008_[1]), .B(_05621_), .Y(_05643_));
NAND_g _26436_ (.A(_09031_), .B(_05642_), .Y(_05644_));
AND_g _26437_ (.A(_00008_[4]), .B(_05643_), .Y(_05645_));
NAND_g _26438_ (.A(_05644_), .B(_05645_), .Y(_05646_));
AND_g _26439_ (.A(_14624_), .B(_05646_), .Y(_05647_));
NAND_g _26440_ (.A(_05600_), .B(_05647_), .Y(_05648_));
NAND_g _26441_ (.A(_05554_), .B(_05648_), .Y(_05649_));
NAND_g _26442_ (.A(_10595_), .B(_05649_), .Y(_05650_));
NAND_g _26443_ (.A(pcpi_rs1[21]), .B(_14481_), .Y(_05651_));
AND_g _26444_ (.A(_05321_), .B(_05651_), .Y(_05652_));
NAND_g _26445_ (.A(pcpi_rs1[26]), .B(_14482_), .Y(_05653_));
AND_g _26446_ (.A(_05319_), .B(_05653_), .Y(_05654_));
NAND_g _26447_ (.A(_13880_), .B(_05654_), .Y(_05655_));
NAND_g _26448_ (.A(_13879_), .B(_05652_), .Y(_05656_));
AND_g _26449_ (.A(_13883_), .B(_05655_), .Y(_05657_));
NAND_g _26450_ (.A(_05656_), .B(_05657_), .Y(_05658_));
AND_g _26451_ (.A(_14488_), .B(_05658_), .Y(_05659_));
AND_g _26452_ (.A(_05650_), .B(_05659_), .Y(_05660_));
XOR_g _26453_ (.A(_14508_), .B(_14594_), .Y(_05661_));
NAND_g _26454_ (.A(_14614_), .B(_05661_), .Y(_05662_));
AND_g _26455_ (.A(_05660_), .B(_05662_), .Y(_05663_));
NOR_g _26456_ (.A(_05553_), .B(_05663_), .Y(_01040_));
NOR_g _26457_ (.A(pcpi_rs1[23]), .B(_14488_), .Y(_05664_));
NAND_g _26458_ (.A(reg_pc[23]), .B(_14617_), .Y(_05665_));
NAND_g _26459_ (.A(cpuregs[7][23]), .B(_00008_[2]), .Y(_05666_));
NAND_g _26460_ (.A(cpuregs[3][23]), .B(_09032_), .Y(_05667_));
AND_g _26461_ (.A(_05666_), .B(_05667_), .Y(_05668_));
NAND_g _26462_ (.A(cpuregs[6][23]), .B(_00008_[2]), .Y(_05669_));
NAND_g _26463_ (.A(cpuregs[2][23]), .B(_09032_), .Y(_05670_));
AND_g _26464_ (.A(_05669_), .B(_05670_), .Y(_05671_));
NAND_g _26465_ (.A(_09030_), .B(_05671_), .Y(_05672_));
NAND_g _26466_ (.A(_00008_[0]), .B(_05668_), .Y(_05673_));
NAND_g _26467_ (.A(_05672_), .B(_05673_), .Y(_05674_));
NAND_g _26468_ (.A(cpuregs[4][23]), .B(_00008_[2]), .Y(_05675_));
NAND_g _26469_ (.A(cpuregs[0][23]), .B(_09032_), .Y(_05676_));
AND_g _26470_ (.A(_09030_), .B(_05676_), .Y(_05677_));
NAND_g _26471_ (.A(_05675_), .B(_05677_), .Y(_05678_));
NAND_g _26472_ (.A(cpuregs[1][23]), .B(_09032_), .Y(_05679_));
NAND_g _26473_ (.A(cpuregs[5][23]), .B(_00008_[2]), .Y(_05680_));
AND_g _26474_ (.A(_00008_[0]), .B(_05680_), .Y(_05681_));
NAND_g _26475_ (.A(_05679_), .B(_05681_), .Y(_05682_));
NAND_g _26476_ (.A(_05678_), .B(_05682_), .Y(_05683_));
NAND_g _26477_ (.A(cpuregs[11][23]), .B(_09032_), .Y(_05684_));
NAND_g _26478_ (.A(cpuregs[15][23]), .B(_00008_[2]), .Y(_05685_));
NAND_g _26479_ (.A(_05684_), .B(_05685_), .Y(_05686_));
NAND_g _26480_ (.A(_00008_[0]), .B(_05686_), .Y(_05687_));
NAND_g _26481_ (.A(cpuregs[14][23]), .B(_00008_[2]), .Y(_05688_));
NAND_g _26482_ (.A(cpuregs[10][23]), .B(_09032_), .Y(_05689_));
NAND_g _26483_ (.A(_05688_), .B(_05689_), .Y(_05690_));
NAND_g _26484_ (.A(_09030_), .B(_05690_), .Y(_05691_));
AND_g _26485_ (.A(_05687_), .B(_05691_), .Y(_05692_));
NAND_g _26486_ (.A(_08882_), .B(_00008_[2]), .Y(_05693_));
NOR_g _26487_ (.A(cpuregs[8][23]), .B(_00008_[2]), .Y(_05694_));
NOR_g _26488_ (.A(_00008_[0]), .B(_05694_), .Y(_05695_));
NAND_g _26489_ (.A(_05693_), .B(_05695_), .Y(_05696_));
NAND_g _26490_ (.A(_08932_), .B(_00008_[2]), .Y(_05697_));
NOR_g _26491_ (.A(cpuregs[9][23]), .B(_00008_[2]), .Y(_05698_));
NOR_g _26492_ (.A(_09030_), .B(_05698_), .Y(_05699_));
NAND_g _26493_ (.A(_05697_), .B(_05699_), .Y(_05700_));
AND_g _26494_ (.A(_05696_), .B(_05700_), .Y(_05701_));
NAND_g _26495_ (.A(_09033_), .B(_05683_), .Y(_05702_));
NAND_g _26496_ (.A(_00008_[3]), .B(_05701_), .Y(_05703_));
AND_g _26497_ (.A(_09031_), .B(_05703_), .Y(_05704_));
NAND_g _26498_ (.A(_05702_), .B(_05704_), .Y(_05705_));
NAND_g _26499_ (.A(_00008_[3]), .B(_05692_), .Y(_05706_));
NAND_g _26500_ (.A(_09033_), .B(_05674_), .Y(_05707_));
AND_g _26501_ (.A(_05706_), .B(_05707_), .Y(_05708_));
AND_g _26502_ (.A(_00008_[1]), .B(_05708_), .Y(_05709_));
NOR_g _26503_ (.A(_00008_[4]), .B(_05709_), .Y(_05710_));
NAND_g _26504_ (.A(_05705_), .B(_05710_), .Y(_05711_));
NAND_g _26505_ (.A(_08899_), .B(_00008_[2]), .Y(_05712_));
NOR_g _26506_ (.A(cpuregs[19][23]), .B(_00008_[2]), .Y(_05713_));
NOR_g _26507_ (.A(cpuregs[18][23]), .B(_00008_[2]), .Y(_05714_));
AND_g _26508_ (.A(_08924_), .B(_00008_[2]), .Y(_05715_));
NOR_g _26509_ (.A(_05714_), .B(_05715_), .Y(_05716_));
NOR_g _26510_ (.A(_09030_), .B(_05713_), .Y(_05717_));
NAND_g _26511_ (.A(_05712_), .B(_05717_), .Y(_05718_));
NAND_g _26512_ (.A(_09030_), .B(_05716_), .Y(_05719_));
AND_g _26513_ (.A(_05718_), .B(_05719_), .Y(_05720_));
NAND_g _26514_ (.A(_00008_[1]), .B(_05720_), .Y(_05721_));
NOR_g _26515_ (.A(cpuregs[17][23]), .B(_00008_[2]), .Y(_05722_));
NAND_g _26516_ (.A(_08998_), .B(_00008_[2]), .Y(_05723_));
NOR_g _26517_ (.A(cpuregs[16][23]), .B(_00008_[2]), .Y(_05724_));
AND_g _26518_ (.A(_08850_), .B(_00008_[2]), .Y(_05725_));
NOR_g _26519_ (.A(_05724_), .B(_05725_), .Y(_05726_));
NOR_g _26520_ (.A(_09030_), .B(_05722_), .Y(_05727_));
NAND_g _26521_ (.A(_05723_), .B(_05727_), .Y(_05728_));
NAND_g _26522_ (.A(_09030_), .B(_05726_), .Y(_05729_));
AND_g _26523_ (.A(_05728_), .B(_05729_), .Y(_05730_));
NAND_g _26524_ (.A(_09031_), .B(_05730_), .Y(_05731_));
NAND_g _26525_ (.A(_05721_), .B(_05731_), .Y(_05732_));
NAND_g _26526_ (.A(_09033_), .B(_05732_), .Y(_05733_));
NAND_g _26527_ (.A(cpuregs[25][23]), .B(_09031_), .Y(_05734_));
NAND_g _26528_ (.A(cpuregs[27][23]), .B(_00008_[1]), .Y(_05735_));
AND_g _26529_ (.A(_09032_), .B(_05735_), .Y(_05736_));
NAND_g _26530_ (.A(_05734_), .B(_05736_), .Y(_05737_));
NAND_g _26531_ (.A(cpuregs[29][23]), .B(_09031_), .Y(_05738_));
NAND_g _26532_ (.A(cpuregs[31][23]), .B(_00008_[1]), .Y(_05739_));
AND_g _26533_ (.A(_00008_[2]), .B(_05739_), .Y(_05740_));
NAND_g _26534_ (.A(_05738_), .B(_05740_), .Y(_05741_));
NAND_g _26535_ (.A(_05737_), .B(_05741_), .Y(_05742_));
NAND_g _26536_ (.A(_00008_[0]), .B(_05742_), .Y(_05743_));
NAND_g _26537_ (.A(cpuregs[24][23]), .B(_09031_), .Y(_05744_));
NAND_g _26538_ (.A(cpuregs[26][23]), .B(_00008_[1]), .Y(_05745_));
AND_g _26539_ (.A(_09032_), .B(_05745_), .Y(_05746_));
NAND_g _26540_ (.A(_05744_), .B(_05746_), .Y(_05747_));
NAND_g _26541_ (.A(cpuregs[28][23]), .B(_09031_), .Y(_05748_));
NAND_g _26542_ (.A(cpuregs[30][23]), .B(_00008_[1]), .Y(_05749_));
AND_g _26543_ (.A(_00008_[2]), .B(_05749_), .Y(_05750_));
NAND_g _26544_ (.A(_05748_), .B(_05750_), .Y(_05751_));
NAND_g _26545_ (.A(_05747_), .B(_05751_), .Y(_05752_));
NAND_g _26546_ (.A(_09030_), .B(_05752_), .Y(_05753_));
NAND_g _26547_ (.A(_05743_), .B(_05753_), .Y(_05754_));
NAND_g _26548_ (.A(_00008_[3]), .B(_05754_), .Y(_05755_));
NAND_g _26549_ (.A(_05733_), .B(_05755_), .Y(_05756_));
NAND_g _26550_ (.A(_00008_[4]), .B(_05756_), .Y(_05757_));
AND_g _26551_ (.A(_14624_), .B(_05711_), .Y(_05758_));
NAND_g _26552_ (.A(_05757_), .B(_05758_), .Y(_05759_));
NAND_g _26553_ (.A(_05665_), .B(_05759_), .Y(_05760_));
NAND_g _26554_ (.A(_10595_), .B(_05760_), .Y(_05761_));
NAND_g _26555_ (.A(pcpi_rs1[22]), .B(_14481_), .Y(_05762_));
AND_g _26556_ (.A(_05433_), .B(_05762_), .Y(_05763_));
NAND_g _26557_ (.A(pcpi_rs1[27]), .B(_14482_), .Y(_05764_));
AND_g _26558_ (.A(_05430_), .B(_05764_), .Y(_05765_));
NAND_g _26559_ (.A(_13880_), .B(_05765_), .Y(_05766_));
NAND_g _26560_ (.A(_13879_), .B(_05763_), .Y(_05767_));
AND_g _26561_ (.A(_13883_), .B(_05766_), .Y(_05768_));
NAND_g _26562_ (.A(_05767_), .B(_05768_), .Y(_05769_));
AND_g _26563_ (.A(_14488_), .B(_05769_), .Y(_05770_));
AND_g _26564_ (.A(_05761_), .B(_05770_), .Y(_05771_));
XOR_g _26565_ (.A(decoded_imm[23]), .B(pcpi_rs1[23]), .Y(_05772_));
XNOR_g _26566_ (.A(_14596_), .B(_05772_), .Y(_05773_));
NAND_g _26567_ (.A(_14614_), .B(_05773_), .Y(_05774_));
AND_g _26568_ (.A(_05771_), .B(_05774_), .Y(_05775_));
NOR_g _26569_ (.A(_05664_), .B(_05775_), .Y(_01041_));
NOR_g _26570_ (.A(pcpi_rs1[24]), .B(_14488_), .Y(_05776_));
XOR_g _26571_ (.A(_14504_), .B(_14598_), .Y(_05777_));
NAND_g _26572_ (.A(_14614_), .B(_05777_), .Y(_05778_));
NAND_g _26573_ (.A(reg_pc[24]), .B(_14617_), .Y(_05779_));
NAND_g _26574_ (.A(_08977_), .B(_00008_[2]), .Y(_05780_));
NOR_g _26575_ (.A(cpuregs[3][24]), .B(_00008_[2]), .Y(_05781_));
NOR_g _26576_ (.A(_09030_), .B(_05781_), .Y(_05782_));
AND_g _26577_ (.A(_05780_), .B(_05782_), .Y(_05783_));
NAND_g _26578_ (.A(cpuregs[6][24]), .B(_00008_[2]), .Y(_05784_));
NAND_g _26579_ (.A(cpuregs[2][24]), .B(_09032_), .Y(_05785_));
AND_g _26580_ (.A(_05784_), .B(_05785_), .Y(_05786_));
NOR_g _26581_ (.A(_00008_[0]), .B(_05786_), .Y(_05787_));
NOR_g _26582_ (.A(_05783_), .B(_05787_), .Y(_05788_));
NAND_g _26583_ (.A(_08959_), .B(_00008_[2]), .Y(_05789_));
NOR_g _26584_ (.A(cpuregs[1][24]), .B(_00008_[2]), .Y(_05790_));
NOR_g _26585_ (.A(_09030_), .B(_05790_), .Y(_05791_));
AND_g _26586_ (.A(_05789_), .B(_05791_), .Y(_05792_));
NAND_g _26587_ (.A(cpuregs[4][24]), .B(_00008_[2]), .Y(_05793_));
NAND_g _26588_ (.A(cpuregs[0][24]), .B(_09032_), .Y(_05794_));
AND_g _26589_ (.A(_05793_), .B(_05794_), .Y(_05795_));
NOR_g _26590_ (.A(_00008_[0]), .B(_05795_), .Y(_05796_));
NOR_g _26591_ (.A(_05792_), .B(_05796_), .Y(_05797_));
NAND_g _26592_ (.A(_00008_[1]), .B(_05788_), .Y(_05798_));
NAND_g _26593_ (.A(_09031_), .B(_05797_), .Y(_05799_));
AND_g _26594_ (.A(_05798_), .B(_05799_), .Y(_05800_));
NAND_g _26595_ (.A(_09033_), .B(_05800_), .Y(_05801_));
NAND_g _26596_ (.A(cpuregs[13][24]), .B(_00008_[0]), .Y(_05802_));
NAND_g _26597_ (.A(cpuregs[12][24]), .B(_09030_), .Y(_05803_));
AND_g _26598_ (.A(_00008_[2]), .B(_05803_), .Y(_05804_));
NAND_g _26599_ (.A(_05802_), .B(_05804_), .Y(_05805_));
NAND_g _26600_ (.A(cpuregs[9][24]), .B(_00008_[0]), .Y(_05806_));
NAND_g _26601_ (.A(cpuregs[8][24]), .B(_09030_), .Y(_05807_));
AND_g _26602_ (.A(_09032_), .B(_05807_), .Y(_05808_));
NAND_g _26603_ (.A(_05806_), .B(_05808_), .Y(_05809_));
AND_g _26604_ (.A(_09031_), .B(_05809_), .Y(_05810_));
NAND_g _26605_ (.A(_05805_), .B(_05810_), .Y(_05811_));
NAND_g _26606_ (.A(cpuregs[15][24]), .B(_00008_[0]), .Y(_05812_));
NAND_g _26607_ (.A(cpuregs[14][24]), .B(_09030_), .Y(_05813_));
AND_g _26608_ (.A(_00008_[2]), .B(_05813_), .Y(_05814_));
NAND_g _26609_ (.A(_05812_), .B(_05814_), .Y(_05815_));
NAND_g _26610_ (.A(cpuregs[11][24]), .B(_00008_[0]), .Y(_05816_));
NAND_g _26611_ (.A(cpuregs[10][24]), .B(_09030_), .Y(_05817_));
AND_g _26612_ (.A(_09032_), .B(_05817_), .Y(_05818_));
NAND_g _26613_ (.A(_05816_), .B(_05818_), .Y(_05819_));
AND_g _26614_ (.A(_00008_[1]), .B(_05819_), .Y(_05820_));
NAND_g _26615_ (.A(_05815_), .B(_05820_), .Y(_05821_));
NAND_g _26616_ (.A(_05811_), .B(_05821_), .Y(_05822_));
AND_g _26617_ (.A(_00008_[3]), .B(_05822_), .Y(_05823_));
NOR_g _26618_ (.A(_00008_[4]), .B(_05823_), .Y(_05824_));
NAND_g _26619_ (.A(_05801_), .B(_05824_), .Y(_05825_));
NAND_g _26620_ (.A(cpuregs[25][24]), .B(_09032_), .Y(_05826_));
NAND_g _26621_ (.A(cpuregs[29][24]), .B(_00008_[2]), .Y(_05827_));
AND_g _26622_ (.A(_09031_), .B(_05827_), .Y(_05828_));
NAND_g _26623_ (.A(_05826_), .B(_05828_), .Y(_05829_));
NAND_g _26624_ (.A(cpuregs[31][24]), .B(_00008_[2]), .Y(_05830_));
NAND_g _26625_ (.A(cpuregs[27][24]), .B(_09032_), .Y(_05831_));
AND_g _26626_ (.A(_00008_[1]), .B(_05831_), .Y(_05832_));
NAND_g _26627_ (.A(_05830_), .B(_05832_), .Y(_05833_));
NAND_g _26628_ (.A(_05829_), .B(_05833_), .Y(_05834_));
NAND_g _26629_ (.A(_00008_[0]), .B(_05834_), .Y(_05835_));
NAND_g _26630_ (.A(cpuregs[24][24]), .B(_09032_), .Y(_05836_));
NAND_g _26631_ (.A(cpuregs[28][24]), .B(_00008_[2]), .Y(_05837_));
AND_g _26632_ (.A(_09031_), .B(_05837_), .Y(_05838_));
NAND_g _26633_ (.A(_05836_), .B(_05838_), .Y(_05839_));
NAND_g _26634_ (.A(cpuregs[26][24]), .B(_09032_), .Y(_05840_));
NAND_g _26635_ (.A(cpuregs[30][24]), .B(_00008_[2]), .Y(_05841_));
AND_g _26636_ (.A(_00008_[1]), .B(_05841_), .Y(_05842_));
NAND_g _26637_ (.A(_05840_), .B(_05842_), .Y(_05843_));
NAND_g _26638_ (.A(_05839_), .B(_05843_), .Y(_05844_));
NAND_g _26639_ (.A(_09030_), .B(_05844_), .Y(_05845_));
NAND_g _26640_ (.A(_05835_), .B(_05845_), .Y(_05846_));
NAND_g _26641_ (.A(_00008_[3]), .B(_05846_), .Y(_05847_));
NAND_g _26642_ (.A(cpuregs[17][24]), .B(_09031_), .Y(_05848_));
NAND_g _26643_ (.A(cpuregs[19][24]), .B(_00008_[1]), .Y(_05849_));
AND_g _26644_ (.A(_09032_), .B(_05849_), .Y(_05850_));
NAND_g _26645_ (.A(_05848_), .B(_05850_), .Y(_05851_));
NAND_g _26646_ (.A(cpuregs[21][24]), .B(_09031_), .Y(_05852_));
NAND_g _26647_ (.A(cpuregs[23][24]), .B(_00008_[1]), .Y(_05853_));
AND_g _26648_ (.A(_00008_[2]), .B(_05853_), .Y(_05854_));
NAND_g _26649_ (.A(_05852_), .B(_05854_), .Y(_05855_));
NAND_g _26650_ (.A(_05851_), .B(_05855_), .Y(_05856_));
NAND_g _26651_ (.A(_00008_[0]), .B(_05856_), .Y(_05857_));
NAND_g _26652_ (.A(cpuregs[16][24]), .B(_09031_), .Y(_05858_));
NAND_g _26653_ (.A(cpuregs[18][24]), .B(_00008_[1]), .Y(_05859_));
AND_g _26654_ (.A(_09032_), .B(_05859_), .Y(_05860_));
NAND_g _26655_ (.A(_05858_), .B(_05860_), .Y(_05861_));
NAND_g _26656_ (.A(cpuregs[20][24]), .B(_09031_), .Y(_05862_));
NAND_g _26657_ (.A(cpuregs[22][24]), .B(_00008_[1]), .Y(_05863_));
AND_g _26658_ (.A(_00008_[2]), .B(_05863_), .Y(_05864_));
NAND_g _26659_ (.A(_05862_), .B(_05864_), .Y(_05865_));
NAND_g _26660_ (.A(_05861_), .B(_05865_), .Y(_05866_));
NAND_g _26661_ (.A(_09030_), .B(_05866_), .Y(_05867_));
NAND_g _26662_ (.A(_05857_), .B(_05867_), .Y(_05868_));
AND_g _26663_ (.A(_09033_), .B(_05868_), .Y(_05869_));
NOT_g _26664_ (.A(_05869_), .Y(_05870_));
NAND_g _26665_ (.A(_05847_), .B(_05870_), .Y(_05871_));
NAND_g _26666_ (.A(_00008_[4]), .B(_05871_), .Y(_05872_));
AND_g _26667_ (.A(_14624_), .B(_05872_), .Y(_05873_));
NAND_g _26668_ (.A(_05825_), .B(_05873_), .Y(_05874_));
NAND_g _26669_ (.A(_05779_), .B(_05874_), .Y(_05875_));
NAND_g _26670_ (.A(_10595_), .B(_05875_), .Y(_05876_));
NAND_g _26671_ (.A(pcpi_rs1[23]), .B(_14481_), .Y(_05877_));
AND_g _26672_ (.A(_05544_), .B(_05877_), .Y(_05878_));
NAND_g _26673_ (.A(pcpi_rs1[28]), .B(_14482_), .Y(_05879_));
AND_g _26674_ (.A(_05542_), .B(_05879_), .Y(_05880_));
NAND_g _26675_ (.A(_13880_), .B(_05880_), .Y(_05881_));
NAND_g _26676_ (.A(_13879_), .B(_05878_), .Y(_05882_));
AND_g _26677_ (.A(_13883_), .B(_05881_), .Y(_05883_));
NAND_g _26678_ (.A(_05882_), .B(_05883_), .Y(_05884_));
AND_g _26679_ (.A(_14488_), .B(_05884_), .Y(_05885_));
AND_g _26680_ (.A(_05876_), .B(_05885_), .Y(_05886_));
AND_g _26681_ (.A(_05778_), .B(_05886_), .Y(_05887_));
NOR_g _26682_ (.A(_05776_), .B(_05887_), .Y(_01042_));
NOR_g _26683_ (.A(pcpi_rs1[25]), .B(_14488_), .Y(_05888_));
XOR_g _26684_ (.A(decoded_imm[25]), .B(pcpi_rs1[25]), .Y(_05889_));
XNOR_g _26685_ (.A(_14600_), .B(_05889_), .Y(_05890_));
NAND_g _26686_ (.A(_14614_), .B(_05890_), .Y(_05891_));
NAND_g _26687_ (.A(reg_pc[25]), .B(_14617_), .Y(_05892_));
NAND_g _26688_ (.A(cpuregs[7][25]), .B(_00008_[2]), .Y(_05893_));
NAND_g _26689_ (.A(cpuregs[3][25]), .B(_09032_), .Y(_05894_));
NAND_g _26690_ (.A(_05893_), .B(_05894_), .Y(_05895_));
NAND_g _26691_ (.A(_00008_[0]), .B(_05895_), .Y(_05896_));
NAND_g _26692_ (.A(cpuregs[6][25]), .B(_00008_[2]), .Y(_05897_));
NAND_g _26693_ (.A(cpuregs[2][25]), .B(_09032_), .Y(_05898_));
NAND_g _26694_ (.A(_05897_), .B(_05898_), .Y(_05899_));
NAND_g _26695_ (.A(_09030_), .B(_05899_), .Y(_05900_));
AND_g _26696_ (.A(_05896_), .B(_05900_), .Y(_05901_));
NAND_g _26697_ (.A(cpuregs[4][25]), .B(_00008_[2]), .Y(_05902_));
NAND_g _26698_ (.A(cpuregs[0][25]), .B(_09032_), .Y(_05903_));
AND_g _26699_ (.A(_05902_), .B(_05903_), .Y(_05904_));
NAND_g _26700_ (.A(_09030_), .B(_05904_), .Y(_05905_));
NAND_g _26701_ (.A(cpuregs[5][25]), .B(_00008_[2]), .Y(_05906_));
NAND_g _26702_ (.A(cpuregs[1][25]), .B(_09032_), .Y(_05907_));
AND_g _26703_ (.A(_00008_[0]), .B(_05907_), .Y(_05908_));
NAND_g _26704_ (.A(_05906_), .B(_05908_), .Y(_05909_));
NAND_g _26705_ (.A(cpuregs[11][25]), .B(_09032_), .Y(_05910_));
NAND_g _26706_ (.A(cpuregs[15][25]), .B(_00008_[2]), .Y(_05911_));
NAND_g _26707_ (.A(_05910_), .B(_05911_), .Y(_05912_));
AND_g _26708_ (.A(_00008_[0]), .B(_05912_), .Y(_05913_));
NAND_g _26709_ (.A(cpuregs[14][25]), .B(_00008_[2]), .Y(_05914_));
NAND_g _26710_ (.A(cpuregs[10][25]), .B(_09032_), .Y(_05915_));
AND_g _26711_ (.A(_05914_), .B(_05915_), .Y(_05916_));
NOR_g _26712_ (.A(_00008_[0]), .B(_05916_), .Y(_05917_));
NOR_g _26713_ (.A(_05913_), .B(_05917_), .Y(_05918_));
NAND_g _26714_ (.A(_08883_), .B(_00008_[2]), .Y(_05919_));
NOR_g _26715_ (.A(cpuregs[8][25]), .B(_00008_[2]), .Y(_05920_));
NOR_g _26716_ (.A(_00008_[0]), .B(_05920_), .Y(_05921_));
NAND_g _26717_ (.A(_05919_), .B(_05921_), .Y(_05922_));
NAND_g _26718_ (.A(_08981_), .B(_09032_), .Y(_05923_));
NAND_g _26719_ (.A(_08933_), .B(_00008_[2]), .Y(_05924_));
AND_g _26720_ (.A(_00008_[0]), .B(_05924_), .Y(_05925_));
NAND_g _26721_ (.A(_05923_), .B(_05925_), .Y(_05926_));
NAND_g _26722_ (.A(_05922_), .B(_05926_), .Y(_05927_));
NAND_g _26723_ (.A(_00008_[3]), .B(_05927_), .Y(_05928_));
AND_g _26724_ (.A(_09033_), .B(_05909_), .Y(_05929_));
NAND_g _26725_ (.A(_05905_), .B(_05929_), .Y(_05930_));
NAND_g _26726_ (.A(_05928_), .B(_05930_), .Y(_05931_));
NAND_g _26727_ (.A(_09031_), .B(_05931_), .Y(_05932_));
NAND_g _26728_ (.A(_00008_[3]), .B(_05918_), .Y(_05933_));
NAND_g _26729_ (.A(_09033_), .B(_05901_), .Y(_05934_));
AND_g _26730_ (.A(_05933_), .B(_05934_), .Y(_05935_));
AND_g _26731_ (.A(_00008_[1]), .B(_05935_), .Y(_05936_));
NOR_g _26732_ (.A(_00008_[4]), .B(_05936_), .Y(_05937_));
NAND_g _26733_ (.A(_05932_), .B(_05937_), .Y(_05938_));
NAND_g _26734_ (.A(_08900_), .B(_00008_[2]), .Y(_05939_));
NOR_g _26735_ (.A(cpuregs[19][25]), .B(_00008_[2]), .Y(_05940_));
NOR_g _26736_ (.A(cpuregs[18][25]), .B(_00008_[2]), .Y(_05941_));
AND_g _26737_ (.A(_08925_), .B(_00008_[2]), .Y(_05942_));
NOR_g _26738_ (.A(_05941_), .B(_05942_), .Y(_05943_));
NOR_g _26739_ (.A(_09030_), .B(_05940_), .Y(_05944_));
NAND_g _26740_ (.A(_05939_), .B(_05944_), .Y(_05945_));
NAND_g _26741_ (.A(_09030_), .B(_05943_), .Y(_05946_));
AND_g _26742_ (.A(_05945_), .B(_05946_), .Y(_05947_));
NAND_g _26743_ (.A(_00008_[1]), .B(_05947_), .Y(_05948_));
NOR_g _26744_ (.A(cpuregs[17][25]), .B(_00008_[2]), .Y(_05949_));
NAND_g _26745_ (.A(_08999_), .B(_00008_[2]), .Y(_05950_));
NOR_g _26746_ (.A(cpuregs[16][25]), .B(_00008_[2]), .Y(_05951_));
AND_g _26747_ (.A(_08851_), .B(_00008_[2]), .Y(_05952_));
NOR_g _26748_ (.A(_05951_), .B(_05952_), .Y(_05953_));
NOR_g _26749_ (.A(_09030_), .B(_05949_), .Y(_05954_));
NAND_g _26750_ (.A(_05950_), .B(_05954_), .Y(_05955_));
NAND_g _26751_ (.A(_09030_), .B(_05953_), .Y(_05956_));
AND_g _26752_ (.A(_05955_), .B(_05956_), .Y(_05957_));
NAND_g _26753_ (.A(_09031_), .B(_05957_), .Y(_05958_));
NAND_g _26754_ (.A(_05948_), .B(_05958_), .Y(_05959_));
NAND_g _26755_ (.A(_09033_), .B(_05959_), .Y(_05960_));
NAND_g _26756_ (.A(cpuregs[25][25]), .B(_09031_), .Y(_05961_));
NAND_g _26757_ (.A(cpuregs[27][25]), .B(_00008_[1]), .Y(_05962_));
AND_g _26758_ (.A(_09032_), .B(_05962_), .Y(_05963_));
NAND_g _26759_ (.A(_05961_), .B(_05963_), .Y(_05964_));
NAND_g _26760_ (.A(cpuregs[29][25]), .B(_09031_), .Y(_05965_));
NAND_g _26761_ (.A(cpuregs[31][25]), .B(_00008_[1]), .Y(_05966_));
AND_g _26762_ (.A(_00008_[2]), .B(_05966_), .Y(_05967_));
NAND_g _26763_ (.A(_05965_), .B(_05967_), .Y(_05968_));
NAND_g _26764_ (.A(_05964_), .B(_05968_), .Y(_05969_));
NAND_g _26765_ (.A(_00008_[0]), .B(_05969_), .Y(_05970_));
NAND_g _26766_ (.A(cpuregs[24][25]), .B(_09031_), .Y(_05971_));
NAND_g _26767_ (.A(cpuregs[26][25]), .B(_00008_[1]), .Y(_05972_));
AND_g _26768_ (.A(_09032_), .B(_05972_), .Y(_05973_));
NAND_g _26769_ (.A(_05971_), .B(_05973_), .Y(_05974_));
NAND_g _26770_ (.A(cpuregs[28][25]), .B(_09031_), .Y(_05975_));
NAND_g _26771_ (.A(cpuregs[30][25]), .B(_00008_[1]), .Y(_05976_));
AND_g _26772_ (.A(_00008_[2]), .B(_05976_), .Y(_05977_));
NAND_g _26773_ (.A(_05975_), .B(_05977_), .Y(_05978_));
NAND_g _26774_ (.A(_05974_), .B(_05978_), .Y(_05979_));
NAND_g _26775_ (.A(_09030_), .B(_05979_), .Y(_05980_));
NAND_g _26776_ (.A(_05970_), .B(_05980_), .Y(_05981_));
NAND_g _26777_ (.A(_00008_[3]), .B(_05981_), .Y(_05982_));
NAND_g _26778_ (.A(_05960_), .B(_05982_), .Y(_05983_));
NAND_g _26779_ (.A(_00008_[4]), .B(_05983_), .Y(_05984_));
AND_g _26780_ (.A(_14624_), .B(_05938_), .Y(_05985_));
NAND_g _26781_ (.A(_05984_), .B(_05985_), .Y(_05986_));
NAND_g _26782_ (.A(_05892_), .B(_05986_), .Y(_05987_));
NAND_g _26783_ (.A(_10595_), .B(_05987_), .Y(_05988_));
NAND_g _26784_ (.A(pcpi_rs1[24]), .B(_14481_), .Y(_05989_));
AND_g _26785_ (.A(_05653_), .B(_05989_), .Y(_05990_));
NAND_g _26786_ (.A(pcpi_rs1[29]), .B(_14482_), .Y(_05991_));
AND_g _26787_ (.A(_05651_), .B(_05991_), .Y(_05992_));
NAND_g _26788_ (.A(_13880_), .B(_05992_), .Y(_05993_));
NAND_g _26789_ (.A(_13879_), .B(_05990_), .Y(_05994_));
AND_g _26790_ (.A(_13883_), .B(_05993_), .Y(_05995_));
NAND_g _26791_ (.A(_05994_), .B(_05995_), .Y(_05996_));
AND_g _26792_ (.A(_14488_), .B(_05996_), .Y(_05997_));
AND_g _26793_ (.A(_05988_), .B(_05997_), .Y(_05998_));
AND_g _26794_ (.A(_05891_), .B(_05998_), .Y(_05999_));
NOR_g _26795_ (.A(_05888_), .B(_05999_), .Y(_01043_));
NOR_g _26796_ (.A(pcpi_rs1[26]), .B(_14488_), .Y(_06000_));
XOR_g _26797_ (.A(_14500_), .B(_14602_), .Y(_06001_));
NAND_g _26798_ (.A(_14614_), .B(_06001_), .Y(_06002_));
NAND_g _26799_ (.A(reg_pc[26]), .B(_14617_), .Y(_06003_));
NAND_g _26800_ (.A(cpuregs[7][26]), .B(_00008_[2]), .Y(_06004_));
NAND_g _26801_ (.A(cpuregs[3][26]), .B(_09032_), .Y(_06005_));
NAND_g _26802_ (.A(_06004_), .B(_06005_), .Y(_06006_));
AND_g _26803_ (.A(_00008_[0]), .B(_06006_), .Y(_06007_));
NAND_g _26804_ (.A(cpuregs[6][26]), .B(_00008_[2]), .Y(_06008_));
NAND_g _26805_ (.A(cpuregs[2][26]), .B(_09032_), .Y(_06009_));
AND_g _26806_ (.A(_06008_), .B(_06009_), .Y(_06010_));
NOR_g _26807_ (.A(_00008_[0]), .B(_06010_), .Y(_06011_));
NOR_g _26808_ (.A(_06007_), .B(_06011_), .Y(_06012_));
NAND_g _26809_ (.A(cpuregs[5][26]), .B(_00008_[2]), .Y(_06013_));
NAND_g _26810_ (.A(cpuregs[1][26]), .B(_09032_), .Y(_06014_));
NAND_g _26811_ (.A(_06013_), .B(_06014_), .Y(_06015_));
NAND_g _26812_ (.A(_00008_[0]), .B(_06015_), .Y(_06016_));
NAND_g _26813_ (.A(cpuregs[4][26]), .B(_00008_[2]), .Y(_06017_));
NAND_g _26814_ (.A(cpuregs[0][26]), .B(_09032_), .Y(_06018_));
AND_g _26815_ (.A(_06017_), .B(_06018_), .Y(_06019_));
NOR_g _26816_ (.A(_00008_[0]), .B(_06019_), .Y(_06020_));
NAND_g _26817_ (.A(_00008_[1]), .B(_06012_), .Y(_06021_));
NOR_g _26818_ (.A(_00008_[1]), .B(_06020_), .Y(_06022_));
NAND_g _26819_ (.A(_06016_), .B(_06022_), .Y(_06023_));
AND_g _26820_ (.A(_09033_), .B(_06023_), .Y(_06024_));
NAND_g _26821_ (.A(_06021_), .B(_06024_), .Y(_06025_));
NAND_g _26822_ (.A(cpuregs[13][26]), .B(_00008_[0]), .Y(_06026_));
NAND_g _26823_ (.A(cpuregs[12][26]), .B(_09030_), .Y(_06027_));
AND_g _26824_ (.A(_00008_[2]), .B(_06027_), .Y(_06028_));
NAND_g _26825_ (.A(_06026_), .B(_06028_), .Y(_06029_));
NAND_g _26826_ (.A(cpuregs[9][26]), .B(_00008_[0]), .Y(_06030_));
NAND_g _26827_ (.A(cpuregs[8][26]), .B(_09030_), .Y(_06031_));
AND_g _26828_ (.A(_09032_), .B(_06031_), .Y(_06032_));
NAND_g _26829_ (.A(_06030_), .B(_06032_), .Y(_06033_));
AND_g _26830_ (.A(_09031_), .B(_06033_), .Y(_06034_));
NAND_g _26831_ (.A(_06029_), .B(_06034_), .Y(_06035_));
NAND_g _26832_ (.A(cpuregs[15][26]), .B(_00008_[0]), .Y(_06036_));
NAND_g _26833_ (.A(cpuregs[14][26]), .B(_09030_), .Y(_06037_));
AND_g _26834_ (.A(_00008_[2]), .B(_06037_), .Y(_06038_));
NAND_g _26835_ (.A(_06036_), .B(_06038_), .Y(_06039_));
NAND_g _26836_ (.A(cpuregs[11][26]), .B(_00008_[0]), .Y(_06040_));
NAND_g _26837_ (.A(cpuregs[10][26]), .B(_09030_), .Y(_06041_));
AND_g _26838_ (.A(_09032_), .B(_06041_), .Y(_06042_));
NAND_g _26839_ (.A(_06040_), .B(_06042_), .Y(_06043_));
AND_g _26840_ (.A(_00008_[1]), .B(_06043_), .Y(_06044_));
NAND_g _26841_ (.A(_06039_), .B(_06044_), .Y(_06045_));
NAND_g _26842_ (.A(_06035_), .B(_06045_), .Y(_06046_));
AND_g _26843_ (.A(_00008_[3]), .B(_06046_), .Y(_06047_));
NOR_g _26844_ (.A(_00008_[4]), .B(_06047_), .Y(_06048_));
NAND_g _26845_ (.A(_06025_), .B(_06048_), .Y(_06049_));
NAND_g _26846_ (.A(cpuregs[25][26]), .B(_09032_), .Y(_06050_));
NAND_g _26847_ (.A(cpuregs[29][26]), .B(_00008_[2]), .Y(_06051_));
AND_g _26848_ (.A(_09031_), .B(_06051_), .Y(_06052_));
NAND_g _26849_ (.A(_06050_), .B(_06052_), .Y(_06053_));
NAND_g _26850_ (.A(cpuregs[31][26]), .B(_00008_[2]), .Y(_06054_));
NAND_g _26851_ (.A(cpuregs[27][26]), .B(_09032_), .Y(_06055_));
AND_g _26852_ (.A(_00008_[1]), .B(_06055_), .Y(_06056_));
NAND_g _26853_ (.A(_06054_), .B(_06056_), .Y(_06057_));
NAND_g _26854_ (.A(_06053_), .B(_06057_), .Y(_06058_));
NAND_g _26855_ (.A(_00008_[0]), .B(_06058_), .Y(_06059_));
NAND_g _26856_ (.A(cpuregs[24][26]), .B(_09032_), .Y(_06060_));
NAND_g _26857_ (.A(cpuregs[28][26]), .B(_00008_[2]), .Y(_06061_));
AND_g _26858_ (.A(_09031_), .B(_06061_), .Y(_06062_));
NAND_g _26859_ (.A(_06060_), .B(_06062_), .Y(_06063_));
NAND_g _26860_ (.A(cpuregs[26][26]), .B(_09032_), .Y(_06064_));
NAND_g _26861_ (.A(cpuregs[30][26]), .B(_00008_[2]), .Y(_06065_));
AND_g _26862_ (.A(_00008_[1]), .B(_06065_), .Y(_06066_));
NAND_g _26863_ (.A(_06064_), .B(_06066_), .Y(_06067_));
NAND_g _26864_ (.A(_06063_), .B(_06067_), .Y(_06068_));
NAND_g _26865_ (.A(_09030_), .B(_06068_), .Y(_06069_));
NAND_g _26866_ (.A(_06059_), .B(_06069_), .Y(_06070_));
NAND_g _26867_ (.A(_00008_[3]), .B(_06070_), .Y(_06071_));
NAND_g _26868_ (.A(cpuregs[17][26]), .B(_09031_), .Y(_06072_));
NAND_g _26869_ (.A(cpuregs[19][26]), .B(_00008_[1]), .Y(_06073_));
AND_g _26870_ (.A(_09032_), .B(_06073_), .Y(_06074_));
NAND_g _26871_ (.A(_06072_), .B(_06074_), .Y(_06075_));
NAND_g _26872_ (.A(cpuregs[21][26]), .B(_09031_), .Y(_06076_));
NAND_g _26873_ (.A(cpuregs[23][26]), .B(_00008_[1]), .Y(_06077_));
AND_g _26874_ (.A(_00008_[2]), .B(_06077_), .Y(_06078_));
NAND_g _26875_ (.A(_06076_), .B(_06078_), .Y(_06079_));
NAND_g _26876_ (.A(_06075_), .B(_06079_), .Y(_06080_));
NAND_g _26877_ (.A(_00008_[0]), .B(_06080_), .Y(_06081_));
NAND_g _26878_ (.A(cpuregs[16][26]), .B(_09031_), .Y(_06082_));
NAND_g _26879_ (.A(cpuregs[18][26]), .B(_00008_[1]), .Y(_06083_));
AND_g _26880_ (.A(_09032_), .B(_06083_), .Y(_06084_));
NAND_g _26881_ (.A(_06082_), .B(_06084_), .Y(_06085_));
NAND_g _26882_ (.A(cpuregs[20][26]), .B(_09031_), .Y(_06086_));
NAND_g _26883_ (.A(cpuregs[22][26]), .B(_00008_[1]), .Y(_06087_));
AND_g _26884_ (.A(_00008_[2]), .B(_06087_), .Y(_06088_));
NAND_g _26885_ (.A(_06086_), .B(_06088_), .Y(_06089_));
NAND_g _26886_ (.A(_06085_), .B(_06089_), .Y(_06090_));
NAND_g _26887_ (.A(_09030_), .B(_06090_), .Y(_06091_));
NAND_g _26888_ (.A(_06081_), .B(_06091_), .Y(_06092_));
AND_g _26889_ (.A(_09033_), .B(_06092_), .Y(_06093_));
NOT_g _26890_ (.A(_06093_), .Y(_06094_));
NAND_g _26891_ (.A(_06071_), .B(_06094_), .Y(_06095_));
NAND_g _26892_ (.A(_00008_[4]), .B(_06095_), .Y(_06096_));
AND_g _26893_ (.A(_14624_), .B(_06096_), .Y(_06097_));
NAND_g _26894_ (.A(_06049_), .B(_06097_), .Y(_06098_));
NAND_g _26895_ (.A(_06003_), .B(_06098_), .Y(_06099_));
NAND_g _26896_ (.A(_10595_), .B(_06099_), .Y(_06100_));
NAND_g _26897_ (.A(pcpi_rs1[25]), .B(_14481_), .Y(_06101_));
AND_g _26898_ (.A(_05764_), .B(_06101_), .Y(_06102_));
NAND_g _26899_ (.A(pcpi_rs1[30]), .B(_14482_), .Y(_06103_));
AND_g _26900_ (.A(_05762_), .B(_06103_), .Y(_06104_));
NAND_g _26901_ (.A(_13880_), .B(_06104_), .Y(_06105_));
NAND_g _26902_ (.A(_13879_), .B(_06102_), .Y(_06106_));
AND_g _26903_ (.A(_13883_), .B(_06105_), .Y(_06107_));
NAND_g _26904_ (.A(_06106_), .B(_06107_), .Y(_06108_));
AND_g _26905_ (.A(_14488_), .B(_06108_), .Y(_06109_));
AND_g _26906_ (.A(_06100_), .B(_06109_), .Y(_06110_));
AND_g _26907_ (.A(_06002_), .B(_06110_), .Y(_06111_));
NOR_g _26908_ (.A(_06000_), .B(_06111_), .Y(_01044_));
NOR_g _26909_ (.A(pcpi_rs1[27]), .B(_14488_), .Y(_06112_));
XNOR_g _26910_ (.A(decoded_imm[27]), .B(pcpi_rs1[27]), .Y(_06113_));
NOR_g _26911_ (.A(_14604_), .B(_06113_), .Y(_06114_));
NAND_g _26912_ (.A(_14604_), .B(_06113_), .Y(_06115_));
NAND_g _26913_ (.A(_14614_), .B(_06115_), .Y(_06116_));
NOR_g _26914_ (.A(_06114_), .B(_06116_), .Y(_06117_));
NAND_g _26915_ (.A(reg_pc[27]), .B(_14617_), .Y(_06118_));
NAND_g _26916_ (.A(_08978_), .B(_00008_[2]), .Y(_06119_));
NOR_g _26917_ (.A(cpuregs[3][27]), .B(_00008_[2]), .Y(_06120_));
NOR_g _26918_ (.A(_09030_), .B(_06120_), .Y(_06121_));
AND_g _26919_ (.A(_06119_), .B(_06121_), .Y(_06122_));
NAND_g _26920_ (.A(cpuregs[6][27]), .B(_00008_[2]), .Y(_06123_));
NAND_g _26921_ (.A(cpuregs[2][27]), .B(_09032_), .Y(_06124_));
AND_g _26922_ (.A(_06123_), .B(_06124_), .Y(_06125_));
NOR_g _26923_ (.A(_00008_[0]), .B(_06125_), .Y(_06126_));
NOR_g _26924_ (.A(_06122_), .B(_06126_), .Y(_06127_));
NAND_g _26925_ (.A(cpuregs[5][27]), .B(_00008_[2]), .Y(_06128_));
NAND_g _26926_ (.A(cpuregs[1][27]), .B(_09032_), .Y(_06129_));
NAND_g _26927_ (.A(_06128_), .B(_06129_), .Y(_06130_));
NAND_g _26928_ (.A(_00008_[0]), .B(_06130_), .Y(_06131_));
NAND_g _26929_ (.A(cpuregs[4][27]), .B(_00008_[2]), .Y(_06132_));
NAND_g _26930_ (.A(cpuregs[0][27]), .B(_09032_), .Y(_06133_));
AND_g _26931_ (.A(_06132_), .B(_06133_), .Y(_06134_));
NOR_g _26932_ (.A(_00008_[0]), .B(_06134_), .Y(_06135_));
NAND_g _26933_ (.A(_00008_[1]), .B(_06127_), .Y(_06136_));
NOR_g _26934_ (.A(_00008_[1]), .B(_06135_), .Y(_06137_));
NAND_g _26935_ (.A(_06131_), .B(_06137_), .Y(_06138_));
AND_g _26936_ (.A(_06136_), .B(_06138_), .Y(_06139_));
NAND_g _26937_ (.A(_09033_), .B(_06139_), .Y(_06140_));
NAND_g _26938_ (.A(cpuregs[13][27]), .B(_00008_[0]), .Y(_06141_));
NAND_g _26939_ (.A(cpuregs[12][27]), .B(_09030_), .Y(_06142_));
AND_g _26940_ (.A(_00008_[2]), .B(_06142_), .Y(_06143_));
NAND_g _26941_ (.A(_06141_), .B(_06143_), .Y(_06144_));
NAND_g _26942_ (.A(cpuregs[9][27]), .B(_00008_[0]), .Y(_06145_));
NAND_g _26943_ (.A(cpuregs[8][27]), .B(_09030_), .Y(_06146_));
AND_g _26944_ (.A(_09032_), .B(_06146_), .Y(_06147_));
NAND_g _26945_ (.A(_06145_), .B(_06147_), .Y(_06148_));
AND_g _26946_ (.A(_09031_), .B(_06148_), .Y(_06149_));
NAND_g _26947_ (.A(_06144_), .B(_06149_), .Y(_06150_));
NAND_g _26948_ (.A(cpuregs[15][27]), .B(_00008_[0]), .Y(_06151_));
NAND_g _26949_ (.A(cpuregs[14][27]), .B(_09030_), .Y(_06152_));
AND_g _26950_ (.A(_00008_[2]), .B(_06152_), .Y(_06153_));
NAND_g _26951_ (.A(_06151_), .B(_06153_), .Y(_06154_));
NAND_g _26952_ (.A(cpuregs[11][27]), .B(_00008_[0]), .Y(_06155_));
NAND_g _26953_ (.A(cpuregs[10][27]), .B(_09030_), .Y(_06156_));
AND_g _26954_ (.A(_09032_), .B(_06156_), .Y(_06157_));
NAND_g _26955_ (.A(_06155_), .B(_06157_), .Y(_06158_));
AND_g _26956_ (.A(_00008_[1]), .B(_06158_), .Y(_06159_));
NAND_g _26957_ (.A(_06154_), .B(_06159_), .Y(_06160_));
NAND_g _26958_ (.A(_06150_), .B(_06160_), .Y(_06161_));
AND_g _26959_ (.A(_00008_[3]), .B(_06161_), .Y(_06162_));
NOR_g _26960_ (.A(_00008_[4]), .B(_06162_), .Y(_06163_));
NAND_g _26961_ (.A(_06140_), .B(_06163_), .Y(_06164_));
NAND_g _26962_ (.A(cpuregs[26][27]), .B(_09032_), .Y(_06165_));
NAND_g _26963_ (.A(cpuregs[30][27]), .B(_00008_[2]), .Y(_06166_));
AND_g _26964_ (.A(_09030_), .B(_06166_), .Y(_06167_));
NAND_g _26965_ (.A(_06165_), .B(_06167_), .Y(_06168_));
NAND_g _26966_ (.A(cpuregs[31][27]), .B(_00008_[2]), .Y(_06169_));
NAND_g _26967_ (.A(cpuregs[27][27]), .B(_09032_), .Y(_06170_));
AND_g _26968_ (.A(_00008_[0]), .B(_06170_), .Y(_06171_));
NAND_g _26969_ (.A(_06169_), .B(_06171_), .Y(_06172_));
NAND_g _26970_ (.A(_06168_), .B(_06172_), .Y(_06173_));
NAND_g _26971_ (.A(_00008_[3]), .B(_06173_), .Y(_06174_));
NAND_g _26972_ (.A(cpuregs[18][27]), .B(_09032_), .Y(_06175_));
NAND_g _26973_ (.A(cpuregs[22][27]), .B(_00008_[2]), .Y(_06176_));
AND_g _26974_ (.A(_09030_), .B(_06176_), .Y(_06177_));
NAND_g _26975_ (.A(_06175_), .B(_06177_), .Y(_06178_));
NAND_g _26976_ (.A(cpuregs[19][27]), .B(_09032_), .Y(_06179_));
NAND_g _26977_ (.A(cpuregs[23][27]), .B(_00008_[2]), .Y(_06180_));
AND_g _26978_ (.A(_00008_[0]), .B(_06180_), .Y(_06181_));
NAND_g _26979_ (.A(_06179_), .B(_06181_), .Y(_06182_));
NAND_g _26980_ (.A(_06178_), .B(_06182_), .Y(_06183_));
NAND_g _26981_ (.A(_09033_), .B(_06183_), .Y(_06184_));
AND_g _26982_ (.A(_06174_), .B(_06184_), .Y(_06185_));
NAND_g _26983_ (.A(cpuregs[24][27]), .B(_09032_), .Y(_06186_));
NAND_g _26984_ (.A(cpuregs[28][27]), .B(_00008_[2]), .Y(_06187_));
AND_g _26985_ (.A(_09030_), .B(_06187_), .Y(_06188_));
NAND_g _26986_ (.A(_06186_), .B(_06188_), .Y(_06189_));
NAND_g _26987_ (.A(cpuregs[29][27]), .B(_00008_[2]), .Y(_06190_));
NAND_g _26988_ (.A(cpuregs[25][27]), .B(_09032_), .Y(_06191_));
AND_g _26989_ (.A(_00008_[0]), .B(_06191_), .Y(_06192_));
NAND_g _26990_ (.A(_06190_), .B(_06192_), .Y(_06193_));
NAND_g _26991_ (.A(_06189_), .B(_06193_), .Y(_06194_));
NAND_g _26992_ (.A(_00008_[3]), .B(_06194_), .Y(_06195_));
NAND_g _26993_ (.A(cpuregs[16][27]), .B(_09032_), .Y(_06196_));
NAND_g _26994_ (.A(cpuregs[20][27]), .B(_00008_[2]), .Y(_06197_));
AND_g _26995_ (.A(_09030_), .B(_06197_), .Y(_06198_));
NAND_g _26996_ (.A(_06196_), .B(_06198_), .Y(_06199_));
NAND_g _26997_ (.A(cpuregs[17][27]), .B(_09032_), .Y(_06200_));
NAND_g _26998_ (.A(cpuregs[21][27]), .B(_00008_[2]), .Y(_06201_));
AND_g _26999_ (.A(_00008_[0]), .B(_06201_), .Y(_06202_));
NAND_g _27000_ (.A(_06200_), .B(_06202_), .Y(_06203_));
NAND_g _27001_ (.A(_06199_), .B(_06203_), .Y(_06204_));
NAND_g _27002_ (.A(_09033_), .B(_06204_), .Y(_06205_));
AND_g _27003_ (.A(_06195_), .B(_06205_), .Y(_06206_));
NAND_g _27004_ (.A(_00008_[1]), .B(_06185_), .Y(_06207_));
NAND_g _27005_ (.A(_09031_), .B(_06206_), .Y(_06208_));
AND_g _27006_ (.A(_00008_[4]), .B(_06207_), .Y(_06209_));
NAND_g _27007_ (.A(_06208_), .B(_06209_), .Y(_06210_));
AND_g _27008_ (.A(_14624_), .B(_06210_), .Y(_06211_));
NAND_g _27009_ (.A(_06164_), .B(_06211_), .Y(_06212_));
NAND_g _27010_ (.A(_06118_), .B(_06212_), .Y(_06213_));
NAND_g _27011_ (.A(_10595_), .B(_06213_), .Y(_06214_));
NAND_g _27012_ (.A(pcpi_rs1[26]), .B(_14481_), .Y(_06215_));
AND_g _27013_ (.A(_05879_), .B(_06215_), .Y(_06216_));
NAND_g _27014_ (.A(pcpi_rs1[31]), .B(_14482_), .Y(_06217_));
AND_g _27015_ (.A(_05877_), .B(_06217_), .Y(_06218_));
NAND_g _27016_ (.A(_13880_), .B(_06218_), .Y(_06219_));
NAND_g _27017_ (.A(_13879_), .B(_06216_), .Y(_06220_));
AND_g _27018_ (.A(_13883_), .B(_06219_), .Y(_06221_));
NAND_g _27019_ (.A(_06220_), .B(_06221_), .Y(_06222_));
AND_g _27020_ (.A(_14488_), .B(_06222_), .Y(_06223_));
NAND_g _27021_ (.A(_06214_), .B(_06223_), .Y(_06224_));
NOR_g _27022_ (.A(_06117_), .B(_06224_), .Y(_06225_));
NOR_g _27023_ (.A(_06112_), .B(_06225_), .Y(_01045_));
NOR_g _27024_ (.A(pcpi_rs1[28]), .B(_14488_), .Y(_06226_));
XOR_g _27025_ (.A(_14496_), .B(_14606_), .Y(_06227_));
NAND_g _27026_ (.A(_14614_), .B(_06227_), .Y(_06228_));
NAND_g _27027_ (.A(reg_pc[28]), .B(_14617_), .Y(_06229_));
NAND_g _27028_ (.A(cpuregs[13][28]), .B(_00008_[2]), .Y(_06230_));
NAND_g _27029_ (.A(cpuregs[9][28]), .B(_09032_), .Y(_06231_));
NAND_g _27030_ (.A(_06230_), .B(_06231_), .Y(_06232_));
NAND_g _27031_ (.A(_00008_[0]), .B(_06232_), .Y(_06233_));
NAND_g _27032_ (.A(cpuregs[12][28]), .B(_00008_[2]), .Y(_06234_));
NAND_g _27033_ (.A(cpuregs[8][28]), .B(_09032_), .Y(_06235_));
AND_g _27034_ (.A(_06234_), .B(_06235_), .Y(_06236_));
NOR_g _27035_ (.A(_00008_[0]), .B(_06236_), .Y(_06237_));
NAND_g _27036_ (.A(_08917_), .B(_00008_[2]), .Y(_06238_));
NOR_g _27037_ (.A(cpuregs[0][28]), .B(_00008_[2]), .Y(_06239_));
NOR_g _27038_ (.A(_00008_[0]), .B(_06239_), .Y(_06240_));
NAND_g _27039_ (.A(_06238_), .B(_06240_), .Y(_06241_));
NAND_g _27040_ (.A(_08960_), .B(_00008_[2]), .Y(_06242_));
NOR_g _27041_ (.A(cpuregs[1][28]), .B(_00008_[2]), .Y(_06243_));
NOR_g _27042_ (.A(_09030_), .B(_06243_), .Y(_06244_));
NAND_g _27043_ (.A(_06242_), .B(_06244_), .Y(_06245_));
NAND_g _27044_ (.A(cpuregs[11][28]), .B(_09032_), .Y(_06246_));
NAND_g _27045_ (.A(cpuregs[15][28]), .B(_00008_[2]), .Y(_06247_));
NAND_g _27046_ (.A(_06246_), .B(_06247_), .Y(_06248_));
AND_g _27047_ (.A(_00008_[0]), .B(_06248_), .Y(_06249_));
NAND_g _27048_ (.A(cpuregs[14][28]), .B(_00008_[2]), .Y(_06250_));
NAND_g _27049_ (.A(cpuregs[10][28]), .B(_09032_), .Y(_06251_));
AND_g _27050_ (.A(_06250_), .B(_06251_), .Y(_06252_));
NOR_g _27051_ (.A(_00008_[0]), .B(_06252_), .Y(_06253_));
NOR_g _27052_ (.A(_06249_), .B(_06253_), .Y(_06254_));
NAND_g _27053_ (.A(_09016_), .B(_00008_[2]), .Y(_06255_));
NOR_g _27054_ (.A(cpuregs[2][28]), .B(_00008_[2]), .Y(_06256_));
NOR_g _27055_ (.A(_00008_[0]), .B(_06256_), .Y(_06257_));
NAND_g _27056_ (.A(_06255_), .B(_06257_), .Y(_06258_));
NAND_g _27057_ (.A(_08979_), .B(_00008_[2]), .Y(_06259_));
NOR_g _27058_ (.A(cpuregs[3][28]), .B(_00008_[2]), .Y(_06260_));
NOR_g _27059_ (.A(_09030_), .B(_06260_), .Y(_06261_));
NAND_g _27060_ (.A(_06259_), .B(_06261_), .Y(_06262_));
AND_g _27061_ (.A(_06258_), .B(_06262_), .Y(_06263_));
AND_g _27062_ (.A(_09031_), .B(_06241_), .Y(_06264_));
NAND_g _27063_ (.A(_06245_), .B(_06264_), .Y(_06265_));
NAND_g _27064_ (.A(_00008_[1]), .B(_06263_), .Y(_06266_));
AND_g _27065_ (.A(_06265_), .B(_06266_), .Y(_06267_));
NAND_g _27066_ (.A(_09033_), .B(_06267_), .Y(_06268_));
NAND_g _27067_ (.A(_00008_[1]), .B(_06254_), .Y(_06269_));
NOR_g _27068_ (.A(_00008_[1]), .B(_06237_), .Y(_06270_));
NAND_g _27069_ (.A(_06233_), .B(_06270_), .Y(_06271_));
AND_g _27070_ (.A(_00008_[3]), .B(_06271_), .Y(_06272_));
AND_g _27071_ (.A(_06269_), .B(_06272_), .Y(_06273_));
NOR_g _27072_ (.A(_00008_[4]), .B(_06273_), .Y(_06274_));
NAND_g _27073_ (.A(_06268_), .B(_06274_), .Y(_06275_));
NAND_g _27074_ (.A(_08902_), .B(_00008_[2]), .Y(_06276_));
NOR_g _27075_ (.A(cpuregs[19][28]), .B(_00008_[2]), .Y(_06277_));
NOR_g _27076_ (.A(cpuregs[18][28]), .B(_00008_[2]), .Y(_06278_));
NOR_g _27077_ (.A(cpuregs[22][28]), .B(_09032_), .Y(_06279_));
NOR_g _27078_ (.A(_06278_), .B(_06279_), .Y(_06280_));
NOR_g _27079_ (.A(_09030_), .B(_06277_), .Y(_06281_));
NAND_g _27080_ (.A(_06276_), .B(_06281_), .Y(_06282_));
NAND_g _27081_ (.A(_09030_), .B(_06280_), .Y(_06283_));
AND_g _27082_ (.A(_06282_), .B(_06283_), .Y(_06284_));
NAND_g _27083_ (.A(_00008_[1]), .B(_06284_), .Y(_06285_));
NOR_g _27084_ (.A(cpuregs[17][28]), .B(_00008_[2]), .Y(_06286_));
NAND_g _27085_ (.A(_09001_), .B(_00008_[2]), .Y(_06287_));
NOR_g _27086_ (.A(cpuregs[16][28]), .B(_00008_[2]), .Y(_06288_));
NOR_g _27087_ (.A(cpuregs[20][28]), .B(_09032_), .Y(_06289_));
NOR_g _27088_ (.A(_06288_), .B(_06289_), .Y(_06290_));
NOR_g _27089_ (.A(_09030_), .B(_06286_), .Y(_06291_));
NAND_g _27090_ (.A(_06287_), .B(_06291_), .Y(_06292_));
NAND_g _27091_ (.A(_09030_), .B(_06290_), .Y(_06293_));
AND_g _27092_ (.A(_06292_), .B(_06293_), .Y(_06294_));
NAND_g _27093_ (.A(_09031_), .B(_06294_), .Y(_06295_));
NAND_g _27094_ (.A(_06285_), .B(_06295_), .Y(_06296_));
NAND_g _27095_ (.A(_09033_), .B(_06296_), .Y(_06297_));
NAND_g _27096_ (.A(cpuregs[25][28]), .B(_09031_), .Y(_06298_));
NAND_g _27097_ (.A(cpuregs[27][28]), .B(_00008_[1]), .Y(_06299_));
AND_g _27098_ (.A(_09032_), .B(_06299_), .Y(_06300_));
NAND_g _27099_ (.A(_06298_), .B(_06300_), .Y(_06301_));
NAND_g _27100_ (.A(cpuregs[29][28]), .B(_09031_), .Y(_06302_));
NAND_g _27101_ (.A(cpuregs[31][28]), .B(_00008_[1]), .Y(_06303_));
AND_g _27102_ (.A(_00008_[2]), .B(_06303_), .Y(_06304_));
NAND_g _27103_ (.A(_06302_), .B(_06304_), .Y(_06305_));
NAND_g _27104_ (.A(_06301_), .B(_06305_), .Y(_06306_));
NAND_g _27105_ (.A(_00008_[0]), .B(_06306_), .Y(_06307_));
NAND_g _27106_ (.A(cpuregs[24][28]), .B(_09031_), .Y(_06308_));
NAND_g _27107_ (.A(cpuregs[26][28]), .B(_00008_[1]), .Y(_06309_));
AND_g _27108_ (.A(_09032_), .B(_06309_), .Y(_06310_));
NAND_g _27109_ (.A(_06308_), .B(_06310_), .Y(_06311_));
NAND_g _27110_ (.A(cpuregs[28][28]), .B(_09031_), .Y(_06312_));
NAND_g _27111_ (.A(cpuregs[30][28]), .B(_00008_[1]), .Y(_06313_));
AND_g _27112_ (.A(_00008_[2]), .B(_06313_), .Y(_06314_));
NAND_g _27113_ (.A(_06312_), .B(_06314_), .Y(_06315_));
NAND_g _27114_ (.A(_06311_), .B(_06315_), .Y(_06316_));
NAND_g _27115_ (.A(_09030_), .B(_06316_), .Y(_06317_));
NAND_g _27116_ (.A(_06307_), .B(_06317_), .Y(_06318_));
NAND_g _27117_ (.A(_00008_[3]), .B(_06318_), .Y(_06319_));
NAND_g _27118_ (.A(_06297_), .B(_06319_), .Y(_06320_));
NAND_g _27119_ (.A(_00008_[4]), .B(_06320_), .Y(_06321_));
AND_g _27120_ (.A(_14624_), .B(_06275_), .Y(_06322_));
NAND_g _27121_ (.A(_06321_), .B(_06322_), .Y(_06323_));
NAND_g _27122_ (.A(_06229_), .B(_06323_), .Y(_06324_));
NAND_g _27123_ (.A(_10595_), .B(_06324_), .Y(_06325_));
NOR_g _27124_ (.A(_13880_), .B(_14721_), .Y(_06326_));
NAND_g _27125_ (.A(_05991_), .B(_06326_), .Y(_06327_));
NAND_g _27126_ (.A(pcpi_rs1[31]), .B(_14477_), .Y(_06328_));
AND_g _27127_ (.A(_13880_), .B(_06328_), .Y(_06329_));
NAND_g _27128_ (.A(_05989_), .B(_06329_), .Y(_06330_));
AND_g _27129_ (.A(_06327_), .B(_06330_), .Y(_06331_));
NAND_g _27130_ (.A(_13883_), .B(_06331_), .Y(_06332_));
AND_g _27131_ (.A(_14488_), .B(_06325_), .Y(_06333_));
AND_g _27132_ (.A(_06332_), .B(_06333_), .Y(_06334_));
AND_g _27133_ (.A(_06228_), .B(_06334_), .Y(_06335_));
NOR_g _27134_ (.A(_06226_), .B(_06335_), .Y(_01046_));
NOR_g _27135_ (.A(pcpi_rs1[29]), .B(_14488_), .Y(_06336_));
XOR_g _27136_ (.A(decoded_imm[29]), .B(pcpi_rs1[29]), .Y(_06337_));
XNOR_g _27137_ (.A(_14608_), .B(_06337_), .Y(_06338_));
NAND_g _27138_ (.A(_14614_), .B(_06338_), .Y(_06339_));
NAND_g _27139_ (.A(reg_pc[29]), .B(_14617_), .Y(_06340_));
NAND_g _27140_ (.A(cpuregs[7][29]), .B(_00008_[2]), .Y(_06341_));
NAND_g _27141_ (.A(cpuregs[3][29]), .B(_09032_), .Y(_06342_));
NAND_g _27142_ (.A(_06341_), .B(_06342_), .Y(_06343_));
AND_g _27143_ (.A(_00008_[0]), .B(_06343_), .Y(_06344_));
NAND_g _27144_ (.A(cpuregs[6][29]), .B(_00008_[2]), .Y(_06345_));
NAND_g _27145_ (.A(cpuregs[2][29]), .B(_09032_), .Y(_06346_));
AND_g _27146_ (.A(_06345_), .B(_06346_), .Y(_06347_));
NOR_g _27147_ (.A(_00008_[0]), .B(_06347_), .Y(_06348_));
NOR_g _27148_ (.A(_06344_), .B(_06348_), .Y(_06349_));
NAND_g _27149_ (.A(cpuregs[5][29]), .B(_00008_[2]), .Y(_06350_));
NAND_g _27150_ (.A(cpuregs[1][29]), .B(_09032_), .Y(_06351_));
NAND_g _27151_ (.A(_06350_), .B(_06351_), .Y(_06352_));
NAND_g _27152_ (.A(_00008_[0]), .B(_06352_), .Y(_06353_));
NAND_g _27153_ (.A(cpuregs[4][29]), .B(_00008_[2]), .Y(_06354_));
NAND_g _27154_ (.A(cpuregs[0][29]), .B(_09032_), .Y(_06355_));
AND_g _27155_ (.A(_06354_), .B(_06355_), .Y(_06356_));
NOR_g _27156_ (.A(_00008_[0]), .B(_06356_), .Y(_06357_));
NAND_g _27157_ (.A(_00008_[1]), .B(_06349_), .Y(_06358_));
NOR_g _27158_ (.A(_00008_[1]), .B(_06357_), .Y(_06359_));
NAND_g _27159_ (.A(_06353_), .B(_06359_), .Y(_06360_));
AND_g _27160_ (.A(_09033_), .B(_06360_), .Y(_06361_));
NAND_g _27161_ (.A(_06358_), .B(_06361_), .Y(_06362_));
NAND_g _27162_ (.A(cpuregs[13][29]), .B(_00008_[0]), .Y(_06363_));
NAND_g _27163_ (.A(cpuregs[12][29]), .B(_09030_), .Y(_06364_));
AND_g _27164_ (.A(_00008_[2]), .B(_06364_), .Y(_06365_));
NAND_g _27165_ (.A(_06363_), .B(_06365_), .Y(_06366_));
NAND_g _27166_ (.A(cpuregs[9][29]), .B(_00008_[0]), .Y(_06367_));
NAND_g _27167_ (.A(cpuregs[8][29]), .B(_09030_), .Y(_06368_));
AND_g _27168_ (.A(_09032_), .B(_06368_), .Y(_06369_));
NAND_g _27169_ (.A(_06367_), .B(_06369_), .Y(_06370_));
AND_g _27170_ (.A(_09031_), .B(_06370_), .Y(_06371_));
NAND_g _27171_ (.A(_06366_), .B(_06371_), .Y(_06372_));
NAND_g _27172_ (.A(cpuregs[15][29]), .B(_00008_[0]), .Y(_06373_));
NAND_g _27173_ (.A(cpuregs[14][29]), .B(_09030_), .Y(_06374_));
AND_g _27174_ (.A(_00008_[2]), .B(_06374_), .Y(_06375_));
NAND_g _27175_ (.A(_06373_), .B(_06375_), .Y(_06376_));
NAND_g _27176_ (.A(cpuregs[11][29]), .B(_00008_[0]), .Y(_06377_));
NAND_g _27177_ (.A(cpuregs[10][29]), .B(_09030_), .Y(_06378_));
AND_g _27178_ (.A(_09032_), .B(_06378_), .Y(_06379_));
NAND_g _27179_ (.A(_06377_), .B(_06379_), .Y(_06380_));
AND_g _27180_ (.A(_00008_[1]), .B(_06380_), .Y(_06381_));
NAND_g _27181_ (.A(_06376_), .B(_06381_), .Y(_06382_));
NAND_g _27182_ (.A(_06372_), .B(_06382_), .Y(_06383_));
AND_g _27183_ (.A(_00008_[3]), .B(_06383_), .Y(_06384_));
NOR_g _27184_ (.A(_00008_[4]), .B(_06384_), .Y(_06385_));
NAND_g _27185_ (.A(_06362_), .B(_06385_), .Y(_06386_));
NAND_g _27186_ (.A(cpuregs[25][29]), .B(_09032_), .Y(_06387_));
NAND_g _27187_ (.A(cpuregs[29][29]), .B(_00008_[2]), .Y(_06388_));
AND_g _27188_ (.A(_09031_), .B(_06388_), .Y(_06389_));
NAND_g _27189_ (.A(_06387_), .B(_06389_), .Y(_06390_));
NAND_g _27190_ (.A(cpuregs[31][29]), .B(_00008_[2]), .Y(_06391_));
NAND_g _27191_ (.A(cpuregs[27][29]), .B(_09032_), .Y(_06392_));
AND_g _27192_ (.A(_00008_[1]), .B(_06392_), .Y(_06393_));
NAND_g _27193_ (.A(_06391_), .B(_06393_), .Y(_06394_));
NAND_g _27194_ (.A(_06390_), .B(_06394_), .Y(_06395_));
NAND_g _27195_ (.A(_00008_[0]), .B(_06395_), .Y(_06396_));
NAND_g _27196_ (.A(cpuregs[24][29]), .B(_09032_), .Y(_06397_));
NAND_g _27197_ (.A(cpuregs[28][29]), .B(_00008_[2]), .Y(_06398_));
AND_g _27198_ (.A(_09031_), .B(_06398_), .Y(_06399_));
NAND_g _27199_ (.A(_06397_), .B(_06399_), .Y(_06400_));
NAND_g _27200_ (.A(cpuregs[26][29]), .B(_09032_), .Y(_06401_));
NAND_g _27201_ (.A(cpuregs[30][29]), .B(_00008_[2]), .Y(_06402_));
AND_g _27202_ (.A(_00008_[1]), .B(_06402_), .Y(_06403_));
NAND_g _27203_ (.A(_06401_), .B(_06403_), .Y(_06404_));
NAND_g _27204_ (.A(_06400_), .B(_06404_), .Y(_06405_));
NAND_g _27205_ (.A(_09030_), .B(_06405_), .Y(_06406_));
NAND_g _27206_ (.A(_06396_), .B(_06406_), .Y(_06407_));
NAND_g _27207_ (.A(_00008_[3]), .B(_06407_), .Y(_06408_));
NAND_g _27208_ (.A(cpuregs[17][29]), .B(_09031_), .Y(_06409_));
NAND_g _27209_ (.A(cpuregs[19][29]), .B(_00008_[1]), .Y(_06410_));
AND_g _27210_ (.A(_09032_), .B(_06410_), .Y(_06411_));
NAND_g _27211_ (.A(_06409_), .B(_06411_), .Y(_06412_));
NAND_g _27212_ (.A(cpuregs[21][29]), .B(_09031_), .Y(_06413_));
NAND_g _27213_ (.A(cpuregs[23][29]), .B(_00008_[1]), .Y(_06414_));
AND_g _27214_ (.A(_00008_[2]), .B(_06414_), .Y(_06415_));
NAND_g _27215_ (.A(_06413_), .B(_06415_), .Y(_06416_));
NAND_g _27216_ (.A(_06412_), .B(_06416_), .Y(_06417_));
NAND_g _27217_ (.A(_00008_[0]), .B(_06417_), .Y(_06418_));
NAND_g _27218_ (.A(cpuregs[16][29]), .B(_09031_), .Y(_06419_));
NAND_g _27219_ (.A(cpuregs[18][29]), .B(_00008_[1]), .Y(_06420_));
AND_g _27220_ (.A(_09032_), .B(_06420_), .Y(_06421_));
NAND_g _27221_ (.A(_06419_), .B(_06421_), .Y(_06422_));
NAND_g _27222_ (.A(cpuregs[20][29]), .B(_09031_), .Y(_06423_));
NAND_g _27223_ (.A(cpuregs[22][29]), .B(_00008_[1]), .Y(_06424_));
AND_g _27224_ (.A(_00008_[2]), .B(_06424_), .Y(_06425_));
NAND_g _27225_ (.A(_06423_), .B(_06425_), .Y(_06426_));
NAND_g _27226_ (.A(_06422_), .B(_06426_), .Y(_06427_));
NAND_g _27227_ (.A(_09030_), .B(_06427_), .Y(_06428_));
NAND_g _27228_ (.A(_06418_), .B(_06428_), .Y(_06429_));
AND_g _27229_ (.A(_09033_), .B(_06429_), .Y(_06430_));
NOT_g _27230_ (.A(_06430_), .Y(_06431_));
NAND_g _27231_ (.A(_06408_), .B(_06431_), .Y(_06432_));
NAND_g _27232_ (.A(_00008_[4]), .B(_06432_), .Y(_06433_));
AND_g _27233_ (.A(_14624_), .B(_06433_), .Y(_06434_));
NAND_g _27234_ (.A(_06386_), .B(_06434_), .Y(_06435_));
NAND_g _27235_ (.A(_06340_), .B(_06435_), .Y(_06436_));
NAND_g _27236_ (.A(_10595_), .B(_06436_), .Y(_06437_));
NAND_g _27237_ (.A(pcpi_rs1[28]), .B(_14481_), .Y(_06438_));
AND_g _27238_ (.A(_13879_), .B(_06438_), .Y(_06439_));
NAND_g _27239_ (.A(_06103_), .B(_06439_), .Y(_06440_));
NAND_g _27240_ (.A(_06101_), .B(_06329_), .Y(_06441_));
AND_g _27241_ (.A(_06440_), .B(_06441_), .Y(_06442_));
NAND_g _27242_ (.A(_13883_), .B(_06442_), .Y(_06443_));
AND_g _27243_ (.A(_14488_), .B(_06443_), .Y(_06444_));
AND_g _27244_ (.A(_06437_), .B(_06444_), .Y(_06445_));
AND_g _27245_ (.A(_06339_), .B(_06445_), .Y(_06446_));
NOR_g _27246_ (.A(_06336_), .B(_06446_), .Y(_01047_));
NOR_g _27247_ (.A(pcpi_rs1[30]), .B(_14488_), .Y(_06447_));
NAND_g _27248_ (.A(reg_pc[30]), .B(_14617_), .Y(_06448_));
NAND_g _27249_ (.A(cpuregs[7][30]), .B(_00008_[2]), .Y(_06449_));
NAND_g _27250_ (.A(cpuregs[3][30]), .B(_09032_), .Y(_06450_));
AND_g _27251_ (.A(_06449_), .B(_06450_), .Y(_06451_));
NAND_g _27252_ (.A(cpuregs[6][30]), .B(_00008_[2]), .Y(_06452_));
NAND_g _27253_ (.A(cpuregs[2][30]), .B(_09032_), .Y(_06453_));
AND_g _27254_ (.A(_06452_), .B(_06453_), .Y(_06454_));
NAND_g _27255_ (.A(_09030_), .B(_06454_), .Y(_06455_));
NAND_g _27256_ (.A(_00008_[0]), .B(_06451_), .Y(_06456_));
AND_g _27257_ (.A(_06455_), .B(_06456_), .Y(_06457_));
NAND_g _27258_ (.A(_00008_[1]), .B(_06457_), .Y(_06458_));
NAND_g _27259_ (.A(cpuregs[4][30]), .B(_00008_[2]), .Y(_06459_));
NAND_g _27260_ (.A(cpuregs[0][30]), .B(_09032_), .Y(_06460_));
AND_g _27261_ (.A(_06459_), .B(_06460_), .Y(_06461_));
NAND_g _27262_ (.A(_09030_), .B(_06461_), .Y(_06462_));
NAND_g _27263_ (.A(cpuregs[5][30]), .B(_00008_[2]), .Y(_06463_));
NAND_g _27264_ (.A(cpuregs[1][30]), .B(_09032_), .Y(_06464_));
AND_g _27265_ (.A(_00008_[0]), .B(_06464_), .Y(_06465_));
NAND_g _27266_ (.A(_06463_), .B(_06465_), .Y(_06466_));
AND_g _27267_ (.A(_06462_), .B(_06466_), .Y(_06467_));
NAND_g _27268_ (.A(_09031_), .B(_06467_), .Y(_06468_));
NAND_g _27269_ (.A(_06458_), .B(_06468_), .Y(_06469_));
NAND_g _27270_ (.A(_09033_), .B(_06469_), .Y(_06470_));
NAND_g _27271_ (.A(cpuregs[11][30]), .B(_09032_), .Y(_06471_));
NAND_g _27272_ (.A(cpuregs[15][30]), .B(_00008_[2]), .Y(_06472_));
NAND_g _27273_ (.A(_06471_), .B(_06472_), .Y(_06473_));
NAND_g _27274_ (.A(_00008_[0]), .B(_06473_), .Y(_06474_));
NAND_g _27275_ (.A(cpuregs[14][30]), .B(_00008_[2]), .Y(_06475_));
NAND_g _27276_ (.A(cpuregs[10][30]), .B(_09032_), .Y(_06476_));
NAND_g _27277_ (.A(_06475_), .B(_06476_), .Y(_06477_));
NAND_g _27278_ (.A(_09030_), .B(_06477_), .Y(_06478_));
NAND_g _27279_ (.A(_06474_), .B(_06478_), .Y(_06479_));
AND_g _27280_ (.A(_00008_[1]), .B(_06479_), .Y(_06480_));
NAND_g _27281_ (.A(_08884_), .B(_00008_[2]), .Y(_06481_));
NOR_g _27282_ (.A(cpuregs[8][30]), .B(_00008_[2]), .Y(_06482_));
NOR_g _27283_ (.A(_00008_[0]), .B(_06482_), .Y(_06483_));
AND_g _27284_ (.A(_06481_), .B(_06483_), .Y(_06484_));
NOR_g _27285_ (.A(cpuregs[9][30]), .B(_00008_[2]), .Y(_06485_));
NAND_g _27286_ (.A(_08935_), .B(_00008_[2]), .Y(_06486_));
NAND_g _27287_ (.A(_00008_[0]), .B(_06486_), .Y(_06487_));
NOR_g _27288_ (.A(_06485_), .B(_06487_), .Y(_06488_));
NOR_g _27289_ (.A(_06484_), .B(_06488_), .Y(_06489_));
NOR_g _27290_ (.A(_00008_[1]), .B(_06489_), .Y(_06490_));
NOR_g _27291_ (.A(_06480_), .B(_06490_), .Y(_06491_));
NOR_g _27292_ (.A(_09033_), .B(_06491_), .Y(_06492_));
NOR_g _27293_ (.A(_00008_[4]), .B(_06492_), .Y(_06493_));
NAND_g _27294_ (.A(_06470_), .B(_06493_), .Y(_06494_));
NAND_g _27295_ (.A(_08903_), .B(_00008_[2]), .Y(_06495_));
NOR_g _27296_ (.A(cpuregs[19][30]), .B(_00008_[2]), .Y(_06496_));
NOR_g _27297_ (.A(cpuregs[18][30]), .B(_00008_[2]), .Y(_06497_));
NOR_g _27298_ (.A(cpuregs[22][30]), .B(_09032_), .Y(_06498_));
NOR_g _27299_ (.A(_06497_), .B(_06498_), .Y(_06499_));
NOR_g _27300_ (.A(_09030_), .B(_06496_), .Y(_06500_));
NAND_g _27301_ (.A(_06495_), .B(_06500_), .Y(_06501_));
NAND_g _27302_ (.A(_09030_), .B(_06499_), .Y(_06502_));
AND_g _27303_ (.A(_06501_), .B(_06502_), .Y(_06503_));
NAND_g _27304_ (.A(_00008_[1]), .B(_06503_), .Y(_06504_));
NOR_g _27305_ (.A(cpuregs[17][30]), .B(_00008_[2]), .Y(_06505_));
NAND_g _27306_ (.A(_09002_), .B(_00008_[2]), .Y(_06506_));
NOR_g _27307_ (.A(cpuregs[16][30]), .B(_00008_[2]), .Y(_06507_));
NOR_g _27308_ (.A(cpuregs[20][30]), .B(_09032_), .Y(_06508_));
NOR_g _27309_ (.A(_06507_), .B(_06508_), .Y(_06509_));
NOR_g _27310_ (.A(_09030_), .B(_06505_), .Y(_06510_));
NAND_g _27311_ (.A(_06506_), .B(_06510_), .Y(_06511_));
NAND_g _27312_ (.A(_09030_), .B(_06509_), .Y(_06512_));
AND_g _27313_ (.A(_06511_), .B(_06512_), .Y(_06513_));
NAND_g _27314_ (.A(_09031_), .B(_06513_), .Y(_06514_));
NAND_g _27315_ (.A(_06504_), .B(_06514_), .Y(_06515_));
NAND_g _27316_ (.A(_09033_), .B(_06515_), .Y(_06516_));
NAND_g _27317_ (.A(cpuregs[25][30]), .B(_09031_), .Y(_06517_));
NAND_g _27318_ (.A(cpuregs[27][30]), .B(_00008_[1]), .Y(_06518_));
AND_g _27319_ (.A(_09032_), .B(_06518_), .Y(_06519_));
NAND_g _27320_ (.A(_06517_), .B(_06519_), .Y(_06520_));
NAND_g _27321_ (.A(cpuregs[29][30]), .B(_09031_), .Y(_06521_));
NAND_g _27322_ (.A(cpuregs[31][30]), .B(_00008_[1]), .Y(_06522_));
AND_g _27323_ (.A(_00008_[2]), .B(_06522_), .Y(_06523_));
NAND_g _27324_ (.A(_06521_), .B(_06523_), .Y(_06524_));
NAND_g _27325_ (.A(_06520_), .B(_06524_), .Y(_06525_));
NAND_g _27326_ (.A(_00008_[0]), .B(_06525_), .Y(_06526_));
NAND_g _27327_ (.A(cpuregs[24][30]), .B(_09031_), .Y(_06527_));
NAND_g _27328_ (.A(cpuregs[26][30]), .B(_00008_[1]), .Y(_06528_));
AND_g _27329_ (.A(_09032_), .B(_06528_), .Y(_06529_));
NAND_g _27330_ (.A(_06527_), .B(_06529_), .Y(_06530_));
NAND_g _27331_ (.A(cpuregs[28][30]), .B(_09031_), .Y(_06531_));
NAND_g _27332_ (.A(cpuregs[30][30]), .B(_00008_[1]), .Y(_06532_));
AND_g _27333_ (.A(_00008_[2]), .B(_06532_), .Y(_06533_));
NAND_g _27334_ (.A(_06531_), .B(_06533_), .Y(_06534_));
NAND_g _27335_ (.A(_06530_), .B(_06534_), .Y(_06535_));
NAND_g _27336_ (.A(_09030_), .B(_06535_), .Y(_06536_));
NAND_g _27337_ (.A(_06526_), .B(_06536_), .Y(_06537_));
NAND_g _27338_ (.A(_00008_[3]), .B(_06537_), .Y(_06538_));
NAND_g _27339_ (.A(_06516_), .B(_06538_), .Y(_06539_));
NAND_g _27340_ (.A(_00008_[4]), .B(_06539_), .Y(_06540_));
AND_g _27341_ (.A(_14624_), .B(_06494_), .Y(_06541_));
NAND_g _27342_ (.A(_06540_), .B(_06541_), .Y(_06542_));
NAND_g _27343_ (.A(_06448_), .B(_06542_), .Y(_06543_));
NAND_g _27344_ (.A(_10595_), .B(_06543_), .Y(_06544_));
NAND_g _27345_ (.A(_06215_), .B(_06329_), .Y(_06545_));
NAND_g _27346_ (.A(pcpi_rs1[29]), .B(_14481_), .Y(_06546_));
AND_g _27347_ (.A(_13879_), .B(_06546_), .Y(_06547_));
NAND_g _27348_ (.A(_06217_), .B(_06547_), .Y(_06548_));
AND_g _27349_ (.A(_06545_), .B(_06548_), .Y(_06549_));
NAND_g _27350_ (.A(_13883_), .B(_06549_), .Y(_06550_));
AND_g _27351_ (.A(_14488_), .B(_06550_), .Y(_06551_));
AND_g _27352_ (.A(_06544_), .B(_06551_), .Y(_06552_));
XOR_g _27353_ (.A(_14492_), .B(_14610_), .Y(_06553_));
NAND_g _27354_ (.A(_14614_), .B(_06553_), .Y(_06554_));
AND_g _27355_ (.A(_06552_), .B(_06554_), .Y(_06555_));
NOR_g _27356_ (.A(_06447_), .B(_06555_), .Y(_01048_));
AND_g _27357_ (.A(_09085_), .B(_02494_), .Y(_06556_));
NAND_g _27358_ (.A(_09085_), .B(_02494_), .Y(_06557_));
NAND_g _27359_ (.A(_09098_), .B(_06556_), .Y(_06558_));
NAND_g _27360_ (.A(cpuregs[7][0]), .B(_06557_), .Y(_06559_));
NAND_g _27361_ (.A(_06558_), .B(_06559_), .Y(_01049_));
NAND_g _27362_ (.A(_09109_), .B(_06556_), .Y(_06560_));
NAND_g _27363_ (.A(cpuregs[7][1]), .B(_06557_), .Y(_06561_));
NAND_g _27364_ (.A(_06560_), .B(_06561_), .Y(_01050_));
NAND_g _27365_ (.A(_09118_), .B(_06556_), .Y(_06562_));
NAND_g _27366_ (.A(cpuregs[7][2]), .B(_06557_), .Y(_06563_));
NAND_g _27367_ (.A(_06562_), .B(_06563_), .Y(_01051_));
NAND_g _27368_ (.A(_09131_), .B(_06556_), .Y(_06564_));
NAND_g _27369_ (.A(cpuregs[7][3]), .B(_06557_), .Y(_06565_));
NAND_g _27370_ (.A(_06564_), .B(_06565_), .Y(_01052_));
NAND_g _27371_ (.A(_09144_), .B(_06556_), .Y(_06566_));
NAND_g _27372_ (.A(cpuregs[7][4]), .B(_06557_), .Y(_06567_));
NAND_g _27373_ (.A(_06566_), .B(_06567_), .Y(_01053_));
NAND_g _27374_ (.A(_09157_), .B(_06556_), .Y(_06568_));
NAND_g _27375_ (.A(cpuregs[7][5]), .B(_06557_), .Y(_06569_));
NAND_g _27376_ (.A(_06568_), .B(_06569_), .Y(_01054_));
NAND_g _27377_ (.A(_09170_), .B(_06556_), .Y(_06570_));
NAND_g _27378_ (.A(cpuregs[7][6]), .B(_06557_), .Y(_06571_));
NAND_g _27379_ (.A(_06570_), .B(_06571_), .Y(_01055_));
NAND_g _27380_ (.A(_09183_), .B(_06556_), .Y(_06572_));
NAND_g _27381_ (.A(cpuregs[7][7]), .B(_06557_), .Y(_06573_));
NAND_g _27382_ (.A(_06572_), .B(_06573_), .Y(_01056_));
NAND_g _27383_ (.A(_09196_), .B(_06556_), .Y(_06574_));
NAND_g _27384_ (.A(cpuregs[7][8]), .B(_06557_), .Y(_06575_));
NAND_g _27385_ (.A(_06574_), .B(_06575_), .Y(_01057_));
NAND_g _27386_ (.A(_09209_), .B(_06556_), .Y(_06576_));
NAND_g _27387_ (.A(cpuregs[7][9]), .B(_06557_), .Y(_06577_));
NAND_g _27388_ (.A(_06576_), .B(_06577_), .Y(_01058_));
NAND_g _27389_ (.A(_09222_), .B(_06556_), .Y(_06578_));
NAND_g _27390_ (.A(cpuregs[7][10]), .B(_06557_), .Y(_06579_));
NAND_g _27391_ (.A(_06578_), .B(_06579_), .Y(_01059_));
NAND_g _27392_ (.A(_09235_), .B(_06556_), .Y(_06580_));
NAND_g _27393_ (.A(cpuregs[7][11]), .B(_06557_), .Y(_06581_));
NAND_g _27394_ (.A(_06580_), .B(_06581_), .Y(_01060_));
NAND_g _27395_ (.A(_09248_), .B(_06556_), .Y(_06582_));
NAND_g _27396_ (.A(cpuregs[7][12]), .B(_06557_), .Y(_06583_));
NAND_g _27397_ (.A(_06582_), .B(_06583_), .Y(_01061_));
NAND_g _27398_ (.A(_09261_), .B(_06556_), .Y(_06584_));
NAND_g _27399_ (.A(cpuregs[7][13]), .B(_06557_), .Y(_06585_));
NAND_g _27400_ (.A(_06584_), .B(_06585_), .Y(_01062_));
NAND_g _27401_ (.A(_09274_), .B(_06556_), .Y(_06586_));
NAND_g _27402_ (.A(cpuregs[7][14]), .B(_06557_), .Y(_06587_));
NAND_g _27403_ (.A(_06586_), .B(_06587_), .Y(_01063_));
NAND_g _27404_ (.A(_09287_), .B(_06556_), .Y(_06588_));
NAND_g _27405_ (.A(cpuregs[7][15]), .B(_06557_), .Y(_06589_));
NAND_g _27406_ (.A(_06588_), .B(_06589_), .Y(_01064_));
NAND_g _27407_ (.A(_09300_), .B(_06556_), .Y(_06590_));
NAND_g _27408_ (.A(cpuregs[7][16]), .B(_06557_), .Y(_06591_));
NAND_g _27409_ (.A(_06590_), .B(_06591_), .Y(_01065_));
NOR_g _27410_ (.A(cpuregs[7][17]), .B(_06556_), .Y(_06592_));
NOR_g _27411_ (.A(_09313_), .B(_06557_), .Y(_06593_));
NOR_g _27412_ (.A(_06592_), .B(_06593_), .Y(_01066_));
AND_g _27413_ (.A(_08972_), .B(_06557_), .Y(_06594_));
NOR_g _27414_ (.A(_09325_), .B(_06557_), .Y(_06595_));
NOR_g _27415_ (.A(_06594_), .B(_06595_), .Y(_01067_));
NAND_g _27416_ (.A(_09338_), .B(_06556_), .Y(_06596_));
NAND_g _27417_ (.A(cpuregs[7][19]), .B(_06557_), .Y(_06597_));
NAND_g _27418_ (.A(_06596_), .B(_06597_), .Y(_01068_));
NAND_g _27419_ (.A(_09351_), .B(_06556_), .Y(_06598_));
NAND_g _27420_ (.A(cpuregs[7][20]), .B(_06557_), .Y(_06599_));
NAND_g _27421_ (.A(_06598_), .B(_06599_), .Y(_01069_));
NAND_g _27422_ (.A(_09364_), .B(_06556_), .Y(_06600_));
NAND_g _27423_ (.A(cpuregs[7][21]), .B(_06557_), .Y(_06601_));
NAND_g _27424_ (.A(_06600_), .B(_06601_), .Y(_01070_));
NAND_g _27425_ (.A(_09377_), .B(_06556_), .Y(_06602_));
NAND_g _27426_ (.A(cpuregs[7][22]), .B(_06557_), .Y(_06603_));
NAND_g _27427_ (.A(_06602_), .B(_06603_), .Y(_01071_));
NAND_g _27428_ (.A(_09390_), .B(_06556_), .Y(_06604_));
NAND_g _27429_ (.A(cpuregs[7][23]), .B(_06557_), .Y(_06605_));
NAND_g _27430_ (.A(_06604_), .B(_06605_), .Y(_01072_));
NAND_g _27431_ (.A(_09403_), .B(_06556_), .Y(_06606_));
NAND_g _27432_ (.A(cpuregs[7][24]), .B(_06557_), .Y(_06607_));
NAND_g _27433_ (.A(_06606_), .B(_06607_), .Y(_01073_));
NAND_g _27434_ (.A(_09416_), .B(_06556_), .Y(_06608_));
NAND_g _27435_ (.A(cpuregs[7][25]), .B(_06557_), .Y(_06609_));
NAND_g _27436_ (.A(_06608_), .B(_06609_), .Y(_01074_));
NAND_g _27437_ (.A(_09429_), .B(_06556_), .Y(_06610_));
NAND_g _27438_ (.A(cpuregs[7][26]), .B(_06557_), .Y(_06611_));
NAND_g _27439_ (.A(_06610_), .B(_06611_), .Y(_01075_));
NAND_g _27440_ (.A(_09442_), .B(_06556_), .Y(_06612_));
NAND_g _27441_ (.A(cpuregs[7][27]), .B(_06557_), .Y(_06613_));
NAND_g _27442_ (.A(_06612_), .B(_06613_), .Y(_01076_));
NAND_g _27443_ (.A(_09455_), .B(_06556_), .Y(_06614_));
NAND_g _27444_ (.A(cpuregs[7][28]), .B(_06557_), .Y(_06615_));
NAND_g _27445_ (.A(_06614_), .B(_06615_), .Y(_01077_));
NAND_g _27446_ (.A(_09468_), .B(_06556_), .Y(_06616_));
NAND_g _27447_ (.A(cpuregs[7][29]), .B(_06557_), .Y(_06617_));
NAND_g _27448_ (.A(_06616_), .B(_06617_), .Y(_01078_));
NAND_g _27449_ (.A(_09481_), .B(_06556_), .Y(_06618_));
NAND_g _27450_ (.A(cpuregs[7][30]), .B(_06557_), .Y(_06619_));
NAND_g _27451_ (.A(_06618_), .B(_06619_), .Y(_01079_));
NAND_g _27452_ (.A(_09493_), .B(_06556_), .Y(_06620_));
NAND_g _27453_ (.A(cpuregs[7][31]), .B(_06557_), .Y(_06621_));
NAND_g _27454_ (.A(_06620_), .B(_06621_), .Y(_01080_));
AND_g _27455_ (.A(_09077_), .B(_09080_), .Y(_06622_));
NAND_g _27456_ (.A(_09077_), .B(_09080_), .Y(_06623_));
NAND_g _27457_ (.A(cpuregs[8][0]), .B(_06623_), .Y(_06624_));
NAND_g _27458_ (.A(_09097_), .B(_06622_), .Y(_06625_));
NAND_g _27459_ (.A(_06624_), .B(_06625_), .Y(_01081_));
NAND_g _27460_ (.A(cpuregs[8][1]), .B(_06623_), .Y(_06626_));
NAND_g _27461_ (.A(_09108_), .B(_06622_), .Y(_06627_));
NAND_g _27462_ (.A(_06626_), .B(_06627_), .Y(_01082_));
NAND_g _27463_ (.A(cpuregs[8][2]), .B(_06623_), .Y(_06628_));
NAND_g _27464_ (.A(_09117_), .B(_06622_), .Y(_06629_));
NAND_g _27465_ (.A(_06628_), .B(_06629_), .Y(_01083_));
NAND_g _27466_ (.A(cpuregs[8][3]), .B(_06623_), .Y(_06630_));
NAND_g _27467_ (.A(_09130_), .B(_06622_), .Y(_06631_));
NAND_g _27468_ (.A(_06630_), .B(_06631_), .Y(_01084_));
NAND_g _27469_ (.A(cpuregs[8][4]), .B(_06623_), .Y(_06632_));
NAND_g _27470_ (.A(_09143_), .B(_06622_), .Y(_06633_));
NAND_g _27471_ (.A(_06632_), .B(_06633_), .Y(_01085_));
NAND_g _27472_ (.A(cpuregs[8][5]), .B(_06623_), .Y(_06634_));
NAND_g _27473_ (.A(_09156_), .B(_06622_), .Y(_06635_));
NAND_g _27474_ (.A(_06634_), .B(_06635_), .Y(_01086_));
NAND_g _27475_ (.A(cpuregs[8][6]), .B(_06623_), .Y(_06636_));
NAND_g _27476_ (.A(_09169_), .B(_06622_), .Y(_06637_));
NAND_g _27477_ (.A(_06636_), .B(_06637_), .Y(_01087_));
NAND_g _27478_ (.A(cpuregs[8][7]), .B(_06623_), .Y(_06638_));
NAND_g _27479_ (.A(_09182_), .B(_06622_), .Y(_06639_));
NAND_g _27480_ (.A(_06638_), .B(_06639_), .Y(_01088_));
NAND_g _27481_ (.A(cpuregs[8][8]), .B(_06623_), .Y(_06640_));
NAND_g _27482_ (.A(_09195_), .B(_06622_), .Y(_06641_));
NAND_g _27483_ (.A(_06640_), .B(_06641_), .Y(_01089_));
NAND_g _27484_ (.A(cpuregs[8][9]), .B(_06623_), .Y(_06642_));
NAND_g _27485_ (.A(_09208_), .B(_06622_), .Y(_06643_));
NAND_g _27486_ (.A(_06642_), .B(_06643_), .Y(_01090_));
NAND_g _27487_ (.A(cpuregs[8][10]), .B(_06623_), .Y(_06644_));
NAND_g _27488_ (.A(_09221_), .B(_06622_), .Y(_06645_));
NAND_g _27489_ (.A(_06644_), .B(_06645_), .Y(_01091_));
NAND_g _27490_ (.A(cpuregs[8][11]), .B(_06623_), .Y(_06646_));
NAND_g _27491_ (.A(_09234_), .B(_06622_), .Y(_06647_));
NAND_g _27492_ (.A(_06646_), .B(_06647_), .Y(_01092_));
NAND_g _27493_ (.A(cpuregs[8][12]), .B(_06623_), .Y(_06648_));
NAND_g _27494_ (.A(_09247_), .B(_06622_), .Y(_06649_));
NAND_g _27495_ (.A(_06648_), .B(_06649_), .Y(_01093_));
NAND_g _27496_ (.A(cpuregs[8][13]), .B(_06623_), .Y(_06650_));
NAND_g _27497_ (.A(_09260_), .B(_06622_), .Y(_06651_));
NAND_g _27498_ (.A(_06650_), .B(_06651_), .Y(_01094_));
NAND_g _27499_ (.A(cpuregs[8][14]), .B(_06623_), .Y(_06652_));
NAND_g _27500_ (.A(_09273_), .B(_06622_), .Y(_06653_));
NAND_g _27501_ (.A(_06652_), .B(_06653_), .Y(_01095_));
NAND_g _27502_ (.A(cpuregs[8][15]), .B(_06623_), .Y(_06654_));
NAND_g _27503_ (.A(_09286_), .B(_06622_), .Y(_06655_));
NAND_g _27504_ (.A(_06654_), .B(_06655_), .Y(_01096_));
NAND_g _27505_ (.A(_09299_), .B(_06622_), .Y(_06656_));
NAND_g _27506_ (.A(cpuregs[8][16]), .B(_06623_), .Y(_06657_));
NAND_g _27507_ (.A(_06656_), .B(_06657_), .Y(_01097_));
NAND_g _27508_ (.A(_09312_), .B(_06622_), .Y(_06658_));
NAND_g _27509_ (.A(cpuregs[8][17]), .B(_06623_), .Y(_06659_));
NAND_g _27510_ (.A(_06658_), .B(_06659_), .Y(_01098_));
NAND_g _27511_ (.A(_09324_), .B(_06622_), .Y(_06660_));
NAND_g _27512_ (.A(cpuregs[8][18]), .B(_06623_), .Y(_06661_));
NAND_g _27513_ (.A(_06660_), .B(_06661_), .Y(_01099_));
NAND_g _27514_ (.A(_09337_), .B(_06622_), .Y(_06662_));
NAND_g _27515_ (.A(cpuregs[8][19]), .B(_06623_), .Y(_06663_));
NAND_g _27516_ (.A(_06662_), .B(_06663_), .Y(_01100_));
NAND_g _27517_ (.A(_09350_), .B(_06622_), .Y(_06664_));
NAND_g _27518_ (.A(cpuregs[8][20]), .B(_06623_), .Y(_06665_));
NAND_g _27519_ (.A(_06664_), .B(_06665_), .Y(_01101_));
NAND_g _27520_ (.A(_09363_), .B(_06622_), .Y(_06666_));
NAND_g _27521_ (.A(cpuregs[8][21]), .B(_06623_), .Y(_06667_));
NAND_g _27522_ (.A(_06666_), .B(_06667_), .Y(_01102_));
NAND_g _27523_ (.A(_09376_), .B(_06622_), .Y(_06668_));
NAND_g _27524_ (.A(cpuregs[8][22]), .B(_06623_), .Y(_06669_));
NAND_g _27525_ (.A(_06668_), .B(_06669_), .Y(_01103_));
NAND_g _27526_ (.A(_09389_), .B(_06622_), .Y(_06670_));
NAND_g _27527_ (.A(cpuregs[8][23]), .B(_06623_), .Y(_06671_));
NAND_g _27528_ (.A(_06670_), .B(_06671_), .Y(_01104_));
NAND_g _27529_ (.A(_09402_), .B(_06622_), .Y(_06672_));
NAND_g _27530_ (.A(cpuregs[8][24]), .B(_06623_), .Y(_06673_));
NAND_g _27531_ (.A(_06672_), .B(_06673_), .Y(_01105_));
NAND_g _27532_ (.A(_09415_), .B(_06622_), .Y(_06674_));
NAND_g _27533_ (.A(cpuregs[8][25]), .B(_06623_), .Y(_06675_));
NAND_g _27534_ (.A(_06674_), .B(_06675_), .Y(_01106_));
NAND_g _27535_ (.A(_09428_), .B(_06622_), .Y(_06676_));
NAND_g _27536_ (.A(cpuregs[8][26]), .B(_06623_), .Y(_06677_));
NAND_g _27537_ (.A(_06676_), .B(_06677_), .Y(_01107_));
NAND_g _27538_ (.A(_09441_), .B(_06622_), .Y(_06678_));
NAND_g _27539_ (.A(cpuregs[8][27]), .B(_06623_), .Y(_06679_));
NAND_g _27540_ (.A(_06678_), .B(_06679_), .Y(_01108_));
NAND_g _27541_ (.A(_09454_), .B(_06622_), .Y(_06680_));
NAND_g _27542_ (.A(cpuregs[8][28]), .B(_06623_), .Y(_06681_));
NAND_g _27543_ (.A(_06680_), .B(_06681_), .Y(_01109_));
NAND_g _27544_ (.A(_09467_), .B(_06622_), .Y(_06682_));
NAND_g _27545_ (.A(cpuregs[8][29]), .B(_06623_), .Y(_06683_));
NAND_g _27546_ (.A(_06682_), .B(_06683_), .Y(_01110_));
NAND_g _27547_ (.A(_09480_), .B(_06622_), .Y(_06684_));
NAND_g _27548_ (.A(cpuregs[8][30]), .B(_06623_), .Y(_06685_));
NAND_g _27549_ (.A(_06684_), .B(_06685_), .Y(_01111_));
NAND_g _27550_ (.A(_09492_), .B(_06622_), .Y(_06686_));
NAND_g _27551_ (.A(cpuregs[8][31]), .B(_06623_), .Y(_06687_));
NAND_g _27552_ (.A(_06686_), .B(_06687_), .Y(_01112_));
NAND_g _27553_ (.A(_14393_), .B(_00442_), .Y(_06688_));
NAND_g _27554_ (.A(decoded_imm_j[8]), .B(_14394_), .Y(_06689_));
NAND_g _27555_ (.A(_06688_), .B(_06689_), .Y(_01145_));
NAND_g _27556_ (.A(_14393_), .B(_00443_), .Y(_06690_));
NAND_g _27557_ (.A(decoded_imm_j[9]), .B(_14394_), .Y(_06691_));
NAND_g _27558_ (.A(_06690_), .B(_06691_), .Y(_01146_));
NOR_g _27559_ (.A(latched_rd[2]), .B(_09498_), .Y(_06692_));
AND_g _27560_ (.A(_09496_), .B(_06692_), .Y(_06693_));
NAND_g _27561_ (.A(_09496_), .B(_06692_), .Y(_06694_));
NAND_g _27562_ (.A(cpuregs[26][0]), .B(_06694_), .Y(_06695_));
NAND_g _27563_ (.A(_09098_), .B(_06693_), .Y(_06696_));
NAND_g _27564_ (.A(_06695_), .B(_06696_), .Y(_01147_));
NAND_g _27565_ (.A(cpuregs[26][1]), .B(_06694_), .Y(_06697_));
NAND_g _27566_ (.A(_09109_), .B(_06693_), .Y(_06698_));
NAND_g _27567_ (.A(_06697_), .B(_06698_), .Y(_01148_));
NAND_g _27568_ (.A(cpuregs[26][2]), .B(_06694_), .Y(_06699_));
NAND_g _27569_ (.A(_09118_), .B(_06693_), .Y(_06700_));
NAND_g _27570_ (.A(_06699_), .B(_06700_), .Y(_01149_));
NAND_g _27571_ (.A(cpuregs[26][3]), .B(_06694_), .Y(_06701_));
NAND_g _27572_ (.A(_09131_), .B(_06693_), .Y(_06702_));
NAND_g _27573_ (.A(_06701_), .B(_06702_), .Y(_01150_));
NAND_g _27574_ (.A(cpuregs[26][4]), .B(_06694_), .Y(_06703_));
NAND_g _27575_ (.A(_09144_), .B(_06693_), .Y(_06704_));
NAND_g _27576_ (.A(_06703_), .B(_06704_), .Y(_01151_));
NAND_g _27577_ (.A(cpuregs[26][5]), .B(_06694_), .Y(_06705_));
NAND_g _27578_ (.A(_09157_), .B(_06693_), .Y(_06706_));
NAND_g _27579_ (.A(_06705_), .B(_06706_), .Y(_01152_));
NAND_g _27580_ (.A(cpuregs[26][6]), .B(_06694_), .Y(_06707_));
NAND_g _27581_ (.A(_09170_), .B(_06693_), .Y(_06708_));
NAND_g _27582_ (.A(_06707_), .B(_06708_), .Y(_01153_));
NAND_g _27583_ (.A(cpuregs[26][7]), .B(_06694_), .Y(_06709_));
NAND_g _27584_ (.A(_09183_), .B(_06693_), .Y(_06710_));
NAND_g _27585_ (.A(_06709_), .B(_06710_), .Y(_01154_));
NAND_g _27586_ (.A(cpuregs[26][8]), .B(_06694_), .Y(_06711_));
NAND_g _27587_ (.A(_09196_), .B(_06693_), .Y(_06712_));
NAND_g _27588_ (.A(_06711_), .B(_06712_), .Y(_01155_));
NAND_g _27589_ (.A(cpuregs[26][9]), .B(_06694_), .Y(_06713_));
NAND_g _27590_ (.A(_09209_), .B(_06693_), .Y(_06714_));
NAND_g _27591_ (.A(_06713_), .B(_06714_), .Y(_01156_));
NAND_g _27592_ (.A(cpuregs[26][10]), .B(_06694_), .Y(_06715_));
NAND_g _27593_ (.A(_09222_), .B(_06693_), .Y(_06716_));
NAND_g _27594_ (.A(_06715_), .B(_06716_), .Y(_01157_));
NAND_g _27595_ (.A(cpuregs[26][11]), .B(_06694_), .Y(_06717_));
NAND_g _27596_ (.A(_09235_), .B(_06693_), .Y(_06718_));
NAND_g _27597_ (.A(_06717_), .B(_06718_), .Y(_01158_));
NAND_g _27598_ (.A(cpuregs[26][12]), .B(_06694_), .Y(_06719_));
NAND_g _27599_ (.A(_09248_), .B(_06693_), .Y(_06720_));
NAND_g _27600_ (.A(_06719_), .B(_06720_), .Y(_01159_));
NAND_g _27601_ (.A(cpuregs[26][13]), .B(_06694_), .Y(_06721_));
NAND_g _27602_ (.A(_09261_), .B(_06693_), .Y(_06722_));
NAND_g _27603_ (.A(_06721_), .B(_06722_), .Y(_01160_));
NAND_g _27604_ (.A(cpuregs[26][14]), .B(_06694_), .Y(_06723_));
NAND_g _27605_ (.A(_09274_), .B(_06693_), .Y(_06724_));
NAND_g _27606_ (.A(_06723_), .B(_06724_), .Y(_01161_));
NAND_g _27607_ (.A(cpuregs[26][15]), .B(_06694_), .Y(_06725_));
NAND_g _27608_ (.A(_09287_), .B(_06693_), .Y(_06726_));
NAND_g _27609_ (.A(_06725_), .B(_06726_), .Y(_01162_));
NAND_g _27610_ (.A(cpuregs[26][16]), .B(_06694_), .Y(_06727_));
NAND_g _27611_ (.A(_09300_), .B(_06693_), .Y(_06728_));
NAND_g _27612_ (.A(_06727_), .B(_06728_), .Y(_01163_));
NOR_g _27613_ (.A(cpuregs[26][17]), .B(_06693_), .Y(_06729_));
NOR_g _27614_ (.A(_09313_), .B(_06694_), .Y(_06730_));
NOR_g _27615_ (.A(_06729_), .B(_06730_), .Y(_01164_));
NAND_g _27616_ (.A(cpuregs[26][18]), .B(_06694_), .Y(_06731_));
NAND_g _27617_ (.A(_09325_), .B(_06693_), .Y(_06732_));
NAND_g _27618_ (.A(_06731_), .B(_06732_), .Y(_01165_));
NAND_g _27619_ (.A(cpuregs[26][19]), .B(_06694_), .Y(_06733_));
NAND_g _27620_ (.A(_09338_), .B(_06693_), .Y(_06734_));
NAND_g _27621_ (.A(_06733_), .B(_06734_), .Y(_01166_));
NAND_g _27622_ (.A(cpuregs[26][20]), .B(_06694_), .Y(_06735_));
NAND_g _27623_ (.A(_09351_), .B(_06693_), .Y(_06736_));
NAND_g _27624_ (.A(_06735_), .B(_06736_), .Y(_01167_));
NAND_g _27625_ (.A(cpuregs[26][21]), .B(_06694_), .Y(_06737_));
NAND_g _27626_ (.A(_09364_), .B(_06693_), .Y(_06738_));
NAND_g _27627_ (.A(_06737_), .B(_06738_), .Y(_01168_));
NAND_g _27628_ (.A(cpuregs[26][22]), .B(_06694_), .Y(_06739_));
NAND_g _27629_ (.A(_09377_), .B(_06693_), .Y(_06740_));
NAND_g _27630_ (.A(_06739_), .B(_06740_), .Y(_01169_));
NAND_g _27631_ (.A(cpuregs[26][23]), .B(_06694_), .Y(_06741_));
NAND_g _27632_ (.A(_09390_), .B(_06693_), .Y(_06742_));
NAND_g _27633_ (.A(_06741_), .B(_06742_), .Y(_01170_));
NAND_g _27634_ (.A(cpuregs[26][24]), .B(_06694_), .Y(_06743_));
NAND_g _27635_ (.A(_09403_), .B(_06693_), .Y(_06744_));
NAND_g _27636_ (.A(_06743_), .B(_06744_), .Y(_01171_));
NAND_g _27637_ (.A(cpuregs[26][25]), .B(_06694_), .Y(_06745_));
NAND_g _27638_ (.A(_09416_), .B(_06693_), .Y(_06746_));
NAND_g _27639_ (.A(_06745_), .B(_06746_), .Y(_01172_));
NAND_g _27640_ (.A(cpuregs[26][26]), .B(_06694_), .Y(_06747_));
NAND_g _27641_ (.A(_09429_), .B(_06693_), .Y(_06748_));
NAND_g _27642_ (.A(_06747_), .B(_06748_), .Y(_01173_));
NAND_g _27643_ (.A(cpuregs[26][27]), .B(_06694_), .Y(_06749_));
NAND_g _27644_ (.A(_09442_), .B(_06693_), .Y(_06750_));
NAND_g _27645_ (.A(_06749_), .B(_06750_), .Y(_01174_));
NAND_g _27646_ (.A(cpuregs[26][28]), .B(_06694_), .Y(_06751_));
NAND_g _27647_ (.A(_09455_), .B(_06693_), .Y(_06752_));
NAND_g _27648_ (.A(_06751_), .B(_06752_), .Y(_01175_));
NAND_g _27649_ (.A(cpuregs[26][29]), .B(_06694_), .Y(_06753_));
NAND_g _27650_ (.A(_09468_), .B(_06693_), .Y(_06754_));
NAND_g _27651_ (.A(_06753_), .B(_06754_), .Y(_01176_));
NAND_g _27652_ (.A(cpuregs[26][30]), .B(_06694_), .Y(_06755_));
NAND_g _27653_ (.A(_09481_), .B(_06693_), .Y(_06756_));
NAND_g _27654_ (.A(_06755_), .B(_06756_), .Y(_01177_));
NAND_g _27655_ (.A(cpuregs[26][31]), .B(_06694_), .Y(_06757_));
NAND_g _27656_ (.A(_09493_), .B(_06693_), .Y(_06758_));
NAND_g _27657_ (.A(_06757_), .B(_06758_), .Y(_01178_));
AND_g _27658_ (.A(_09085_), .B(_09499_), .Y(_06759_));
NAND_g _27659_ (.A(_09085_), .B(_09499_), .Y(_06760_));
NAND_g _27660_ (.A(_09098_), .B(_06759_), .Y(_06761_));
NAND_g _27661_ (.A(cpuregs[31][0]), .B(_06760_), .Y(_06762_));
NAND_g _27662_ (.A(_06761_), .B(_06762_), .Y(_01179_));
NAND_g _27663_ (.A(_09109_), .B(_06759_), .Y(_06763_));
NAND_g _27664_ (.A(cpuregs[31][1]), .B(_06760_), .Y(_06764_));
NAND_g _27665_ (.A(_06763_), .B(_06764_), .Y(_01180_));
NAND_g _27666_ (.A(_09118_), .B(_06759_), .Y(_06765_));
NAND_g _27667_ (.A(cpuregs[31][2]), .B(_06760_), .Y(_06766_));
NAND_g _27668_ (.A(_06765_), .B(_06766_), .Y(_01181_));
NAND_g _27669_ (.A(_09131_), .B(_06759_), .Y(_06767_));
NAND_g _27670_ (.A(cpuregs[31][3]), .B(_06760_), .Y(_06768_));
NAND_g _27671_ (.A(_06767_), .B(_06768_), .Y(_01182_));
NAND_g _27672_ (.A(_09144_), .B(_06759_), .Y(_06769_));
NAND_g _27673_ (.A(cpuregs[31][4]), .B(_06760_), .Y(_06770_));
NAND_g _27674_ (.A(_06769_), .B(_06770_), .Y(_01183_));
NAND_g _27675_ (.A(_09157_), .B(_06759_), .Y(_06771_));
NAND_g _27676_ (.A(cpuregs[31][5]), .B(_06760_), .Y(_06772_));
NAND_g _27677_ (.A(_06771_), .B(_06772_), .Y(_01184_));
NAND_g _27678_ (.A(_09170_), .B(_06759_), .Y(_06773_));
NAND_g _27679_ (.A(cpuregs[31][6]), .B(_06760_), .Y(_06774_));
NAND_g _27680_ (.A(_06773_), .B(_06774_), .Y(_01185_));
NAND_g _27681_ (.A(_09183_), .B(_06759_), .Y(_06775_));
NAND_g _27682_ (.A(cpuregs[31][7]), .B(_06760_), .Y(_06776_));
NAND_g _27683_ (.A(_06775_), .B(_06776_), .Y(_01186_));
NAND_g _27684_ (.A(_09196_), .B(_06759_), .Y(_06777_));
NAND_g _27685_ (.A(cpuregs[31][8]), .B(_06760_), .Y(_06778_));
NAND_g _27686_ (.A(_06777_), .B(_06778_), .Y(_01187_));
NAND_g _27687_ (.A(_09209_), .B(_06759_), .Y(_06779_));
NAND_g _27688_ (.A(cpuregs[31][9]), .B(_06760_), .Y(_06780_));
NAND_g _27689_ (.A(_06779_), .B(_06780_), .Y(_01188_));
NAND_g _27690_ (.A(_09222_), .B(_06759_), .Y(_06781_));
NAND_g _27691_ (.A(cpuregs[31][10]), .B(_06760_), .Y(_06782_));
NAND_g _27692_ (.A(_06781_), .B(_06782_), .Y(_01189_));
NAND_g _27693_ (.A(_09235_), .B(_06759_), .Y(_06783_));
NAND_g _27694_ (.A(cpuregs[31][11]), .B(_06760_), .Y(_06784_));
NAND_g _27695_ (.A(_06783_), .B(_06784_), .Y(_01190_));
NAND_g _27696_ (.A(_09248_), .B(_06759_), .Y(_06785_));
NAND_g _27697_ (.A(cpuregs[31][12]), .B(_06760_), .Y(_06786_));
NAND_g _27698_ (.A(_06785_), .B(_06786_), .Y(_01191_));
NAND_g _27699_ (.A(_09261_), .B(_06759_), .Y(_06787_));
NAND_g _27700_ (.A(cpuregs[31][13]), .B(_06760_), .Y(_06788_));
NAND_g _27701_ (.A(_06787_), .B(_06788_), .Y(_01192_));
NAND_g _27702_ (.A(_09274_), .B(_06759_), .Y(_06789_));
NAND_g _27703_ (.A(cpuregs[31][14]), .B(_06760_), .Y(_06790_));
NAND_g _27704_ (.A(_06789_), .B(_06790_), .Y(_01193_));
NAND_g _27705_ (.A(_09287_), .B(_06759_), .Y(_06791_));
NAND_g _27706_ (.A(cpuregs[31][15]), .B(_06760_), .Y(_06792_));
NAND_g _27707_ (.A(_06791_), .B(_06792_), .Y(_01194_));
NAND_g _27708_ (.A(_09300_), .B(_06759_), .Y(_06793_));
NAND_g _27709_ (.A(cpuregs[31][16]), .B(_06760_), .Y(_06794_));
NAND_g _27710_ (.A(_06793_), .B(_06794_), .Y(_01195_));
NOR_g _27711_ (.A(cpuregs[31][17]), .B(_06759_), .Y(_06795_));
NOR_g _27712_ (.A(_09313_), .B(_06760_), .Y(_06796_));
NOR_g _27713_ (.A(_06795_), .B(_06796_), .Y(_01196_));
NAND_g _27714_ (.A(_09325_), .B(_06759_), .Y(_06797_));
NAND_g _27715_ (.A(cpuregs[31][18]), .B(_06760_), .Y(_06798_));
NAND_g _27716_ (.A(_06797_), .B(_06798_), .Y(_01197_));
NAND_g _27717_ (.A(_09338_), .B(_06759_), .Y(_06799_));
NAND_g _27718_ (.A(cpuregs[31][19]), .B(_06760_), .Y(_06800_));
NAND_g _27719_ (.A(_06799_), .B(_06800_), .Y(_01198_));
NAND_g _27720_ (.A(_09351_), .B(_06759_), .Y(_06801_));
NAND_g _27721_ (.A(cpuregs[31][20]), .B(_06760_), .Y(_06802_));
NAND_g _27722_ (.A(_06801_), .B(_06802_), .Y(_01199_));
NAND_g _27723_ (.A(_09364_), .B(_06759_), .Y(_06803_));
NAND_g _27724_ (.A(cpuregs[31][21]), .B(_06760_), .Y(_06804_));
NAND_g _27725_ (.A(_06803_), .B(_06804_), .Y(_01200_));
NAND_g _27726_ (.A(_09377_), .B(_06759_), .Y(_06805_));
NAND_g _27727_ (.A(cpuregs[31][22]), .B(_06760_), .Y(_06806_));
NAND_g _27728_ (.A(_06805_), .B(_06806_), .Y(_01201_));
NAND_g _27729_ (.A(_09390_), .B(_06759_), .Y(_06807_));
NAND_g _27730_ (.A(cpuregs[31][23]), .B(_06760_), .Y(_06808_));
NAND_g _27731_ (.A(_06807_), .B(_06808_), .Y(_01202_));
NAND_g _27732_ (.A(_09403_), .B(_06759_), .Y(_06809_));
NAND_g _27733_ (.A(cpuregs[31][24]), .B(_06760_), .Y(_06810_));
NAND_g _27734_ (.A(_06809_), .B(_06810_), .Y(_01203_));
NAND_g _27735_ (.A(_09416_), .B(_06759_), .Y(_06811_));
NAND_g _27736_ (.A(cpuregs[31][25]), .B(_06760_), .Y(_06812_));
NAND_g _27737_ (.A(_06811_), .B(_06812_), .Y(_01204_));
NAND_g _27738_ (.A(_09429_), .B(_06759_), .Y(_06813_));
NAND_g _27739_ (.A(cpuregs[31][26]), .B(_06760_), .Y(_06814_));
NAND_g _27740_ (.A(_06813_), .B(_06814_), .Y(_01205_));
NAND_g _27741_ (.A(_09442_), .B(_06759_), .Y(_06815_));
NAND_g _27742_ (.A(cpuregs[31][27]), .B(_06760_), .Y(_06816_));
NAND_g _27743_ (.A(_06815_), .B(_06816_), .Y(_01206_));
NAND_g _27744_ (.A(_09455_), .B(_06759_), .Y(_06817_));
NAND_g _27745_ (.A(cpuregs[31][28]), .B(_06760_), .Y(_06818_));
NAND_g _27746_ (.A(_06817_), .B(_06818_), .Y(_01207_));
NAND_g _27747_ (.A(_09468_), .B(_06759_), .Y(_06819_));
NAND_g _27748_ (.A(cpuregs[31][29]), .B(_06760_), .Y(_06820_));
NAND_g _27749_ (.A(_06819_), .B(_06820_), .Y(_01208_));
NAND_g _27750_ (.A(_09481_), .B(_06759_), .Y(_06821_));
NAND_g _27751_ (.A(cpuregs[31][30]), .B(_06760_), .Y(_06822_));
NAND_g _27752_ (.A(_06821_), .B(_06822_), .Y(_01209_));
NAND_g _27753_ (.A(_09493_), .B(_06759_), .Y(_06823_));
NAND_g _27754_ (.A(cpuregs[31][31]), .B(_06760_), .Y(_06824_));
NAND_g _27755_ (.A(_06823_), .B(_06824_), .Y(_01210_));
AND_g _27756_ (.A(_09085_), .B(_02760_), .Y(_06825_));
NAND_g _27757_ (.A(_09085_), .B(_02760_), .Y(_06826_));
NAND_g _27758_ (.A(_09098_), .B(_06825_), .Y(_06827_));
NAND_g _27759_ (.A(cpuregs[19][0]), .B(_06826_), .Y(_06828_));
NAND_g _27760_ (.A(_06827_), .B(_06828_), .Y(_01211_));
NAND_g _27761_ (.A(_09109_), .B(_06825_), .Y(_06829_));
NAND_g _27762_ (.A(cpuregs[19][1]), .B(_06826_), .Y(_06830_));
NAND_g _27763_ (.A(_06829_), .B(_06830_), .Y(_01212_));
NAND_g _27764_ (.A(_09118_), .B(_06825_), .Y(_06831_));
NAND_g _27765_ (.A(cpuregs[19][2]), .B(_06826_), .Y(_06832_));
NAND_g _27766_ (.A(_06831_), .B(_06832_), .Y(_01213_));
NAND_g _27767_ (.A(_09131_), .B(_06825_), .Y(_06833_));
NAND_g _27768_ (.A(cpuregs[19][3]), .B(_06826_), .Y(_06834_));
NAND_g _27769_ (.A(_06833_), .B(_06834_), .Y(_01214_));
NAND_g _27770_ (.A(_09144_), .B(_06825_), .Y(_06835_));
NAND_g _27771_ (.A(cpuregs[19][4]), .B(_06826_), .Y(_06836_));
NAND_g _27772_ (.A(_06835_), .B(_06836_), .Y(_01215_));
NAND_g _27773_ (.A(_09157_), .B(_06825_), .Y(_06837_));
NAND_g _27774_ (.A(cpuregs[19][5]), .B(_06826_), .Y(_06838_));
NAND_g _27775_ (.A(_06837_), .B(_06838_), .Y(_01216_));
NAND_g _27776_ (.A(_09170_), .B(_06825_), .Y(_06839_));
NAND_g _27777_ (.A(cpuregs[19][6]), .B(_06826_), .Y(_06840_));
NAND_g _27778_ (.A(_06839_), .B(_06840_), .Y(_01217_));
NAND_g _27779_ (.A(_09183_), .B(_06825_), .Y(_06841_));
NAND_g _27780_ (.A(cpuregs[19][7]), .B(_06826_), .Y(_06842_));
NAND_g _27781_ (.A(_06841_), .B(_06842_), .Y(_01218_));
NAND_g _27782_ (.A(_09196_), .B(_06825_), .Y(_06843_));
NAND_g _27783_ (.A(cpuregs[19][8]), .B(_06826_), .Y(_06844_));
NAND_g _27784_ (.A(_06843_), .B(_06844_), .Y(_01219_));
NAND_g _27785_ (.A(_09209_), .B(_06825_), .Y(_06845_));
NAND_g _27786_ (.A(cpuregs[19][9]), .B(_06826_), .Y(_06846_));
NAND_g _27787_ (.A(_06845_), .B(_06846_), .Y(_01220_));
NAND_g _27788_ (.A(_09222_), .B(_06825_), .Y(_06847_));
NAND_g _27789_ (.A(cpuregs[19][10]), .B(_06826_), .Y(_06848_));
NAND_g _27790_ (.A(_06847_), .B(_06848_), .Y(_01221_));
NAND_g _27791_ (.A(_09235_), .B(_06825_), .Y(_06849_));
NAND_g _27792_ (.A(cpuregs[19][11]), .B(_06826_), .Y(_06850_));
NAND_g _27793_ (.A(_06849_), .B(_06850_), .Y(_01222_));
NAND_g _27794_ (.A(_09248_), .B(_06825_), .Y(_06851_));
NAND_g _27795_ (.A(cpuregs[19][12]), .B(_06826_), .Y(_06852_));
NAND_g _27796_ (.A(_06851_), .B(_06852_), .Y(_01223_));
NAND_g _27797_ (.A(_09261_), .B(_06825_), .Y(_06853_));
NAND_g _27798_ (.A(cpuregs[19][13]), .B(_06826_), .Y(_06854_));
NAND_g _27799_ (.A(_06853_), .B(_06854_), .Y(_01224_));
NAND_g _27800_ (.A(_09274_), .B(_06825_), .Y(_06855_));
NAND_g _27801_ (.A(cpuregs[19][14]), .B(_06826_), .Y(_06856_));
NAND_g _27802_ (.A(_06855_), .B(_06856_), .Y(_01225_));
NAND_g _27803_ (.A(_09287_), .B(_06825_), .Y(_06857_));
NAND_g _27804_ (.A(cpuregs[19][15]), .B(_06826_), .Y(_06858_));
NAND_g _27805_ (.A(_06857_), .B(_06858_), .Y(_01226_));
NAND_g _27806_ (.A(_09300_), .B(_06825_), .Y(_06859_));
NAND_g _27807_ (.A(cpuregs[19][16]), .B(_06826_), .Y(_06860_));
NAND_g _27808_ (.A(_06859_), .B(_06860_), .Y(_01227_));
NOR_g _27809_ (.A(cpuregs[19][17]), .B(_06825_), .Y(_06861_));
NOR_g _27810_ (.A(_09313_), .B(_06826_), .Y(_06862_));
NOR_g _27811_ (.A(_06861_), .B(_06862_), .Y(_01228_));
NOR_g _27812_ (.A(cpuregs[19][18]), .B(_06825_), .Y(_06863_));
NOR_g _27813_ (.A(_09325_), .B(_06826_), .Y(_06864_));
NOR_g _27814_ (.A(_06863_), .B(_06864_), .Y(_01229_));
NAND_g _27815_ (.A(_09338_), .B(_06825_), .Y(_06865_));
NAND_g _27816_ (.A(cpuregs[19][19]), .B(_06826_), .Y(_06866_));
NAND_g _27817_ (.A(_06865_), .B(_06866_), .Y(_01230_));
NAND_g _27818_ (.A(_09351_), .B(_06825_), .Y(_06867_));
NAND_g _27819_ (.A(cpuregs[19][20]), .B(_06826_), .Y(_06868_));
NAND_g _27820_ (.A(_06867_), .B(_06868_), .Y(_01231_));
NAND_g _27821_ (.A(_09364_), .B(_06825_), .Y(_06869_));
NAND_g _27822_ (.A(cpuregs[19][21]), .B(_06826_), .Y(_06870_));
NAND_g _27823_ (.A(_06869_), .B(_06870_), .Y(_01232_));
NAND_g _27824_ (.A(_09377_), .B(_06825_), .Y(_06871_));
NAND_g _27825_ (.A(cpuregs[19][22]), .B(_06826_), .Y(_06872_));
NAND_g _27826_ (.A(_06871_), .B(_06872_), .Y(_01233_));
NAND_g _27827_ (.A(_09390_), .B(_06825_), .Y(_06873_));
NAND_g _27828_ (.A(cpuregs[19][23]), .B(_06826_), .Y(_06874_));
NAND_g _27829_ (.A(_06873_), .B(_06874_), .Y(_01234_));
NAND_g _27830_ (.A(_09403_), .B(_06825_), .Y(_06875_));
NAND_g _27831_ (.A(cpuregs[19][24]), .B(_06826_), .Y(_06876_));
NAND_g _27832_ (.A(_06875_), .B(_06876_), .Y(_01235_));
NAND_g _27833_ (.A(_09416_), .B(_06825_), .Y(_06877_));
NAND_g _27834_ (.A(cpuregs[19][25]), .B(_06826_), .Y(_06878_));
NAND_g _27835_ (.A(_06877_), .B(_06878_), .Y(_01236_));
NAND_g _27836_ (.A(_09429_), .B(_06825_), .Y(_06879_));
NAND_g _27837_ (.A(cpuregs[19][26]), .B(_06826_), .Y(_06880_));
NAND_g _27838_ (.A(_06879_), .B(_06880_), .Y(_01237_));
NAND_g _27839_ (.A(_09442_), .B(_06825_), .Y(_06881_));
NAND_g _27840_ (.A(cpuregs[19][27]), .B(_06826_), .Y(_06882_));
NAND_g _27841_ (.A(_06881_), .B(_06882_), .Y(_01238_));
NAND_g _27842_ (.A(_09455_), .B(_06825_), .Y(_06883_));
NAND_g _27843_ (.A(cpuregs[19][28]), .B(_06826_), .Y(_06884_));
NAND_g _27844_ (.A(_06883_), .B(_06884_), .Y(_01239_));
NAND_g _27845_ (.A(_09468_), .B(_06825_), .Y(_06885_));
NAND_g _27846_ (.A(cpuregs[19][29]), .B(_06826_), .Y(_06886_));
NAND_g _27847_ (.A(_06885_), .B(_06886_), .Y(_01240_));
NAND_g _27848_ (.A(_09481_), .B(_06825_), .Y(_06887_));
NAND_g _27849_ (.A(cpuregs[19][30]), .B(_06826_), .Y(_06888_));
NAND_g _27850_ (.A(_06887_), .B(_06888_), .Y(_01241_));
NAND_g _27851_ (.A(_09493_), .B(_06825_), .Y(_06889_));
NAND_g _27852_ (.A(cpuregs[19][31]), .B(_06826_), .Y(_06890_));
NAND_g _27853_ (.A(_06889_), .B(_06890_), .Y(_01242_));
NAND_g _27854_ (.A(_14393_), .B(_00440_), .Y(_06891_));
NAND_g _27855_ (.A(decoded_imm_j[6]), .B(_14394_), .Y(_06892_));
NAND_g _27856_ (.A(_06891_), .B(_06892_), .Y(_01243_));
AND_g _27857_ (.A(_09825_), .B(_06692_), .Y(_06893_));
NAND_g _27858_ (.A(_09825_), .B(_06692_), .Y(_06894_));
NAND_g _27859_ (.A(cpuregs[25][0]), .B(_06894_), .Y(_06895_));
NAND_g _27860_ (.A(_09098_), .B(_06893_), .Y(_06896_));
NAND_g _27861_ (.A(_06895_), .B(_06896_), .Y(_01244_));
NAND_g _27862_ (.A(cpuregs[25][1]), .B(_06894_), .Y(_06897_));
NAND_g _27863_ (.A(_09109_), .B(_06893_), .Y(_06898_));
NAND_g _27864_ (.A(_06897_), .B(_06898_), .Y(_01245_));
NAND_g _27865_ (.A(cpuregs[25][2]), .B(_06894_), .Y(_06899_));
NAND_g _27866_ (.A(_09118_), .B(_06893_), .Y(_06900_));
NAND_g _27867_ (.A(_06899_), .B(_06900_), .Y(_01246_));
NAND_g _27868_ (.A(cpuregs[25][3]), .B(_06894_), .Y(_06901_));
NAND_g _27869_ (.A(_09131_), .B(_06893_), .Y(_06902_));
NAND_g _27870_ (.A(_06901_), .B(_06902_), .Y(_01247_));
NAND_g _27871_ (.A(cpuregs[25][4]), .B(_06894_), .Y(_06903_));
NAND_g _27872_ (.A(_09144_), .B(_06893_), .Y(_06904_));
NAND_g _27873_ (.A(_06903_), .B(_06904_), .Y(_01248_));
NAND_g _27874_ (.A(cpuregs[25][5]), .B(_06894_), .Y(_06905_));
NAND_g _27875_ (.A(_09157_), .B(_06893_), .Y(_06906_));
NAND_g _27876_ (.A(_06905_), .B(_06906_), .Y(_01249_));
NAND_g _27877_ (.A(cpuregs[25][6]), .B(_06894_), .Y(_06907_));
NAND_g _27878_ (.A(_09170_), .B(_06893_), .Y(_06908_));
NAND_g _27879_ (.A(_06907_), .B(_06908_), .Y(_01250_));
NAND_g _27880_ (.A(cpuregs[25][7]), .B(_06894_), .Y(_06909_));
NAND_g _27881_ (.A(_09183_), .B(_06893_), .Y(_06910_));
NAND_g _27882_ (.A(_06909_), .B(_06910_), .Y(_01251_));
NAND_g _27883_ (.A(cpuregs[25][8]), .B(_06894_), .Y(_06911_));
NAND_g _27884_ (.A(_09196_), .B(_06893_), .Y(_06912_));
NAND_g _27885_ (.A(_06911_), .B(_06912_), .Y(_01252_));
NAND_g _27886_ (.A(cpuregs[25][9]), .B(_06894_), .Y(_06913_));
NAND_g _27887_ (.A(_09209_), .B(_06893_), .Y(_06914_));
NAND_g _27888_ (.A(_06913_), .B(_06914_), .Y(_01253_));
NAND_g _27889_ (.A(cpuregs[25][10]), .B(_06894_), .Y(_06915_));
NAND_g _27890_ (.A(_09222_), .B(_06893_), .Y(_06916_));
NAND_g _27891_ (.A(_06915_), .B(_06916_), .Y(_01254_));
NAND_g _27892_ (.A(cpuregs[25][11]), .B(_06894_), .Y(_06917_));
NAND_g _27893_ (.A(_09235_), .B(_06893_), .Y(_06918_));
NAND_g _27894_ (.A(_06917_), .B(_06918_), .Y(_01255_));
NAND_g _27895_ (.A(cpuregs[25][12]), .B(_06894_), .Y(_06919_));
NAND_g _27896_ (.A(_09248_), .B(_06893_), .Y(_06920_));
NAND_g _27897_ (.A(_06919_), .B(_06920_), .Y(_01256_));
NAND_g _27898_ (.A(cpuregs[25][13]), .B(_06894_), .Y(_06921_));
NAND_g _27899_ (.A(_09261_), .B(_06893_), .Y(_06922_));
NAND_g _27900_ (.A(_06921_), .B(_06922_), .Y(_01257_));
NAND_g _27901_ (.A(cpuregs[25][14]), .B(_06894_), .Y(_06923_));
NAND_g _27902_ (.A(_09274_), .B(_06893_), .Y(_06924_));
NAND_g _27903_ (.A(_06923_), .B(_06924_), .Y(_01258_));
NAND_g _27904_ (.A(cpuregs[25][15]), .B(_06894_), .Y(_06925_));
NAND_g _27905_ (.A(_09287_), .B(_06893_), .Y(_06926_));
NAND_g _27906_ (.A(_06925_), .B(_06926_), .Y(_01259_));
NAND_g _27907_ (.A(cpuregs[25][16]), .B(_06894_), .Y(_06927_));
NAND_g _27908_ (.A(_09300_), .B(_06893_), .Y(_06928_));
NAND_g _27909_ (.A(_06927_), .B(_06928_), .Y(_01260_));
NOR_g _27910_ (.A(cpuregs[25][17]), .B(_06893_), .Y(_06929_));
NOR_g _27911_ (.A(_09313_), .B(_06894_), .Y(_06930_));
NOR_g _27912_ (.A(_06929_), .B(_06930_), .Y(_01261_));
NAND_g _27913_ (.A(cpuregs[25][18]), .B(_06894_), .Y(_06931_));
NAND_g _27914_ (.A(_09325_), .B(_06893_), .Y(_06932_));
NAND_g _27915_ (.A(_06931_), .B(_06932_), .Y(_01262_));
NAND_g _27916_ (.A(cpuregs[25][19]), .B(_06894_), .Y(_06933_));
NAND_g _27917_ (.A(_09338_), .B(_06893_), .Y(_06934_));
NAND_g _27918_ (.A(_06933_), .B(_06934_), .Y(_01263_));
NAND_g _27919_ (.A(cpuregs[25][20]), .B(_06894_), .Y(_06935_));
NAND_g _27920_ (.A(_09351_), .B(_06893_), .Y(_06936_));
NAND_g _27921_ (.A(_06935_), .B(_06936_), .Y(_01264_));
NAND_g _27922_ (.A(cpuregs[25][21]), .B(_06894_), .Y(_06937_));
NAND_g _27923_ (.A(_09364_), .B(_06893_), .Y(_06938_));
NAND_g _27924_ (.A(_06937_), .B(_06938_), .Y(_01265_));
NAND_g _27925_ (.A(cpuregs[25][22]), .B(_06894_), .Y(_06939_));
NAND_g _27926_ (.A(_09377_), .B(_06893_), .Y(_06940_));
NAND_g _27927_ (.A(_06939_), .B(_06940_), .Y(_01266_));
NAND_g _27928_ (.A(cpuregs[25][23]), .B(_06894_), .Y(_06941_));
NAND_g _27929_ (.A(_09390_), .B(_06893_), .Y(_06942_));
NAND_g _27930_ (.A(_06941_), .B(_06942_), .Y(_01267_));
NAND_g _27931_ (.A(cpuregs[25][24]), .B(_06894_), .Y(_06943_));
NAND_g _27932_ (.A(_09403_), .B(_06893_), .Y(_06944_));
NAND_g _27933_ (.A(_06943_), .B(_06944_), .Y(_01268_));
NAND_g _27934_ (.A(cpuregs[25][25]), .B(_06894_), .Y(_06945_));
NAND_g _27935_ (.A(_09416_), .B(_06893_), .Y(_06946_));
NAND_g _27936_ (.A(_06945_), .B(_06946_), .Y(_01269_));
NAND_g _27937_ (.A(cpuregs[25][26]), .B(_06894_), .Y(_06947_));
NAND_g _27938_ (.A(_09429_), .B(_06893_), .Y(_06948_));
NAND_g _27939_ (.A(_06947_), .B(_06948_), .Y(_01270_));
NAND_g _27940_ (.A(cpuregs[25][27]), .B(_06894_), .Y(_06949_));
NAND_g _27941_ (.A(_09442_), .B(_06893_), .Y(_06950_));
NAND_g _27942_ (.A(_06949_), .B(_06950_), .Y(_01271_));
NAND_g _27943_ (.A(cpuregs[25][28]), .B(_06894_), .Y(_06951_));
NAND_g _27944_ (.A(_09455_), .B(_06893_), .Y(_06952_));
NAND_g _27945_ (.A(_06951_), .B(_06952_), .Y(_01272_));
NAND_g _27946_ (.A(cpuregs[25][29]), .B(_06894_), .Y(_06953_));
NAND_g _27947_ (.A(_09468_), .B(_06893_), .Y(_06954_));
NAND_g _27948_ (.A(_06953_), .B(_06954_), .Y(_01273_));
NAND_g _27949_ (.A(cpuregs[25][30]), .B(_06894_), .Y(_06955_));
NAND_g _27950_ (.A(_09481_), .B(_06893_), .Y(_06956_));
NAND_g _27951_ (.A(_06955_), .B(_06956_), .Y(_01274_));
NAND_g _27952_ (.A(cpuregs[25][31]), .B(_06894_), .Y(_06957_));
NAND_g _27953_ (.A(_09493_), .B(_06893_), .Y(_06958_));
NAND_g _27954_ (.A(_06957_), .B(_06958_), .Y(_01275_));
AND_g _27955_ (.A(_09825_), .B(_02693_), .Y(_06959_));
NAND_g _27956_ (.A(_09825_), .B(_02693_), .Y(_06960_));
NAND_g _27957_ (.A(_09098_), .B(_06959_), .Y(_06961_));
NAND_g _27958_ (.A(cpuregs[9][0]), .B(_06960_), .Y(_06962_));
NAND_g _27959_ (.A(_06961_), .B(_06962_), .Y(_01276_));
NAND_g _27960_ (.A(_09109_), .B(_06959_), .Y(_06963_));
NAND_g _27961_ (.A(cpuregs[9][1]), .B(_06960_), .Y(_06964_));
NAND_g _27962_ (.A(_06963_), .B(_06964_), .Y(_01277_));
NAND_g _27963_ (.A(_09118_), .B(_06959_), .Y(_06965_));
NAND_g _27964_ (.A(cpuregs[9][2]), .B(_06960_), .Y(_06966_));
NAND_g _27965_ (.A(_06965_), .B(_06966_), .Y(_01278_));
NAND_g _27966_ (.A(_09131_), .B(_06959_), .Y(_06967_));
NAND_g _27967_ (.A(cpuregs[9][3]), .B(_06960_), .Y(_06968_));
NAND_g _27968_ (.A(_06967_), .B(_06968_), .Y(_01279_));
NAND_g _27969_ (.A(_09144_), .B(_06959_), .Y(_06969_));
NAND_g _27970_ (.A(cpuregs[9][4]), .B(_06960_), .Y(_06970_));
NAND_g _27971_ (.A(_06969_), .B(_06970_), .Y(_01280_));
NAND_g _27972_ (.A(_09157_), .B(_06959_), .Y(_06971_));
NAND_g _27973_ (.A(cpuregs[9][5]), .B(_06960_), .Y(_06972_));
NAND_g _27974_ (.A(_06971_), .B(_06972_), .Y(_01281_));
NAND_g _27975_ (.A(_09170_), .B(_06959_), .Y(_06973_));
NAND_g _27976_ (.A(cpuregs[9][6]), .B(_06960_), .Y(_06974_));
NAND_g _27977_ (.A(_06973_), .B(_06974_), .Y(_01282_));
NAND_g _27978_ (.A(_09183_), .B(_06959_), .Y(_06975_));
NAND_g _27979_ (.A(cpuregs[9][7]), .B(_06960_), .Y(_06976_));
NAND_g _27980_ (.A(_06975_), .B(_06976_), .Y(_01283_));
NAND_g _27981_ (.A(_09196_), .B(_06959_), .Y(_06977_));
NAND_g _27982_ (.A(cpuregs[9][8]), .B(_06960_), .Y(_06978_));
NAND_g _27983_ (.A(_06977_), .B(_06978_), .Y(_01284_));
NAND_g _27984_ (.A(_09209_), .B(_06959_), .Y(_06979_));
NAND_g _27985_ (.A(cpuregs[9][9]), .B(_06960_), .Y(_06980_));
NAND_g _27986_ (.A(_06979_), .B(_06980_), .Y(_01285_));
NAND_g _27987_ (.A(_09222_), .B(_06959_), .Y(_06981_));
NAND_g _27988_ (.A(cpuregs[9][10]), .B(_06960_), .Y(_06982_));
NAND_g _27989_ (.A(_06981_), .B(_06982_), .Y(_01286_));
NAND_g _27990_ (.A(_09235_), .B(_06959_), .Y(_06983_));
NAND_g _27991_ (.A(cpuregs[9][11]), .B(_06960_), .Y(_06984_));
NAND_g _27992_ (.A(_06983_), .B(_06984_), .Y(_01287_));
NAND_g _27993_ (.A(_09248_), .B(_06959_), .Y(_06985_));
NAND_g _27994_ (.A(cpuregs[9][12]), .B(_06960_), .Y(_06986_));
NAND_g _27995_ (.A(_06985_), .B(_06986_), .Y(_01288_));
NAND_g _27996_ (.A(_09261_), .B(_06959_), .Y(_06987_));
NAND_g _27997_ (.A(cpuregs[9][13]), .B(_06960_), .Y(_06988_));
NAND_g _27998_ (.A(_06987_), .B(_06988_), .Y(_01289_));
NAND_g _27999_ (.A(_09274_), .B(_06959_), .Y(_06989_));
NAND_g _28000_ (.A(cpuregs[9][14]), .B(_06960_), .Y(_06990_));
NAND_g _28001_ (.A(_06989_), .B(_06990_), .Y(_01290_));
NAND_g _28002_ (.A(_09287_), .B(_06959_), .Y(_06991_));
NAND_g _28003_ (.A(cpuregs[9][15]), .B(_06960_), .Y(_06992_));
NAND_g _28004_ (.A(_06991_), .B(_06992_), .Y(_01291_));
NOR_g _28005_ (.A(cpuregs[9][16]), .B(_06959_), .Y(_06993_));
NOR_g _28006_ (.A(_09300_), .B(_06960_), .Y(_06994_));
NOR_g _28007_ (.A(_06993_), .B(_06994_), .Y(_01292_));
NOR_g _28008_ (.A(cpuregs[9][17]), .B(_06959_), .Y(_06995_));
NOR_g _28009_ (.A(_09313_), .B(_06960_), .Y(_06996_));
NOR_g _28010_ (.A(_06995_), .B(_06996_), .Y(_01293_));
NAND_g _28011_ (.A(_09325_), .B(_06959_), .Y(_06997_));
NAND_g _28012_ (.A(cpuregs[9][18]), .B(_06960_), .Y(_06998_));
NAND_g _28013_ (.A(_06997_), .B(_06998_), .Y(_01294_));
NAND_g _28014_ (.A(_09338_), .B(_06959_), .Y(_06999_));
NAND_g _28015_ (.A(cpuregs[9][19]), .B(_06960_), .Y(_07000_));
NAND_g _28016_ (.A(_06999_), .B(_07000_), .Y(_01295_));
NAND_g _28017_ (.A(_09351_), .B(_06959_), .Y(_07001_));
NAND_g _28018_ (.A(cpuregs[9][20]), .B(_06960_), .Y(_07002_));
NAND_g _28019_ (.A(_07001_), .B(_07002_), .Y(_01296_));
NAND_g _28020_ (.A(_09364_), .B(_06959_), .Y(_07003_));
NAND_g _28021_ (.A(cpuregs[9][21]), .B(_06960_), .Y(_07004_));
NAND_g _28022_ (.A(_07003_), .B(_07004_), .Y(_01297_));
NAND_g _28023_ (.A(_09377_), .B(_06959_), .Y(_07005_));
NAND_g _28024_ (.A(cpuregs[9][22]), .B(_06960_), .Y(_07006_));
NAND_g _28025_ (.A(_07005_), .B(_07006_), .Y(_01298_));
NAND_g _28026_ (.A(_09390_), .B(_06959_), .Y(_07007_));
NAND_g _28027_ (.A(cpuregs[9][23]), .B(_06960_), .Y(_07008_));
NAND_g _28028_ (.A(_07007_), .B(_07008_), .Y(_01299_));
NAND_g _28029_ (.A(_09403_), .B(_06959_), .Y(_07009_));
NAND_g _28030_ (.A(cpuregs[9][24]), .B(_06960_), .Y(_07010_));
NAND_g _28031_ (.A(_07009_), .B(_07010_), .Y(_01300_));
NAND_g _28032_ (.A(_09416_), .B(_06959_), .Y(_07011_));
NAND_g _28033_ (.A(cpuregs[9][25]), .B(_06960_), .Y(_07012_));
NAND_g _28034_ (.A(_07011_), .B(_07012_), .Y(_01301_));
NAND_g _28035_ (.A(_09429_), .B(_06959_), .Y(_07013_));
NAND_g _28036_ (.A(cpuregs[9][26]), .B(_06960_), .Y(_07014_));
NAND_g _28037_ (.A(_07013_), .B(_07014_), .Y(_01302_));
NAND_g _28038_ (.A(_09442_), .B(_06959_), .Y(_07015_));
NAND_g _28039_ (.A(cpuregs[9][27]), .B(_06960_), .Y(_07016_));
NAND_g _28040_ (.A(_07015_), .B(_07016_), .Y(_01303_));
NAND_g _28041_ (.A(_09455_), .B(_06959_), .Y(_07017_));
NAND_g _28042_ (.A(cpuregs[9][28]), .B(_06960_), .Y(_07018_));
NAND_g _28043_ (.A(_07017_), .B(_07018_), .Y(_01304_));
NAND_g _28044_ (.A(_09468_), .B(_06959_), .Y(_07019_));
NAND_g _28045_ (.A(cpuregs[9][29]), .B(_06960_), .Y(_07020_));
NAND_g _28046_ (.A(_07019_), .B(_07020_), .Y(_01305_));
NAND_g _28047_ (.A(_09481_), .B(_06959_), .Y(_07021_));
NAND_g _28048_ (.A(cpuregs[9][30]), .B(_06960_), .Y(_07022_));
NAND_g _28049_ (.A(_07021_), .B(_07022_), .Y(_01306_));
NAND_g _28050_ (.A(_09493_), .B(_06959_), .Y(_07023_));
NAND_g _28051_ (.A(cpuregs[9][31]), .B(_06960_), .Y(_07024_));
NAND_g _28052_ (.A(_07023_), .B(_07024_), .Y(_01307_));
AND_g _28053_ (.A(_09825_), .B(_14285_), .Y(_07025_));
NAND_g _28054_ (.A(_09825_), .B(_14285_), .Y(_07026_));
NAND_g _28055_ (.A(_09098_), .B(_07025_), .Y(_07027_));
NAND_g _28056_ (.A(cpuregs[21][0]), .B(_07026_), .Y(_07028_));
NAND_g _28057_ (.A(_07027_), .B(_07028_), .Y(_01308_));
NAND_g _28058_ (.A(_09109_), .B(_07025_), .Y(_07029_));
NAND_g _28059_ (.A(cpuregs[21][1]), .B(_07026_), .Y(_07030_));
NAND_g _28060_ (.A(_07029_), .B(_07030_), .Y(_01309_));
NAND_g _28061_ (.A(_09118_), .B(_07025_), .Y(_07031_));
NAND_g _28062_ (.A(cpuregs[21][2]), .B(_07026_), .Y(_07032_));
NAND_g _28063_ (.A(_07031_), .B(_07032_), .Y(_01310_));
NAND_g _28064_ (.A(_09131_), .B(_07025_), .Y(_07033_));
NAND_g _28065_ (.A(cpuregs[21][3]), .B(_07026_), .Y(_07034_));
NAND_g _28066_ (.A(_07033_), .B(_07034_), .Y(_01311_));
NAND_g _28067_ (.A(_09144_), .B(_07025_), .Y(_07035_));
NAND_g _28068_ (.A(cpuregs[21][4]), .B(_07026_), .Y(_07036_));
NAND_g _28069_ (.A(_07035_), .B(_07036_), .Y(_01312_));
NAND_g _28070_ (.A(_09157_), .B(_07025_), .Y(_07037_));
NAND_g _28071_ (.A(cpuregs[21][5]), .B(_07026_), .Y(_07038_));
NAND_g _28072_ (.A(_07037_), .B(_07038_), .Y(_01313_));
NAND_g _28073_ (.A(_09170_), .B(_07025_), .Y(_07039_));
NAND_g _28074_ (.A(cpuregs[21][6]), .B(_07026_), .Y(_07040_));
NAND_g _28075_ (.A(_07039_), .B(_07040_), .Y(_01314_));
NAND_g _28076_ (.A(_09183_), .B(_07025_), .Y(_07041_));
NAND_g _28077_ (.A(cpuregs[21][7]), .B(_07026_), .Y(_07042_));
NAND_g _28078_ (.A(_07041_), .B(_07042_), .Y(_01315_));
NAND_g _28079_ (.A(_09196_), .B(_07025_), .Y(_07043_));
NAND_g _28080_ (.A(cpuregs[21][8]), .B(_07026_), .Y(_07044_));
NAND_g _28081_ (.A(_07043_), .B(_07044_), .Y(_01316_));
NAND_g _28082_ (.A(_09209_), .B(_07025_), .Y(_07045_));
NAND_g _28083_ (.A(cpuregs[21][9]), .B(_07026_), .Y(_07046_));
NAND_g _28084_ (.A(_07045_), .B(_07046_), .Y(_01317_));
NAND_g _28085_ (.A(_09222_), .B(_07025_), .Y(_07047_));
NAND_g _28086_ (.A(cpuregs[21][10]), .B(_07026_), .Y(_07048_));
NAND_g _28087_ (.A(_07047_), .B(_07048_), .Y(_01318_));
NAND_g _28088_ (.A(_09235_), .B(_07025_), .Y(_07049_));
NAND_g _28089_ (.A(cpuregs[21][11]), .B(_07026_), .Y(_07050_));
NAND_g _28090_ (.A(_07049_), .B(_07050_), .Y(_01319_));
NAND_g _28091_ (.A(_09248_), .B(_07025_), .Y(_07051_));
NAND_g _28092_ (.A(cpuregs[21][12]), .B(_07026_), .Y(_07052_));
NAND_g _28093_ (.A(_07051_), .B(_07052_), .Y(_01320_));
NAND_g _28094_ (.A(_09261_), .B(_07025_), .Y(_07053_));
NAND_g _28095_ (.A(cpuregs[21][13]), .B(_07026_), .Y(_07054_));
NAND_g _28096_ (.A(_07053_), .B(_07054_), .Y(_01321_));
NAND_g _28097_ (.A(_09274_), .B(_07025_), .Y(_07055_));
NAND_g _28098_ (.A(cpuregs[21][14]), .B(_07026_), .Y(_07056_));
NAND_g _28099_ (.A(_07055_), .B(_07056_), .Y(_01322_));
NAND_g _28100_ (.A(_09287_), .B(_07025_), .Y(_07057_));
NAND_g _28101_ (.A(cpuregs[21][15]), .B(_07026_), .Y(_07058_));
NAND_g _28102_ (.A(_07057_), .B(_07058_), .Y(_01323_));
NAND_g _28103_ (.A(_09300_), .B(_07025_), .Y(_07059_));
NAND_g _28104_ (.A(cpuregs[21][16]), .B(_07026_), .Y(_07060_));
NAND_g _28105_ (.A(_07059_), .B(_07060_), .Y(_01324_));
NOR_g _28106_ (.A(cpuregs[21][17]), .B(_07025_), .Y(_07061_));
NOR_g _28107_ (.A(_09313_), .B(_07026_), .Y(_07062_));
NOR_g _28108_ (.A(_07061_), .B(_07062_), .Y(_01325_));
NOR_g _28109_ (.A(cpuregs[21][18]), .B(_07025_), .Y(_07063_));
NOR_g _28110_ (.A(_09325_), .B(_07026_), .Y(_07064_));
NOR_g _28111_ (.A(_07063_), .B(_07064_), .Y(_01326_));
NAND_g _28112_ (.A(_09338_), .B(_07025_), .Y(_07065_));
NAND_g _28113_ (.A(cpuregs[21][19]), .B(_07026_), .Y(_07066_));
NAND_g _28114_ (.A(_07065_), .B(_07066_), .Y(_01327_));
NAND_g _28115_ (.A(_09351_), .B(_07025_), .Y(_07067_));
NAND_g _28116_ (.A(cpuregs[21][20]), .B(_07026_), .Y(_07068_));
NAND_g _28117_ (.A(_07067_), .B(_07068_), .Y(_01328_));
NAND_g _28118_ (.A(_09364_), .B(_07025_), .Y(_07069_));
NAND_g _28119_ (.A(cpuregs[21][21]), .B(_07026_), .Y(_07070_));
NAND_g _28120_ (.A(_07069_), .B(_07070_), .Y(_01329_));
NAND_g _28121_ (.A(_09377_), .B(_07025_), .Y(_07071_));
NAND_g _28122_ (.A(cpuregs[21][22]), .B(_07026_), .Y(_07072_));
NAND_g _28123_ (.A(_07071_), .B(_07072_), .Y(_01330_));
NAND_g _28124_ (.A(_09390_), .B(_07025_), .Y(_07073_));
NAND_g _28125_ (.A(cpuregs[21][23]), .B(_07026_), .Y(_07074_));
NAND_g _28126_ (.A(_07073_), .B(_07074_), .Y(_01331_));
NAND_g _28127_ (.A(_09403_), .B(_07025_), .Y(_07075_));
NAND_g _28128_ (.A(cpuregs[21][24]), .B(_07026_), .Y(_07076_));
NAND_g _28129_ (.A(_07075_), .B(_07076_), .Y(_01332_));
NAND_g _28130_ (.A(_09416_), .B(_07025_), .Y(_07077_));
NAND_g _28131_ (.A(cpuregs[21][25]), .B(_07026_), .Y(_07078_));
NAND_g _28132_ (.A(_07077_), .B(_07078_), .Y(_01333_));
NAND_g _28133_ (.A(_09429_), .B(_07025_), .Y(_07079_));
NAND_g _28134_ (.A(cpuregs[21][26]), .B(_07026_), .Y(_07080_));
NAND_g _28135_ (.A(_07079_), .B(_07080_), .Y(_01334_));
NAND_g _28136_ (.A(_09442_), .B(_07025_), .Y(_07081_));
NAND_g _28137_ (.A(cpuregs[21][27]), .B(_07026_), .Y(_07082_));
NAND_g _28138_ (.A(_07081_), .B(_07082_), .Y(_01335_));
NAND_g _28139_ (.A(_09455_), .B(_07025_), .Y(_07083_));
NAND_g _28140_ (.A(cpuregs[21][28]), .B(_07026_), .Y(_07084_));
NAND_g _28141_ (.A(_07083_), .B(_07084_), .Y(_01336_));
NAND_g _28142_ (.A(_09468_), .B(_07025_), .Y(_07085_));
NAND_g _28143_ (.A(cpuregs[21][29]), .B(_07026_), .Y(_07086_));
NAND_g _28144_ (.A(_07085_), .B(_07086_), .Y(_01337_));
NAND_g _28145_ (.A(_09481_), .B(_07025_), .Y(_07087_));
NAND_g _28146_ (.A(cpuregs[21][30]), .B(_07026_), .Y(_07088_));
NAND_g _28147_ (.A(_07087_), .B(_07088_), .Y(_01338_));
NAND_g _28148_ (.A(_09493_), .B(_07025_), .Y(_07089_));
NAND_g _28149_ (.A(cpuregs[21][31]), .B(_07026_), .Y(_07090_));
NAND_g _28150_ (.A(_07089_), .B(_07090_), .Y(_01339_));
AND_g _28151_ (.A(_09496_), .B(_02494_), .Y(_07091_));
NAND_g _28152_ (.A(_09496_), .B(_02494_), .Y(_07092_));
NAND_g _28153_ (.A(_09098_), .B(_07091_), .Y(_07093_));
NAND_g _28154_ (.A(cpuregs[6][0]), .B(_07092_), .Y(_07094_));
NAND_g _28155_ (.A(_07093_), .B(_07094_), .Y(_01340_));
NAND_g _28156_ (.A(_09109_), .B(_07091_), .Y(_07095_));
NAND_g _28157_ (.A(cpuregs[6][1]), .B(_07092_), .Y(_07096_));
NAND_g _28158_ (.A(_07095_), .B(_07096_), .Y(_01341_));
NAND_g _28159_ (.A(_09118_), .B(_07091_), .Y(_07097_));
NAND_g _28160_ (.A(cpuregs[6][2]), .B(_07092_), .Y(_07098_));
NAND_g _28161_ (.A(_07097_), .B(_07098_), .Y(_01342_));
NAND_g _28162_ (.A(_09131_), .B(_07091_), .Y(_07099_));
NAND_g _28163_ (.A(cpuregs[6][3]), .B(_07092_), .Y(_07100_));
NAND_g _28164_ (.A(_07099_), .B(_07100_), .Y(_01343_));
NAND_g _28165_ (.A(_09144_), .B(_07091_), .Y(_07101_));
NAND_g _28166_ (.A(cpuregs[6][4]), .B(_07092_), .Y(_07102_));
NAND_g _28167_ (.A(_07101_), .B(_07102_), .Y(_01344_));
NAND_g _28168_ (.A(_09157_), .B(_07091_), .Y(_07103_));
NAND_g _28169_ (.A(cpuregs[6][5]), .B(_07092_), .Y(_07104_));
NAND_g _28170_ (.A(_07103_), .B(_07104_), .Y(_01345_));
NAND_g _28171_ (.A(_09170_), .B(_07091_), .Y(_07105_));
NAND_g _28172_ (.A(cpuregs[6][6]), .B(_07092_), .Y(_07106_));
NAND_g _28173_ (.A(_07105_), .B(_07106_), .Y(_01346_));
NAND_g _28174_ (.A(_09183_), .B(_07091_), .Y(_07107_));
NAND_g _28175_ (.A(cpuregs[6][7]), .B(_07092_), .Y(_07108_));
NAND_g _28176_ (.A(_07107_), .B(_07108_), .Y(_01347_));
NAND_g _28177_ (.A(_09196_), .B(_07091_), .Y(_07109_));
NAND_g _28178_ (.A(cpuregs[6][8]), .B(_07092_), .Y(_07110_));
NAND_g _28179_ (.A(_07109_), .B(_07110_), .Y(_01348_));
NAND_g _28180_ (.A(_09209_), .B(_07091_), .Y(_07111_));
NAND_g _28181_ (.A(cpuregs[6][9]), .B(_07092_), .Y(_07112_));
NAND_g _28182_ (.A(_07111_), .B(_07112_), .Y(_01349_));
NAND_g _28183_ (.A(_09222_), .B(_07091_), .Y(_07113_));
NAND_g _28184_ (.A(cpuregs[6][10]), .B(_07092_), .Y(_07114_));
NAND_g _28185_ (.A(_07113_), .B(_07114_), .Y(_01350_));
NAND_g _28186_ (.A(_09235_), .B(_07091_), .Y(_07115_));
NAND_g _28187_ (.A(cpuregs[6][11]), .B(_07092_), .Y(_07116_));
NAND_g _28188_ (.A(_07115_), .B(_07116_), .Y(_01351_));
NAND_g _28189_ (.A(_09248_), .B(_07091_), .Y(_07117_));
NAND_g _28190_ (.A(cpuregs[6][12]), .B(_07092_), .Y(_07118_));
NAND_g _28191_ (.A(_07117_), .B(_07118_), .Y(_01352_));
NAND_g _28192_ (.A(_09261_), .B(_07091_), .Y(_07119_));
NAND_g _28193_ (.A(cpuregs[6][13]), .B(_07092_), .Y(_07120_));
NAND_g _28194_ (.A(_07119_), .B(_07120_), .Y(_01353_));
NAND_g _28195_ (.A(_09274_), .B(_07091_), .Y(_07121_));
NAND_g _28196_ (.A(cpuregs[6][14]), .B(_07092_), .Y(_07122_));
NAND_g _28197_ (.A(_07121_), .B(_07122_), .Y(_01354_));
NAND_g _28198_ (.A(_09287_), .B(_07091_), .Y(_07123_));
NAND_g _28199_ (.A(cpuregs[6][15]), .B(_07092_), .Y(_07124_));
NAND_g _28200_ (.A(_07123_), .B(_07124_), .Y(_01355_));
NAND_g _28201_ (.A(_09300_), .B(_07091_), .Y(_07125_));
NAND_g _28202_ (.A(cpuregs[6][16]), .B(_07092_), .Y(_07126_));
NAND_g _28203_ (.A(_07125_), .B(_07126_), .Y(_01356_));
NOR_g _28204_ (.A(cpuregs[6][17]), .B(_07091_), .Y(_07127_));
NOR_g _28205_ (.A(_09313_), .B(_07092_), .Y(_07128_));
NOR_g _28206_ (.A(_07127_), .B(_07128_), .Y(_01357_));
AND_g _28207_ (.A(_09012_), .B(_07092_), .Y(_07129_));
NOR_g _28208_ (.A(_09325_), .B(_07092_), .Y(_07130_));
NOR_g _28209_ (.A(_07129_), .B(_07130_), .Y(_01358_));
NAND_g _28210_ (.A(_09338_), .B(_07091_), .Y(_07131_));
NAND_g _28211_ (.A(cpuregs[6][19]), .B(_07092_), .Y(_07132_));
NAND_g _28212_ (.A(_07131_), .B(_07132_), .Y(_01359_));
NAND_g _28213_ (.A(_09351_), .B(_07091_), .Y(_07133_));
NAND_g _28214_ (.A(cpuregs[6][20]), .B(_07092_), .Y(_07134_));
NAND_g _28215_ (.A(_07133_), .B(_07134_), .Y(_01360_));
NAND_g _28216_ (.A(_09364_), .B(_07091_), .Y(_07135_));
NAND_g _28217_ (.A(cpuregs[6][21]), .B(_07092_), .Y(_07136_));
NAND_g _28218_ (.A(_07135_), .B(_07136_), .Y(_01361_));
NAND_g _28219_ (.A(_09377_), .B(_07091_), .Y(_07137_));
NAND_g _28220_ (.A(cpuregs[6][22]), .B(_07092_), .Y(_07138_));
NAND_g _28221_ (.A(_07137_), .B(_07138_), .Y(_01362_));
NAND_g _28222_ (.A(_09390_), .B(_07091_), .Y(_07139_));
NAND_g _28223_ (.A(cpuregs[6][23]), .B(_07092_), .Y(_07140_));
NAND_g _28224_ (.A(_07139_), .B(_07140_), .Y(_01363_));
NAND_g _28225_ (.A(_09403_), .B(_07091_), .Y(_07141_));
NAND_g _28226_ (.A(cpuregs[6][24]), .B(_07092_), .Y(_07142_));
NAND_g _28227_ (.A(_07141_), .B(_07142_), .Y(_01364_));
NAND_g _28228_ (.A(_09416_), .B(_07091_), .Y(_07143_));
NAND_g _28229_ (.A(cpuregs[6][25]), .B(_07092_), .Y(_07144_));
NAND_g _28230_ (.A(_07143_), .B(_07144_), .Y(_01365_));
NAND_g _28231_ (.A(_09429_), .B(_07091_), .Y(_07145_));
NAND_g _28232_ (.A(cpuregs[6][26]), .B(_07092_), .Y(_07146_));
NAND_g _28233_ (.A(_07145_), .B(_07146_), .Y(_01366_));
NAND_g _28234_ (.A(_09442_), .B(_07091_), .Y(_07147_));
NAND_g _28235_ (.A(cpuregs[6][27]), .B(_07092_), .Y(_07148_));
NAND_g _28236_ (.A(_07147_), .B(_07148_), .Y(_01367_));
NAND_g _28237_ (.A(_09455_), .B(_07091_), .Y(_07149_));
NAND_g _28238_ (.A(cpuregs[6][28]), .B(_07092_), .Y(_07150_));
NAND_g _28239_ (.A(_07149_), .B(_07150_), .Y(_01368_));
NAND_g _28240_ (.A(_09468_), .B(_07091_), .Y(_07151_));
NAND_g _28241_ (.A(cpuregs[6][29]), .B(_07092_), .Y(_07152_));
NAND_g _28242_ (.A(_07151_), .B(_07152_), .Y(_01369_));
NAND_g _28243_ (.A(_09481_), .B(_07091_), .Y(_07153_));
NAND_g _28244_ (.A(cpuregs[6][30]), .B(_07092_), .Y(_07154_));
NAND_g _28245_ (.A(_07153_), .B(_07154_), .Y(_01370_));
NAND_g _28246_ (.A(_09493_), .B(_07091_), .Y(_07155_));
NAND_g _28247_ (.A(cpuregs[6][31]), .B(_07092_), .Y(_07156_));
NAND_g _28248_ (.A(_07155_), .B(_07156_), .Y(_01371_));
AND_g _28249_ (.A(_09496_), .B(_02693_), .Y(_07157_));
NAND_g _28250_ (.A(_09496_), .B(_02693_), .Y(_07158_));
NAND_g _28251_ (.A(_09098_), .B(_07157_), .Y(_07159_));
NAND_g _28252_ (.A(cpuregs[10][0]), .B(_07158_), .Y(_07160_));
NAND_g _28253_ (.A(_07159_), .B(_07160_), .Y(_01372_));
NAND_g _28254_ (.A(_09109_), .B(_07157_), .Y(_07161_));
NAND_g _28255_ (.A(cpuregs[10][1]), .B(_07158_), .Y(_07162_));
NAND_g _28256_ (.A(_07161_), .B(_07162_), .Y(_01373_));
NAND_g _28257_ (.A(_09118_), .B(_07157_), .Y(_07163_));
NAND_g _28258_ (.A(cpuregs[10][2]), .B(_07158_), .Y(_07164_));
NAND_g _28259_ (.A(_07163_), .B(_07164_), .Y(_01374_));
NAND_g _28260_ (.A(_09131_), .B(_07157_), .Y(_07165_));
NAND_g _28261_ (.A(cpuregs[10][3]), .B(_07158_), .Y(_07166_));
NAND_g _28262_ (.A(_07165_), .B(_07166_), .Y(_01375_));
NAND_g _28263_ (.A(_09144_), .B(_07157_), .Y(_07167_));
NAND_g _28264_ (.A(cpuregs[10][4]), .B(_07158_), .Y(_07168_));
NAND_g _28265_ (.A(_07167_), .B(_07168_), .Y(_01376_));
NAND_g _28266_ (.A(_09157_), .B(_07157_), .Y(_07169_));
NAND_g _28267_ (.A(cpuregs[10][5]), .B(_07158_), .Y(_07170_));
NAND_g _28268_ (.A(_07169_), .B(_07170_), .Y(_01377_));
NAND_g _28269_ (.A(_09170_), .B(_07157_), .Y(_07171_));
NAND_g _28270_ (.A(cpuregs[10][6]), .B(_07158_), .Y(_07172_));
NAND_g _28271_ (.A(_07171_), .B(_07172_), .Y(_01378_));
NAND_g _28272_ (.A(_09183_), .B(_07157_), .Y(_07173_));
NAND_g _28273_ (.A(cpuregs[10][7]), .B(_07158_), .Y(_07174_));
NAND_g _28274_ (.A(_07173_), .B(_07174_), .Y(_01379_));
NAND_g _28275_ (.A(_09196_), .B(_07157_), .Y(_07175_));
NAND_g _28276_ (.A(cpuregs[10][8]), .B(_07158_), .Y(_07176_));
NAND_g _28277_ (.A(_07175_), .B(_07176_), .Y(_01380_));
NAND_g _28278_ (.A(_09209_), .B(_07157_), .Y(_07177_));
NAND_g _28279_ (.A(cpuregs[10][9]), .B(_07158_), .Y(_07178_));
NAND_g _28280_ (.A(_07177_), .B(_07178_), .Y(_01381_));
NAND_g _28281_ (.A(_09222_), .B(_07157_), .Y(_07179_));
NAND_g _28282_ (.A(cpuregs[10][10]), .B(_07158_), .Y(_07180_));
NAND_g _28283_ (.A(_07179_), .B(_07180_), .Y(_01382_));
NAND_g _28284_ (.A(_09235_), .B(_07157_), .Y(_07181_));
NAND_g _28285_ (.A(cpuregs[10][11]), .B(_07158_), .Y(_07182_));
NAND_g _28286_ (.A(_07181_), .B(_07182_), .Y(_01383_));
NAND_g _28287_ (.A(_09248_), .B(_07157_), .Y(_07183_));
NAND_g _28288_ (.A(cpuregs[10][12]), .B(_07158_), .Y(_07184_));
NAND_g _28289_ (.A(_07183_), .B(_07184_), .Y(_01384_));
NAND_g _28290_ (.A(_09261_), .B(_07157_), .Y(_07185_));
NAND_g _28291_ (.A(cpuregs[10][13]), .B(_07158_), .Y(_07186_));
NAND_g _28292_ (.A(_07185_), .B(_07186_), .Y(_01385_));
NAND_g _28293_ (.A(_09274_), .B(_07157_), .Y(_07187_));
NAND_g _28294_ (.A(cpuregs[10][14]), .B(_07158_), .Y(_07188_));
NAND_g _28295_ (.A(_07187_), .B(_07188_), .Y(_01386_));
NAND_g _28296_ (.A(_09287_), .B(_07157_), .Y(_07189_));
NAND_g _28297_ (.A(cpuregs[10][15]), .B(_07158_), .Y(_07190_));
NAND_g _28298_ (.A(_07189_), .B(_07190_), .Y(_01387_));
NOR_g _28299_ (.A(cpuregs[10][16]), .B(_07157_), .Y(_07191_));
NOR_g _28300_ (.A(_09300_), .B(_07158_), .Y(_07192_));
NOR_g _28301_ (.A(_07191_), .B(_07192_), .Y(_01388_));
NOR_g _28302_ (.A(cpuregs[10][17]), .B(_07157_), .Y(_07193_));
NOR_g _28303_ (.A(_09313_), .B(_07158_), .Y(_07194_));
NOR_g _28304_ (.A(_07193_), .B(_07194_), .Y(_01389_));
NAND_g _28305_ (.A(_09325_), .B(_07157_), .Y(_07195_));
NAND_g _28306_ (.A(cpuregs[10][18]), .B(_07158_), .Y(_07196_));
NAND_g _28307_ (.A(_07195_), .B(_07196_), .Y(_01390_));
NAND_g _28308_ (.A(_09338_), .B(_07157_), .Y(_07197_));
NAND_g _28309_ (.A(cpuregs[10][19]), .B(_07158_), .Y(_07198_));
NAND_g _28310_ (.A(_07197_), .B(_07198_), .Y(_01391_));
NAND_g _28311_ (.A(_09351_), .B(_07157_), .Y(_07199_));
NAND_g _28312_ (.A(cpuregs[10][20]), .B(_07158_), .Y(_07200_));
NAND_g _28313_ (.A(_07199_), .B(_07200_), .Y(_01392_));
NAND_g _28314_ (.A(_09364_), .B(_07157_), .Y(_07201_));
NAND_g _28315_ (.A(cpuregs[10][21]), .B(_07158_), .Y(_07202_));
NAND_g _28316_ (.A(_07201_), .B(_07202_), .Y(_01393_));
NAND_g _28317_ (.A(_09377_), .B(_07157_), .Y(_07203_));
NAND_g _28318_ (.A(cpuregs[10][22]), .B(_07158_), .Y(_07204_));
NAND_g _28319_ (.A(_07203_), .B(_07204_), .Y(_01394_));
NAND_g _28320_ (.A(_09390_), .B(_07157_), .Y(_07205_));
NAND_g _28321_ (.A(cpuregs[10][23]), .B(_07158_), .Y(_07206_));
NAND_g _28322_ (.A(_07205_), .B(_07206_), .Y(_01395_));
NAND_g _28323_ (.A(_09403_), .B(_07157_), .Y(_07207_));
NAND_g _28324_ (.A(cpuregs[10][24]), .B(_07158_), .Y(_07208_));
NAND_g _28325_ (.A(_07207_), .B(_07208_), .Y(_01396_));
NAND_g _28326_ (.A(_09416_), .B(_07157_), .Y(_07209_));
NAND_g _28327_ (.A(cpuregs[10][25]), .B(_07158_), .Y(_07210_));
NAND_g _28328_ (.A(_07209_), .B(_07210_), .Y(_01397_));
NAND_g _28329_ (.A(_09429_), .B(_07157_), .Y(_07211_));
NAND_g _28330_ (.A(cpuregs[10][26]), .B(_07158_), .Y(_07212_));
NAND_g _28331_ (.A(_07211_), .B(_07212_), .Y(_01398_));
NAND_g _28332_ (.A(_09442_), .B(_07157_), .Y(_07213_));
NAND_g _28333_ (.A(cpuregs[10][27]), .B(_07158_), .Y(_07214_));
NAND_g _28334_ (.A(_07213_), .B(_07214_), .Y(_01399_));
NAND_g _28335_ (.A(_09455_), .B(_07157_), .Y(_07215_));
NAND_g _28336_ (.A(cpuregs[10][28]), .B(_07158_), .Y(_07216_));
NAND_g _28337_ (.A(_07215_), .B(_07216_), .Y(_01400_));
NAND_g _28338_ (.A(_09468_), .B(_07157_), .Y(_07217_));
NAND_g _28339_ (.A(cpuregs[10][29]), .B(_07158_), .Y(_07218_));
NAND_g _28340_ (.A(_07217_), .B(_07218_), .Y(_01401_));
NAND_g _28341_ (.A(_09481_), .B(_07157_), .Y(_07219_));
NAND_g _28342_ (.A(cpuregs[10][30]), .B(_07158_), .Y(_07220_));
NAND_g _28343_ (.A(_07219_), .B(_07220_), .Y(_01402_));
NAND_g _28344_ (.A(_09493_), .B(_07157_), .Y(_07221_));
NAND_g _28345_ (.A(cpuregs[10][31]), .B(_07158_), .Y(_07222_));
NAND_g _28346_ (.A(_07221_), .B(_07222_), .Y(_01403_));
AND_g _28347_ (.A(_14286_), .B(_06692_), .Y(_07223_));
NAND_g _28348_ (.A(_14286_), .B(_06692_), .Y(_07224_));
NAND_g _28349_ (.A(cpuregs[24][0]), .B(_07224_), .Y(_07225_));
NAND_g _28350_ (.A(_09098_), .B(_07223_), .Y(_07226_));
NAND_g _28351_ (.A(_07225_), .B(_07226_), .Y(_01404_));
NAND_g _28352_ (.A(cpuregs[24][1]), .B(_07224_), .Y(_07227_));
NAND_g _28353_ (.A(_09109_), .B(_07223_), .Y(_07228_));
NAND_g _28354_ (.A(_07227_), .B(_07228_), .Y(_01405_));
NAND_g _28355_ (.A(cpuregs[24][2]), .B(_07224_), .Y(_07229_));
NAND_g _28356_ (.A(_09118_), .B(_07223_), .Y(_07230_));
NAND_g _28357_ (.A(_07229_), .B(_07230_), .Y(_01406_));
NAND_g _28358_ (.A(cpuregs[24][3]), .B(_07224_), .Y(_07231_));
NAND_g _28359_ (.A(_09131_), .B(_07223_), .Y(_07232_));
NAND_g _28360_ (.A(_07231_), .B(_07232_), .Y(_01407_));
NAND_g _28361_ (.A(cpuregs[24][4]), .B(_07224_), .Y(_07233_));
NAND_g _28362_ (.A(_09144_), .B(_07223_), .Y(_07234_));
NAND_g _28363_ (.A(_07233_), .B(_07234_), .Y(_01408_));
NAND_g _28364_ (.A(cpuregs[24][5]), .B(_07224_), .Y(_07235_));
NAND_g _28365_ (.A(_09157_), .B(_07223_), .Y(_07236_));
NAND_g _28366_ (.A(_07235_), .B(_07236_), .Y(_01409_));
NAND_g _28367_ (.A(cpuregs[24][6]), .B(_07224_), .Y(_07237_));
NAND_g _28368_ (.A(_09170_), .B(_07223_), .Y(_07238_));
NAND_g _28369_ (.A(_07237_), .B(_07238_), .Y(_01410_));
NAND_g _28370_ (.A(cpuregs[24][7]), .B(_07224_), .Y(_07239_));
NAND_g _28371_ (.A(_09183_), .B(_07223_), .Y(_07240_));
NAND_g _28372_ (.A(_07239_), .B(_07240_), .Y(_01411_));
NAND_g _28373_ (.A(cpuregs[24][8]), .B(_07224_), .Y(_07241_));
NAND_g _28374_ (.A(_09196_), .B(_07223_), .Y(_07242_));
NAND_g _28375_ (.A(_07241_), .B(_07242_), .Y(_01412_));
NAND_g _28376_ (.A(cpuregs[24][9]), .B(_07224_), .Y(_07243_));
NAND_g _28377_ (.A(_09209_), .B(_07223_), .Y(_07244_));
NAND_g _28378_ (.A(_07243_), .B(_07244_), .Y(_01413_));
NAND_g _28379_ (.A(cpuregs[24][10]), .B(_07224_), .Y(_07245_));
NAND_g _28380_ (.A(_09222_), .B(_07223_), .Y(_07246_));
NAND_g _28381_ (.A(_07245_), .B(_07246_), .Y(_01414_));
NAND_g _28382_ (.A(cpuregs[24][11]), .B(_07224_), .Y(_07247_));
NAND_g _28383_ (.A(_09235_), .B(_07223_), .Y(_07248_));
NAND_g _28384_ (.A(_07247_), .B(_07248_), .Y(_01415_));
NAND_g _28385_ (.A(cpuregs[24][12]), .B(_07224_), .Y(_07249_));
NAND_g _28386_ (.A(_09248_), .B(_07223_), .Y(_07250_));
NAND_g _28387_ (.A(_07249_), .B(_07250_), .Y(_01416_));
NAND_g _28388_ (.A(cpuregs[24][13]), .B(_07224_), .Y(_07251_));
NAND_g _28389_ (.A(_09261_), .B(_07223_), .Y(_07252_));
NAND_g _28390_ (.A(_07251_), .B(_07252_), .Y(_01417_));
NAND_g _28391_ (.A(cpuregs[24][14]), .B(_07224_), .Y(_07253_));
NAND_g _28392_ (.A(_09274_), .B(_07223_), .Y(_07254_));
NAND_g _28393_ (.A(_07253_), .B(_07254_), .Y(_01418_));
NAND_g _28394_ (.A(cpuregs[24][15]), .B(_07224_), .Y(_07255_));
NAND_g _28395_ (.A(_09287_), .B(_07223_), .Y(_07256_));
NAND_g _28396_ (.A(_07255_), .B(_07256_), .Y(_01419_));
NAND_g _28397_ (.A(cpuregs[24][16]), .B(_07224_), .Y(_07257_));
NAND_g _28398_ (.A(_09300_), .B(_07223_), .Y(_07258_));
NAND_g _28399_ (.A(_07257_), .B(_07258_), .Y(_01420_));
NOR_g _28400_ (.A(cpuregs[24][17]), .B(_07223_), .Y(_07259_));
NOR_g _28401_ (.A(_09313_), .B(_07224_), .Y(_07260_));
NOR_g _28402_ (.A(_07259_), .B(_07260_), .Y(_01421_));
NAND_g _28403_ (.A(cpuregs[24][18]), .B(_07224_), .Y(_07261_));
NAND_g _28404_ (.A(_09325_), .B(_07223_), .Y(_07262_));
NAND_g _28405_ (.A(_07261_), .B(_07262_), .Y(_01422_));
NAND_g _28406_ (.A(cpuregs[24][19]), .B(_07224_), .Y(_07263_));
NAND_g _28407_ (.A(_09338_), .B(_07223_), .Y(_07264_));
NAND_g _28408_ (.A(_07263_), .B(_07264_), .Y(_01423_));
NAND_g _28409_ (.A(cpuregs[24][20]), .B(_07224_), .Y(_07265_));
NAND_g _28410_ (.A(_09351_), .B(_07223_), .Y(_07266_));
NAND_g _28411_ (.A(_07265_), .B(_07266_), .Y(_01424_));
NAND_g _28412_ (.A(cpuregs[24][21]), .B(_07224_), .Y(_07267_));
NAND_g _28413_ (.A(_09364_), .B(_07223_), .Y(_07268_));
NAND_g _28414_ (.A(_07267_), .B(_07268_), .Y(_01425_));
NAND_g _28415_ (.A(cpuregs[24][22]), .B(_07224_), .Y(_07269_));
NAND_g _28416_ (.A(_09377_), .B(_07223_), .Y(_07270_));
NAND_g _28417_ (.A(_07269_), .B(_07270_), .Y(_01426_));
NAND_g _28418_ (.A(cpuregs[24][23]), .B(_07224_), .Y(_07271_));
NAND_g _28419_ (.A(_09390_), .B(_07223_), .Y(_07272_));
NAND_g _28420_ (.A(_07271_), .B(_07272_), .Y(_01427_));
NAND_g _28421_ (.A(cpuregs[24][24]), .B(_07224_), .Y(_07273_));
NAND_g _28422_ (.A(_09403_), .B(_07223_), .Y(_07274_));
NAND_g _28423_ (.A(_07273_), .B(_07274_), .Y(_01428_));
NAND_g _28424_ (.A(cpuregs[24][25]), .B(_07224_), .Y(_07275_));
NAND_g _28425_ (.A(_09416_), .B(_07223_), .Y(_07276_));
NAND_g _28426_ (.A(_07275_), .B(_07276_), .Y(_01429_));
NAND_g _28427_ (.A(cpuregs[24][26]), .B(_07224_), .Y(_07277_));
NAND_g _28428_ (.A(_09429_), .B(_07223_), .Y(_07278_));
NAND_g _28429_ (.A(_07277_), .B(_07278_), .Y(_01430_));
NAND_g _28430_ (.A(cpuregs[24][27]), .B(_07224_), .Y(_07279_));
NAND_g _28431_ (.A(_09442_), .B(_07223_), .Y(_07280_));
NAND_g _28432_ (.A(_07279_), .B(_07280_), .Y(_01431_));
NAND_g _28433_ (.A(cpuregs[24][28]), .B(_07224_), .Y(_07281_));
NAND_g _28434_ (.A(_09455_), .B(_07223_), .Y(_07282_));
NAND_g _28435_ (.A(_07281_), .B(_07282_), .Y(_01432_));
NAND_g _28436_ (.A(cpuregs[24][29]), .B(_07224_), .Y(_07283_));
NAND_g _28437_ (.A(_09468_), .B(_07223_), .Y(_07284_));
NAND_g _28438_ (.A(_07283_), .B(_07284_), .Y(_01433_));
NAND_g _28439_ (.A(cpuregs[24][30]), .B(_07224_), .Y(_07285_));
NAND_g _28440_ (.A(_09481_), .B(_07223_), .Y(_07286_));
NAND_g _28441_ (.A(_07285_), .B(_07286_), .Y(_01434_));
NAND_g _28442_ (.A(cpuregs[24][31]), .B(_07224_), .Y(_07287_));
NAND_g _28443_ (.A(_09493_), .B(_07223_), .Y(_07288_));
NAND_g _28444_ (.A(_07287_), .B(_07288_), .Y(_01435_));
NAND_g _28445_ (.A(_14393_), .B(_00445_), .Y(_07289_));
NAND_g _28446_ (.A(decoded_imm_j[31]), .B(_14394_), .Y(_07290_));
NAND_g _28447_ (.A(_07289_), .B(_07290_), .Y(_01436_));
NAND_g _28448_ (.A(_14393_), .B(_00439_), .Y(_07291_));
NAND_g _28449_ (.A(decoded_imm_j[5]), .B(_14394_), .Y(_07292_));
NAND_g _28450_ (.A(_07291_), .B(_07292_), .Y(_01437_));
NAND_g _28451_ (.A(_14393_), .B(_00441_), .Y(_07293_));
NAND_g _28452_ (.A(decoded_imm_j[7]), .B(_14394_), .Y(_07294_));
NAND_g _28453_ (.A(_07293_), .B(_07294_), .Y(_01438_));
AND_g _28454_ (.A(_14286_), .B(_02760_), .Y(_07295_));
NAND_g _28455_ (.A(_14286_), .B(_02760_), .Y(_07296_));
NAND_g _28456_ (.A(_09098_), .B(_07295_), .Y(_07297_));
NAND_g _28457_ (.A(cpuregs[16][0]), .B(_07296_), .Y(_07298_));
NAND_g _28458_ (.A(_07297_), .B(_07298_), .Y(_01439_));
NAND_g _28459_ (.A(_09109_), .B(_07295_), .Y(_07299_));
NAND_g _28460_ (.A(cpuregs[16][1]), .B(_07296_), .Y(_07300_));
NAND_g _28461_ (.A(_07299_), .B(_07300_), .Y(_01440_));
NAND_g _28462_ (.A(_09118_), .B(_07295_), .Y(_07301_));
NAND_g _28463_ (.A(cpuregs[16][2]), .B(_07296_), .Y(_07302_));
NAND_g _28464_ (.A(_07301_), .B(_07302_), .Y(_01441_));
NAND_g _28465_ (.A(_09131_), .B(_07295_), .Y(_07303_));
NAND_g _28466_ (.A(cpuregs[16][3]), .B(_07296_), .Y(_07304_));
NAND_g _28467_ (.A(_07303_), .B(_07304_), .Y(_01442_));
NAND_g _28468_ (.A(_09144_), .B(_07295_), .Y(_07305_));
NAND_g _28469_ (.A(cpuregs[16][4]), .B(_07296_), .Y(_07306_));
NAND_g _28470_ (.A(_07305_), .B(_07306_), .Y(_01443_));
NAND_g _28471_ (.A(_09157_), .B(_07295_), .Y(_07307_));
NAND_g _28472_ (.A(cpuregs[16][5]), .B(_07296_), .Y(_07308_));
NAND_g _28473_ (.A(_07307_), .B(_07308_), .Y(_01444_));
NAND_g _28474_ (.A(_09170_), .B(_07295_), .Y(_07309_));
NAND_g _28475_ (.A(cpuregs[16][6]), .B(_07296_), .Y(_07310_));
NAND_g _28476_ (.A(_07309_), .B(_07310_), .Y(_01445_));
NAND_g _28477_ (.A(_09183_), .B(_07295_), .Y(_07311_));
NAND_g _28478_ (.A(cpuregs[16][7]), .B(_07296_), .Y(_07312_));
NAND_g _28479_ (.A(_07311_), .B(_07312_), .Y(_01446_));
NAND_g _28480_ (.A(_09196_), .B(_07295_), .Y(_07313_));
NAND_g _28481_ (.A(cpuregs[16][8]), .B(_07296_), .Y(_07314_));
NAND_g _28482_ (.A(_07313_), .B(_07314_), .Y(_01447_));
NAND_g _28483_ (.A(_09209_), .B(_07295_), .Y(_07315_));
NAND_g _28484_ (.A(cpuregs[16][9]), .B(_07296_), .Y(_07316_));
NAND_g _28485_ (.A(_07315_), .B(_07316_), .Y(_01448_));
NAND_g _28486_ (.A(_09222_), .B(_07295_), .Y(_07317_));
NAND_g _28487_ (.A(cpuregs[16][10]), .B(_07296_), .Y(_07318_));
NAND_g _28488_ (.A(_07317_), .B(_07318_), .Y(_01449_));
NAND_g _28489_ (.A(_09235_), .B(_07295_), .Y(_07319_));
NAND_g _28490_ (.A(cpuregs[16][11]), .B(_07296_), .Y(_07320_));
NAND_g _28491_ (.A(_07319_), .B(_07320_), .Y(_01450_));
NAND_g _28492_ (.A(_09248_), .B(_07295_), .Y(_07321_));
NAND_g _28493_ (.A(cpuregs[16][12]), .B(_07296_), .Y(_07322_));
NAND_g _28494_ (.A(_07321_), .B(_07322_), .Y(_01451_));
NAND_g _28495_ (.A(_09261_), .B(_07295_), .Y(_07323_));
NAND_g _28496_ (.A(cpuregs[16][13]), .B(_07296_), .Y(_07324_));
NAND_g _28497_ (.A(_07323_), .B(_07324_), .Y(_01452_));
NAND_g _28498_ (.A(_09274_), .B(_07295_), .Y(_07325_));
NAND_g _28499_ (.A(cpuregs[16][14]), .B(_07296_), .Y(_07326_));
NAND_g _28500_ (.A(_07325_), .B(_07326_), .Y(_01453_));
NAND_g _28501_ (.A(_09287_), .B(_07295_), .Y(_07327_));
NAND_g _28502_ (.A(cpuregs[16][15]), .B(_07296_), .Y(_07328_));
NAND_g _28503_ (.A(_07327_), .B(_07328_), .Y(_01454_));
NAND_g _28504_ (.A(_09300_), .B(_07295_), .Y(_07329_));
NAND_g _28505_ (.A(cpuregs[16][16]), .B(_07296_), .Y(_07330_));
NAND_g _28506_ (.A(_07329_), .B(_07330_), .Y(_01455_));
NOR_g _28507_ (.A(cpuregs[16][17]), .B(_07295_), .Y(_07331_));
NOR_g _28508_ (.A(_09313_), .B(_07296_), .Y(_07332_));
NOR_g _28509_ (.A(_07331_), .B(_07332_), .Y(_01456_));
NOR_g _28510_ (.A(cpuregs[16][18]), .B(_07295_), .Y(_07333_));
NOR_g _28511_ (.A(_09325_), .B(_07296_), .Y(_07334_));
NOR_g _28512_ (.A(_07333_), .B(_07334_), .Y(_01457_));
NAND_g _28513_ (.A(_09338_), .B(_07295_), .Y(_07335_));
NAND_g _28514_ (.A(cpuregs[16][19]), .B(_07296_), .Y(_07336_));
NAND_g _28515_ (.A(_07335_), .B(_07336_), .Y(_01458_));
NAND_g _28516_ (.A(_09351_), .B(_07295_), .Y(_07337_));
NAND_g _28517_ (.A(cpuregs[16][20]), .B(_07296_), .Y(_07338_));
NAND_g _28518_ (.A(_07337_), .B(_07338_), .Y(_01459_));
NAND_g _28519_ (.A(_09364_), .B(_07295_), .Y(_07339_));
NAND_g _28520_ (.A(cpuregs[16][21]), .B(_07296_), .Y(_07340_));
NAND_g _28521_ (.A(_07339_), .B(_07340_), .Y(_01460_));
NAND_g _28522_ (.A(_09377_), .B(_07295_), .Y(_07341_));
NAND_g _28523_ (.A(cpuregs[16][22]), .B(_07296_), .Y(_07342_));
NAND_g _28524_ (.A(_07341_), .B(_07342_), .Y(_01461_));
NAND_g _28525_ (.A(_09390_), .B(_07295_), .Y(_07343_));
NAND_g _28526_ (.A(cpuregs[16][23]), .B(_07296_), .Y(_07344_));
NAND_g _28527_ (.A(_07343_), .B(_07344_), .Y(_01462_));
NAND_g _28528_ (.A(_09403_), .B(_07295_), .Y(_07345_));
NAND_g _28529_ (.A(cpuregs[16][24]), .B(_07296_), .Y(_07346_));
NAND_g _28530_ (.A(_07345_), .B(_07346_), .Y(_01463_));
NAND_g _28531_ (.A(_09416_), .B(_07295_), .Y(_07347_));
NAND_g _28532_ (.A(cpuregs[16][25]), .B(_07296_), .Y(_07348_));
NAND_g _28533_ (.A(_07347_), .B(_07348_), .Y(_01464_));
NAND_g _28534_ (.A(_09429_), .B(_07295_), .Y(_07349_));
NAND_g _28535_ (.A(cpuregs[16][26]), .B(_07296_), .Y(_07350_));
NAND_g _28536_ (.A(_07349_), .B(_07350_), .Y(_01465_));
NAND_g _28537_ (.A(_09442_), .B(_07295_), .Y(_07351_));
NAND_g _28538_ (.A(cpuregs[16][27]), .B(_07296_), .Y(_07352_));
NAND_g _28539_ (.A(_07351_), .B(_07352_), .Y(_01466_));
NAND_g _28540_ (.A(_09455_), .B(_07295_), .Y(_07353_));
NAND_g _28541_ (.A(cpuregs[16][28]), .B(_07296_), .Y(_07354_));
NAND_g _28542_ (.A(_07353_), .B(_07354_), .Y(_01467_));
NAND_g _28543_ (.A(_09468_), .B(_07295_), .Y(_07355_));
NAND_g _28544_ (.A(cpuregs[16][29]), .B(_07296_), .Y(_07356_));
NAND_g _28545_ (.A(_07355_), .B(_07356_), .Y(_01468_));
NAND_g _28546_ (.A(_09481_), .B(_07295_), .Y(_07357_));
NAND_g _28547_ (.A(cpuregs[16][30]), .B(_07296_), .Y(_07358_));
NAND_g _28548_ (.A(_07357_), .B(_07358_), .Y(_01469_));
NAND_g _28549_ (.A(_09493_), .B(_07295_), .Y(_07359_));
NAND_g _28550_ (.A(cpuregs[16][31]), .B(_07296_), .Y(_07360_));
NAND_g _28551_ (.A(_07359_), .B(_07360_), .Y(_01470_));
AND_g _28552_ (.A(_09085_), .B(_06692_), .Y(_07361_));
NAND_g _28553_ (.A(_09085_), .B(_06692_), .Y(_07362_));
NAND_g _28554_ (.A(cpuregs[27][0]), .B(_07362_), .Y(_07363_));
NAND_g _28555_ (.A(_09098_), .B(_07361_), .Y(_07364_));
NAND_g _28556_ (.A(_07363_), .B(_07364_), .Y(_01471_));
NAND_g _28557_ (.A(cpuregs[27][1]), .B(_07362_), .Y(_07365_));
NAND_g _28558_ (.A(_09109_), .B(_07361_), .Y(_07366_));
NAND_g _28559_ (.A(_07365_), .B(_07366_), .Y(_01472_));
NAND_g _28560_ (.A(cpuregs[27][2]), .B(_07362_), .Y(_07367_));
NAND_g _28561_ (.A(_09118_), .B(_07361_), .Y(_07368_));
NAND_g _28562_ (.A(_07367_), .B(_07368_), .Y(_01473_));
NAND_g _28563_ (.A(cpuregs[27][3]), .B(_07362_), .Y(_07369_));
NAND_g _28564_ (.A(_09131_), .B(_07361_), .Y(_07370_));
NAND_g _28565_ (.A(_07369_), .B(_07370_), .Y(_01474_));
NAND_g _28566_ (.A(cpuregs[27][4]), .B(_07362_), .Y(_07371_));
NAND_g _28567_ (.A(_09144_), .B(_07361_), .Y(_07372_));
NAND_g _28568_ (.A(_07371_), .B(_07372_), .Y(_01475_));
NAND_g _28569_ (.A(cpuregs[27][5]), .B(_07362_), .Y(_07373_));
NAND_g _28570_ (.A(_09157_), .B(_07361_), .Y(_07374_));
NAND_g _28571_ (.A(_07373_), .B(_07374_), .Y(_01476_));
NAND_g _28572_ (.A(cpuregs[27][6]), .B(_07362_), .Y(_07375_));
NAND_g _28573_ (.A(_09170_), .B(_07361_), .Y(_07376_));
NAND_g _28574_ (.A(_07375_), .B(_07376_), .Y(_01477_));
NAND_g _28575_ (.A(cpuregs[27][7]), .B(_07362_), .Y(_07377_));
NAND_g _28576_ (.A(_09183_), .B(_07361_), .Y(_07378_));
NAND_g _28577_ (.A(_07377_), .B(_07378_), .Y(_01478_));
NAND_g _28578_ (.A(cpuregs[27][8]), .B(_07362_), .Y(_07379_));
NAND_g _28579_ (.A(_09196_), .B(_07361_), .Y(_07380_));
NAND_g _28580_ (.A(_07379_), .B(_07380_), .Y(_01479_));
NAND_g _28581_ (.A(cpuregs[27][9]), .B(_07362_), .Y(_07381_));
NAND_g _28582_ (.A(_09209_), .B(_07361_), .Y(_07382_));
NAND_g _28583_ (.A(_07381_), .B(_07382_), .Y(_01480_));
NAND_g _28584_ (.A(cpuregs[27][10]), .B(_07362_), .Y(_07383_));
NAND_g _28585_ (.A(_09222_), .B(_07361_), .Y(_07384_));
NAND_g _28586_ (.A(_07383_), .B(_07384_), .Y(_01481_));
NAND_g _28587_ (.A(cpuregs[27][11]), .B(_07362_), .Y(_07385_));
NAND_g _28588_ (.A(_09235_), .B(_07361_), .Y(_07386_));
NAND_g _28589_ (.A(_07385_), .B(_07386_), .Y(_01482_));
NAND_g _28590_ (.A(cpuregs[27][12]), .B(_07362_), .Y(_07387_));
NAND_g _28591_ (.A(_09248_), .B(_07361_), .Y(_07388_));
NAND_g _28592_ (.A(_07387_), .B(_07388_), .Y(_01483_));
NAND_g _28593_ (.A(cpuregs[27][13]), .B(_07362_), .Y(_07389_));
NAND_g _28594_ (.A(_09261_), .B(_07361_), .Y(_07390_));
NAND_g _28595_ (.A(_07389_), .B(_07390_), .Y(_01484_));
NAND_g _28596_ (.A(cpuregs[27][14]), .B(_07362_), .Y(_07391_));
NAND_g _28597_ (.A(_09274_), .B(_07361_), .Y(_07392_));
NAND_g _28598_ (.A(_07391_), .B(_07392_), .Y(_01485_));
NAND_g _28599_ (.A(cpuregs[27][15]), .B(_07362_), .Y(_07393_));
NAND_g _28600_ (.A(_09287_), .B(_07361_), .Y(_07394_));
NAND_g _28601_ (.A(_07393_), .B(_07394_), .Y(_01486_));
NAND_g _28602_ (.A(cpuregs[27][16]), .B(_07362_), .Y(_07395_));
NAND_g _28603_ (.A(_09300_), .B(_07361_), .Y(_07396_));
NAND_g _28604_ (.A(_07395_), .B(_07396_), .Y(_01487_));
NOR_g _28605_ (.A(cpuregs[27][17]), .B(_07361_), .Y(_07397_));
NOR_g _28606_ (.A(_09313_), .B(_07362_), .Y(_07398_));
NOR_g _28607_ (.A(_07397_), .B(_07398_), .Y(_01488_));
NAND_g _28608_ (.A(cpuregs[27][18]), .B(_07362_), .Y(_07399_));
NAND_g _28609_ (.A(_09325_), .B(_07361_), .Y(_07400_));
NAND_g _28610_ (.A(_07399_), .B(_07400_), .Y(_01489_));
NAND_g _28611_ (.A(cpuregs[27][19]), .B(_07362_), .Y(_07401_));
NAND_g _28612_ (.A(_09338_), .B(_07361_), .Y(_07402_));
NAND_g _28613_ (.A(_07401_), .B(_07402_), .Y(_01490_));
NAND_g _28614_ (.A(cpuregs[27][20]), .B(_07362_), .Y(_07403_));
NAND_g _28615_ (.A(_09351_), .B(_07361_), .Y(_07404_));
NAND_g _28616_ (.A(_07403_), .B(_07404_), .Y(_01491_));
NAND_g _28617_ (.A(cpuregs[27][21]), .B(_07362_), .Y(_07405_));
NAND_g _28618_ (.A(_09364_), .B(_07361_), .Y(_07406_));
NAND_g _28619_ (.A(_07405_), .B(_07406_), .Y(_01492_));
NAND_g _28620_ (.A(cpuregs[27][22]), .B(_07362_), .Y(_07407_));
NAND_g _28621_ (.A(_09377_), .B(_07361_), .Y(_07408_));
NAND_g _28622_ (.A(_07407_), .B(_07408_), .Y(_01493_));
NAND_g _28623_ (.A(cpuregs[27][23]), .B(_07362_), .Y(_07409_));
NAND_g _28624_ (.A(_09390_), .B(_07361_), .Y(_07410_));
NAND_g _28625_ (.A(_07409_), .B(_07410_), .Y(_01494_));
NAND_g _28626_ (.A(cpuregs[27][24]), .B(_07362_), .Y(_07411_));
NAND_g _28627_ (.A(_09403_), .B(_07361_), .Y(_07412_));
NAND_g _28628_ (.A(_07411_), .B(_07412_), .Y(_01495_));
NAND_g _28629_ (.A(cpuregs[27][25]), .B(_07362_), .Y(_07413_));
NAND_g _28630_ (.A(_09416_), .B(_07361_), .Y(_07414_));
NAND_g _28631_ (.A(_07413_), .B(_07414_), .Y(_01496_));
NAND_g _28632_ (.A(cpuregs[27][26]), .B(_07362_), .Y(_07415_));
NAND_g _28633_ (.A(_09429_), .B(_07361_), .Y(_07416_));
NAND_g _28634_ (.A(_07415_), .B(_07416_), .Y(_01497_));
NAND_g _28635_ (.A(cpuregs[27][27]), .B(_07362_), .Y(_07417_));
NAND_g _28636_ (.A(_09442_), .B(_07361_), .Y(_07418_));
NAND_g _28637_ (.A(_07417_), .B(_07418_), .Y(_01498_));
NAND_g _28638_ (.A(cpuregs[27][28]), .B(_07362_), .Y(_07419_));
NAND_g _28639_ (.A(_09455_), .B(_07361_), .Y(_07420_));
NAND_g _28640_ (.A(_07419_), .B(_07420_), .Y(_01499_));
NAND_g _28641_ (.A(cpuregs[27][29]), .B(_07362_), .Y(_07421_));
NAND_g _28642_ (.A(_09468_), .B(_07361_), .Y(_07422_));
NAND_g _28643_ (.A(_07421_), .B(_07422_), .Y(_01500_));
NAND_g _28644_ (.A(cpuregs[27][30]), .B(_07362_), .Y(_07423_));
NAND_g _28645_ (.A(_09481_), .B(_07361_), .Y(_07424_));
NAND_g _28646_ (.A(_07423_), .B(_07424_), .Y(_01501_));
NAND_g _28647_ (.A(cpuregs[27][31]), .B(_07362_), .Y(_07425_));
NAND_g _28648_ (.A(_09493_), .B(_07361_), .Y(_07426_));
NAND_g _28649_ (.A(_07425_), .B(_07426_), .Y(_01502_));
AND_g _28650_ (.A(_09499_), .B(_14286_), .Y(_07427_));
NAND_g _28651_ (.A(_09499_), .B(_14286_), .Y(_07428_));
NAND_g _28652_ (.A(_09098_), .B(_07427_), .Y(_07429_));
NAND_g _28653_ (.A(cpuregs[28][0]), .B(_07428_), .Y(_07430_));
NAND_g _28654_ (.A(_07429_), .B(_07430_), .Y(_01503_));
NAND_g _28655_ (.A(_09109_), .B(_07427_), .Y(_07431_));
NAND_g _28656_ (.A(cpuregs[28][1]), .B(_07428_), .Y(_07432_));
NAND_g _28657_ (.A(_07431_), .B(_07432_), .Y(_01504_));
NAND_g _28658_ (.A(_09118_), .B(_07427_), .Y(_07433_));
NAND_g _28659_ (.A(cpuregs[28][2]), .B(_07428_), .Y(_07434_));
NAND_g _28660_ (.A(_07433_), .B(_07434_), .Y(_01505_));
NAND_g _28661_ (.A(_09131_), .B(_07427_), .Y(_07435_));
NAND_g _28662_ (.A(cpuregs[28][3]), .B(_07428_), .Y(_07436_));
NAND_g _28663_ (.A(_07435_), .B(_07436_), .Y(_01506_));
NAND_g _28664_ (.A(_09144_), .B(_07427_), .Y(_07437_));
NAND_g _28665_ (.A(cpuregs[28][4]), .B(_07428_), .Y(_07438_));
NAND_g _28666_ (.A(_07437_), .B(_07438_), .Y(_01507_));
NAND_g _28667_ (.A(_09157_), .B(_07427_), .Y(_07439_));
NAND_g _28668_ (.A(cpuregs[28][5]), .B(_07428_), .Y(_07440_));
NAND_g _28669_ (.A(_07439_), .B(_07440_), .Y(_01508_));
NAND_g _28670_ (.A(_09170_), .B(_07427_), .Y(_07441_));
NAND_g _28671_ (.A(cpuregs[28][6]), .B(_07428_), .Y(_07442_));
NAND_g _28672_ (.A(_07441_), .B(_07442_), .Y(_01509_));
NAND_g _28673_ (.A(_09183_), .B(_07427_), .Y(_07443_));
NAND_g _28674_ (.A(cpuregs[28][7]), .B(_07428_), .Y(_07444_));
NAND_g _28675_ (.A(_07443_), .B(_07444_), .Y(_01510_));
NAND_g _28676_ (.A(_09196_), .B(_07427_), .Y(_07445_));
NAND_g _28677_ (.A(cpuregs[28][8]), .B(_07428_), .Y(_07446_));
NAND_g _28678_ (.A(_07445_), .B(_07446_), .Y(_01511_));
NAND_g _28679_ (.A(_09209_), .B(_07427_), .Y(_07447_));
NAND_g _28680_ (.A(cpuregs[28][9]), .B(_07428_), .Y(_07448_));
NAND_g _28681_ (.A(_07447_), .B(_07448_), .Y(_01512_));
NAND_g _28682_ (.A(_09222_), .B(_07427_), .Y(_07449_));
NAND_g _28683_ (.A(cpuregs[28][10]), .B(_07428_), .Y(_07450_));
NAND_g _28684_ (.A(_07449_), .B(_07450_), .Y(_01513_));
NAND_g _28685_ (.A(_09235_), .B(_07427_), .Y(_07451_));
NAND_g _28686_ (.A(cpuregs[28][11]), .B(_07428_), .Y(_07452_));
NAND_g _28687_ (.A(_07451_), .B(_07452_), .Y(_01514_));
NAND_g _28688_ (.A(_09248_), .B(_07427_), .Y(_07453_));
NAND_g _28689_ (.A(cpuregs[28][12]), .B(_07428_), .Y(_07454_));
NAND_g _28690_ (.A(_07453_), .B(_07454_), .Y(_01515_));
NAND_g _28691_ (.A(_09261_), .B(_07427_), .Y(_07455_));
NAND_g _28692_ (.A(cpuregs[28][13]), .B(_07428_), .Y(_07456_));
NAND_g _28693_ (.A(_07455_), .B(_07456_), .Y(_01516_));
NAND_g _28694_ (.A(_09274_), .B(_07427_), .Y(_07457_));
NAND_g _28695_ (.A(cpuregs[28][14]), .B(_07428_), .Y(_07458_));
NAND_g _28696_ (.A(_07457_), .B(_07458_), .Y(_01517_));
NAND_g _28697_ (.A(_09287_), .B(_07427_), .Y(_07459_));
NAND_g _28698_ (.A(cpuregs[28][15]), .B(_07428_), .Y(_07460_));
NAND_g _28699_ (.A(_07459_), .B(_07460_), .Y(_01518_));
NAND_g _28700_ (.A(_09300_), .B(_07427_), .Y(_07461_));
NAND_g _28701_ (.A(cpuregs[28][16]), .B(_07428_), .Y(_07462_));
NAND_g _28702_ (.A(_07461_), .B(_07462_), .Y(_01519_));
NOR_g _28703_ (.A(cpuregs[28][17]), .B(_07427_), .Y(_07463_));
NOR_g _28704_ (.A(_09313_), .B(_07428_), .Y(_07464_));
NOR_g _28705_ (.A(_07463_), .B(_07464_), .Y(_01520_));
NAND_g _28706_ (.A(_09325_), .B(_07427_), .Y(_07465_));
NAND_g _28707_ (.A(cpuregs[28][18]), .B(_07428_), .Y(_07466_));
NAND_g _28708_ (.A(_07465_), .B(_07466_), .Y(_01521_));
NAND_g _28709_ (.A(_09338_), .B(_07427_), .Y(_07467_));
NAND_g _28710_ (.A(cpuregs[28][19]), .B(_07428_), .Y(_07468_));
NAND_g _28711_ (.A(_07467_), .B(_07468_), .Y(_01522_));
NAND_g _28712_ (.A(_09351_), .B(_07427_), .Y(_07469_));
NAND_g _28713_ (.A(cpuregs[28][20]), .B(_07428_), .Y(_07470_));
NAND_g _28714_ (.A(_07469_), .B(_07470_), .Y(_01523_));
NAND_g _28715_ (.A(_09364_), .B(_07427_), .Y(_07471_));
NAND_g _28716_ (.A(cpuregs[28][21]), .B(_07428_), .Y(_07472_));
NAND_g _28717_ (.A(_07471_), .B(_07472_), .Y(_01524_));
NAND_g _28718_ (.A(_09377_), .B(_07427_), .Y(_07473_));
NAND_g _28719_ (.A(cpuregs[28][22]), .B(_07428_), .Y(_07474_));
NAND_g _28720_ (.A(_07473_), .B(_07474_), .Y(_01525_));
NAND_g _28721_ (.A(_09390_), .B(_07427_), .Y(_07475_));
NAND_g _28722_ (.A(cpuregs[28][23]), .B(_07428_), .Y(_07476_));
NAND_g _28723_ (.A(_07475_), .B(_07476_), .Y(_01526_));
NAND_g _28724_ (.A(_09403_), .B(_07427_), .Y(_07477_));
NAND_g _28725_ (.A(cpuregs[28][24]), .B(_07428_), .Y(_07478_));
NAND_g _28726_ (.A(_07477_), .B(_07478_), .Y(_01527_));
NAND_g _28727_ (.A(_09416_), .B(_07427_), .Y(_07479_));
NAND_g _28728_ (.A(cpuregs[28][25]), .B(_07428_), .Y(_07480_));
NAND_g _28729_ (.A(_07479_), .B(_07480_), .Y(_01528_));
NAND_g _28730_ (.A(_09429_), .B(_07427_), .Y(_07481_));
NAND_g _28731_ (.A(cpuregs[28][26]), .B(_07428_), .Y(_07482_));
NAND_g _28732_ (.A(_07481_), .B(_07482_), .Y(_01529_));
NAND_g _28733_ (.A(_09442_), .B(_07427_), .Y(_07483_));
NAND_g _28734_ (.A(cpuregs[28][27]), .B(_07428_), .Y(_07484_));
NAND_g _28735_ (.A(_07483_), .B(_07484_), .Y(_01530_));
NAND_g _28736_ (.A(_09455_), .B(_07427_), .Y(_07485_));
NAND_g _28737_ (.A(cpuregs[28][28]), .B(_07428_), .Y(_07486_));
NAND_g _28738_ (.A(_07485_), .B(_07486_), .Y(_01531_));
NAND_g _28739_ (.A(_09468_), .B(_07427_), .Y(_07487_));
NAND_g _28740_ (.A(cpuregs[28][29]), .B(_07428_), .Y(_07488_));
NAND_g _28741_ (.A(_07487_), .B(_07488_), .Y(_01532_));
NAND_g _28742_ (.A(_09481_), .B(_07427_), .Y(_07489_));
NAND_g _28743_ (.A(cpuregs[28][30]), .B(_07428_), .Y(_07490_));
NAND_g _28744_ (.A(_07489_), .B(_07490_), .Y(_01533_));
NAND_g _28745_ (.A(_09493_), .B(_07427_), .Y(_07491_));
NAND_g _28746_ (.A(cpuregs[28][31]), .B(_07428_), .Y(_07492_));
NAND_g _28747_ (.A(_07491_), .B(_07492_), .Y(_01534_));
NAND_g _28748_ (.A(_08798_), .B(_10717_), .Y(_00003_));
NAND_g _28749_ (.A(_08797_), .B(_10718_), .Y(_00004_));
NAND_g _28750_ (.A(_08858_), .B(_10722_), .Y(_00001_));
NAND_g _28751_ (.A(is_compare), .B(_14212_), .Y(_07493_));
AND_g _28752_ (.A(_09023_), .B(_10742_), .Y(_07494_));
NOT_g _28753_ (.A(_07494_), .Y(_07495_));
NOR_g _28754_ (.A(instr_or), .B(instr_ori), .Y(_07496_));
NOR_g _28755_ (.A(instr_and), .B(instr_andi), .Y(_07497_));
NOR_g _28756_ (.A(_14075_), .B(_07497_), .Y(_07498_));
NAND_g _28757_ (.A(_14075_), .B(_07495_), .Y(_07499_));
AND_g _28758_ (.A(_07496_), .B(_07499_), .Y(_07500_));
NOR_g _28759_ (.A(_14074_), .B(_07500_), .Y(_07501_));
NOR_g _28760_ (.A(_07498_), .B(_07501_), .Y(_07502_));
NAND_g _28761_ (.A(_07493_), .B(_07502_), .Y(alu_out[0]));
NAND_g _28762_ (.A(_08794_), .B(_14075_), .Y(_07503_));
NAND_g _28763_ (.A(instr_sub), .B(_14077_), .Y(_07504_));
AND_g _28764_ (.A(_07503_), .B(_07504_), .Y(_07505_));
NAND_g _28765_ (.A(_14072_), .B(_07505_), .Y(_07506_));
NOR_g _28766_ (.A(_14072_), .B(_07505_), .Y(_07507_));
NOR_g _28767_ (.A(_09023_), .B(_07507_), .Y(_07508_));
NAND_g _28768_ (.A(_07506_), .B(_07508_), .Y(_07509_));
NAND_g _28769_ (.A(_10743_), .B(_14072_), .Y(_07510_));
NOR_g _28770_ (.A(_14071_), .B(_07497_), .Y(_07511_));
NOR_g _28771_ (.A(_14069_), .B(_07496_), .Y(_07512_));
NOR_g _28772_ (.A(_07511_), .B(_07512_), .Y(_07513_));
AND_g _28773_ (.A(_07510_), .B(_07513_), .Y(_07514_));
NAND_g _28774_ (.A(_07509_), .B(_07514_), .Y(alu_out[1]));
NOR_g _28775_ (.A(_08794_), .B(_14079_), .Y(_07515_));
NOR_g _28776_ (.A(_14069_), .B(_14075_), .Y(_07516_));
NOR_g _28777_ (.A(_14070_), .B(_07516_), .Y(_07517_));
NOR_g _28778_ (.A(instr_sub), .B(_07517_), .Y(_07518_));
NOR_g _28779_ (.A(_07515_), .B(_07518_), .Y(_07519_));
XNOR_g _28780_ (.A(_14066_), .B(_07519_), .Y(_07520_));
NAND_g _28781_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07520_), .Y(_07521_));
NAND_g _28782_ (.A(_10743_), .B(_14066_), .Y(_07522_));
NOR_g _28783_ (.A(_14063_), .B(_07496_), .Y(_07523_));
NOR_g _28784_ (.A(_14065_), .B(_07497_), .Y(_07524_));
NOR_g _28785_ (.A(_07523_), .B(_07524_), .Y(_07525_));
AND_g _28786_ (.A(_07522_), .B(_07525_), .Y(_07526_));
NAND_g _28787_ (.A(_07521_), .B(_07526_), .Y(alu_out[2]));
NOR_g _28788_ (.A(_14063_), .B(_07517_), .Y(_07527_));
NOR_g _28789_ (.A(_14064_), .B(_07527_), .Y(_07528_));
NAND_g _28790_ (.A(_08794_), .B(_07528_), .Y(_07529_));
NAND_g _28791_ (.A(instr_sub), .B(_14081_), .Y(_07530_));
AND_g _28792_ (.A(_07529_), .B(_07530_), .Y(_07531_));
XNOR_g _28793_ (.A(_14192_), .B(_07531_), .Y(_07532_));
NAND_g _28794_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07532_), .Y(_07533_));
NAND_g _28795_ (.A(_10743_), .B(_14191_), .Y(_07534_));
NOR_g _28796_ (.A(_14188_), .B(_07496_), .Y(_07535_));
NOR_g _28797_ (.A(_14190_), .B(_07497_), .Y(_07536_));
NOR_g _28798_ (.A(_07535_), .B(_07536_), .Y(_07537_));
AND_g _28799_ (.A(_07534_), .B(_07537_), .Y(_07538_));
NAND_g _28800_ (.A(_07533_), .B(_07538_), .Y(alu_out[3]));
NOR_g _28801_ (.A(_14188_), .B(_07528_), .Y(_07539_));
NOR_g _28802_ (.A(_14189_), .B(_07539_), .Y(_07540_));
NAND_g _28803_ (.A(_08794_), .B(_07540_), .Y(_07541_));
NAND_g _28804_ (.A(instr_sub), .B(_14085_), .Y(_07542_));
AND_g _28805_ (.A(_07541_), .B(_07542_), .Y(_07543_));
XNOR_g _28806_ (.A(_14061_), .B(_07543_), .Y(_07544_));
NAND_g _28807_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07544_), .Y(_07545_));
NAND_g _28808_ (.A(_10743_), .B(_14060_), .Y(_07546_));
NOR_g _28809_ (.A(_14057_), .B(_07496_), .Y(_07547_));
NOR_g _28810_ (.A(_14059_), .B(_07497_), .Y(_07548_));
NOR_g _28811_ (.A(_07547_), .B(_07548_), .Y(_07549_));
AND_g _28812_ (.A(_07546_), .B(_07549_), .Y(_07550_));
NAND_g _28813_ (.A(_07545_), .B(_07550_), .Y(alu_out[4]));
NOR_g _28814_ (.A(_14057_), .B(_07540_), .Y(_07551_));
NOR_g _28815_ (.A(_14058_), .B(_07551_), .Y(_07552_));
NAND_g _28816_ (.A(_08794_), .B(_07552_), .Y(_07553_));
NAND_g _28817_ (.A(instr_sub), .B(_14088_), .Y(_07554_));
NAND_g _28818_ (.A(_07553_), .B(_07554_), .Y(_07555_));
XOR_g _28819_ (.A(_14056_), .B(_07555_), .Y(_07556_));
NAND_g _28820_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07556_), .Y(_07557_));
NOR_g _28821_ (.A(_14055_), .B(_07497_), .Y(_07558_));
NAND_g _28822_ (.A(_10743_), .B(_14055_), .Y(_07559_));
AND_g _28823_ (.A(_07496_), .B(_07559_), .Y(_07560_));
NOR_g _28824_ (.A(_14053_), .B(_07560_), .Y(_07561_));
NOR_g _28825_ (.A(_07558_), .B(_07561_), .Y(_07562_));
NAND_g _28826_ (.A(_07557_), .B(_07562_), .Y(alu_out[5]));
NOR_g _28827_ (.A(_14053_), .B(_07552_), .Y(_07563_));
NOR_g _28828_ (.A(_14054_), .B(_07563_), .Y(_07564_));
NAND_g _28829_ (.A(_08794_), .B(_07564_), .Y(_07565_));
NAND_g _28830_ (.A(instr_sub), .B(_14090_), .Y(_07566_));
NAND_g _28831_ (.A(_07565_), .B(_07566_), .Y(_07567_));
XNOR_g _28832_ (.A(_14050_), .B(_07567_), .Y(_07568_));
NAND_g _28833_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07568_), .Y(_07569_));
NAND_g _28834_ (.A(_10743_), .B(_14050_), .Y(_07570_));
NOR_g _28835_ (.A(_14047_), .B(_07496_), .Y(_07571_));
NOR_g _28836_ (.A(_14049_), .B(_07497_), .Y(_07572_));
NOR_g _28837_ (.A(_07571_), .B(_07572_), .Y(_07573_));
AND_g _28838_ (.A(_07570_), .B(_07573_), .Y(_07574_));
NAND_g _28839_ (.A(_07569_), .B(_07574_), .Y(alu_out[6]));
NOR_g _28840_ (.A(_14047_), .B(_07564_), .Y(_07575_));
NOR_g _28841_ (.A(_14048_), .B(_07575_), .Y(_07576_));
NOR_g _28842_ (.A(instr_sub), .B(_07576_), .Y(_07577_));
AND_g _28843_ (.A(instr_sub), .B(_14092_), .Y(_07578_));
AND_g _28844_ (.A(_14091_), .B(_07578_), .Y(_07579_));
NOR_g _28845_ (.A(_07577_), .B(_07579_), .Y(_07580_));
XNOR_g _28846_ (.A(_14195_), .B(_07580_), .Y(_07581_));
NAND_g _28847_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07581_), .Y(_07582_));
NAND_g _28848_ (.A(_10743_), .B(_14195_), .Y(_07583_));
NOR_g _28849_ (.A(_14193_), .B(_07496_), .Y(_07584_));
NOR_g _28850_ (.A(_14194_), .B(_07497_), .Y(_07585_));
NOR_g _28851_ (.A(_07584_), .B(_07585_), .Y(_07586_));
AND_g _28852_ (.A(_07583_), .B(_07586_), .Y(_07587_));
NAND_g _28853_ (.A(_07582_), .B(_07587_), .Y(alu_out[7]));
AND_g _28854_ (.A(_14194_), .B(_07576_), .Y(_07588_));
NOR_g _28855_ (.A(_14193_), .B(_07588_), .Y(_07589_));
NOR_g _28856_ (.A(instr_sub), .B(_07589_), .Y(_07590_));
AND_g _28857_ (.A(instr_sub), .B(_14096_), .Y(_07591_));
NOR_g _28858_ (.A(_07590_), .B(_07591_), .Y(_07592_));
XNOR_g _28859_ (.A(_14023_), .B(_07592_), .Y(_07593_));
NAND_g _28860_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07593_), .Y(_07594_));
NAND_g _28861_ (.A(_10743_), .B(_14022_), .Y(_07595_));
NOR_g _28862_ (.A(_14021_), .B(_07497_), .Y(_07596_));
NOR_g _28863_ (.A(_14020_), .B(_07496_), .Y(_07597_));
NOR_g _28864_ (.A(_07596_), .B(_07597_), .Y(_07598_));
AND_g _28865_ (.A(_07595_), .B(_07598_), .Y(_07599_));
NAND_g _28866_ (.A(_07594_), .B(_07599_), .Y(alu_out[8]));
NAND_g _28867_ (.A(_14022_), .B(_07589_), .Y(_07600_));
AND_g _28868_ (.A(_14021_), .B(_07600_), .Y(_07601_));
NAND_g _28869_ (.A(_14023_), .B(_14096_), .Y(_07602_));
NAND_g _28870_ (.A(_14104_), .B(_07602_), .Y(_07603_));
NAND_g _28871_ (.A(instr_sub), .B(_07603_), .Y(_07604_));
NAND_g _28872_ (.A(_08794_), .B(_07601_), .Y(_07605_));
AND_g _28873_ (.A(_07604_), .B(_07605_), .Y(_07606_));
XNOR_g _28874_ (.A(_14019_), .B(_07606_), .Y(_07607_));
NAND_g _28875_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07607_), .Y(_07608_));
NAND_g _28876_ (.A(_10743_), .B(_14018_), .Y(_07609_));
NOR_g _28877_ (.A(_14016_), .B(_07496_), .Y(_07610_));
NOR_g _28878_ (.A(_14017_), .B(_07497_), .Y(_07611_));
NOR_g _28879_ (.A(_07610_), .B(_07611_), .Y(_07612_));
AND_g _28880_ (.A(_07609_), .B(_07612_), .Y(_07613_));
NAND_g _28881_ (.A(_07608_), .B(_07613_), .Y(alu_out[9]));
NAND_g _28882_ (.A(_14019_), .B(_07603_), .Y(_07614_));
NAND_g _28883_ (.A(_14103_), .B(_07614_), .Y(_07615_));
AND_g _28884_ (.A(_14017_), .B(_07601_), .Y(_07616_));
NOR_g _28885_ (.A(_14016_), .B(_07616_), .Y(_07617_));
NOR_g _28886_ (.A(instr_sub), .B(_07617_), .Y(_07618_));
AND_g _28887_ (.A(instr_sub), .B(_07615_), .Y(_07619_));
NOR_g _28888_ (.A(_07618_), .B(_07619_), .Y(_07620_));
XNOR_g _28889_ (.A(_14014_), .B(_07620_), .Y(_07621_));
NAND_g _28890_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07621_), .Y(_07622_));
NOR_g _28891_ (.A(_14013_), .B(_07497_), .Y(_07623_));
NAND_g _28892_ (.A(_10743_), .B(_14013_), .Y(_07624_));
AND_g _28893_ (.A(_07496_), .B(_07624_), .Y(_07625_));
NOR_g _28894_ (.A(_14011_), .B(_07625_), .Y(_07626_));
NOR_g _28895_ (.A(_07623_), .B(_07626_), .Y(_07627_));
NAND_g _28896_ (.A(_07622_), .B(_07627_), .Y(alu_out[10]));
NOR_g _28897_ (.A(_14012_), .B(_07617_), .Y(_07628_));
NOR_g _28898_ (.A(_14011_), .B(_07628_), .Y(_07629_));
NAND_g _28899_ (.A(_08794_), .B(_07629_), .Y(_07630_));
NAND_g _28900_ (.A(_14014_), .B(_07615_), .Y(_07631_));
NOR_g _28901_ (.A(_08794_), .B(_14109_), .Y(_07632_));
NAND_g _28902_ (.A(_07631_), .B(_07632_), .Y(_07633_));
AND_g _28903_ (.A(_07630_), .B(_07633_), .Y(_07634_));
XNOR_g _28904_ (.A(_14009_), .B(_07634_), .Y(_07635_));
NAND_g _28905_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07635_), .Y(_07636_));
NAND_g _28906_ (.A(_10743_), .B(_14009_), .Y(_07637_));
NOR_g _28907_ (.A(_14006_), .B(_07496_), .Y(_07638_));
NOR_g _28908_ (.A(_14008_), .B(_07497_), .Y(_07639_));
NOR_g _28909_ (.A(_07638_), .B(_07639_), .Y(_07640_));
AND_g _28910_ (.A(_07637_), .B(_07640_), .Y(_07641_));
NAND_g _28911_ (.A(_07636_), .B(_07641_), .Y(alu_out[11]));
NAND_g _28912_ (.A(_14025_), .B(_14096_), .Y(_07642_));
NAND_g _28913_ (.A(_14113_), .B(_07642_), .Y(_07643_));
NOR_g _28914_ (.A(_14007_), .B(_07629_), .Y(_07644_));
NOR_g _28915_ (.A(_14006_), .B(_07644_), .Y(_07645_));
NOR_g _28916_ (.A(instr_sub), .B(_07645_), .Y(_07646_));
AND_g _28917_ (.A(instr_sub), .B(_07643_), .Y(_07647_));
NOR_g _28918_ (.A(_07646_), .B(_07647_), .Y(_07648_));
XNOR_g _28919_ (.A(_14033_), .B(_07648_), .Y(_07649_));
NAND_g _28920_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07649_), .Y(_07650_));
NAND_g _28921_ (.A(_10743_), .B(_14032_), .Y(_07651_));
NOR_g _28922_ (.A(_14031_), .B(_07497_), .Y(_07652_));
NOR_g _28923_ (.A(_14030_), .B(_07496_), .Y(_07653_));
NOR_g _28924_ (.A(_07652_), .B(_07653_), .Y(_07654_));
AND_g _28925_ (.A(_07651_), .B(_07654_), .Y(_07655_));
NAND_g _28926_ (.A(_07650_), .B(_07655_), .Y(alu_out[12]));
AND_g _28927_ (.A(_14033_), .B(_07643_), .Y(_07656_));
NAND_g _28928_ (.A(_14033_), .B(_07643_), .Y(_07657_));
NAND_g _28929_ (.A(_14100_), .B(_07657_), .Y(_07658_));
NAND_g _28930_ (.A(instr_sub), .B(_07658_), .Y(_07659_));
NAND_g _28931_ (.A(_14032_), .B(_07645_), .Y(_07660_));
AND_g _28932_ (.A(_08794_), .B(_14031_), .Y(_07661_));
NAND_g _28933_ (.A(_07660_), .B(_07661_), .Y(_07662_));
AND_g _28934_ (.A(_07659_), .B(_07662_), .Y(_07663_));
XNOR_g _28935_ (.A(_14029_), .B(_07663_), .Y(_07664_));
NAND_g _28936_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07664_), .Y(_07665_));
NAND_g _28937_ (.A(_10743_), .B(_14028_), .Y(_07666_));
NOR_g _28938_ (.A(_14026_), .B(_07496_), .Y(_07667_));
NOR_g _28939_ (.A(_14027_), .B(_07497_), .Y(_07668_));
NOR_g _28940_ (.A(_07667_), .B(_07668_), .Y(_07669_));
AND_g _28941_ (.A(_07666_), .B(_07669_), .Y(_07670_));
NAND_g _28942_ (.A(_07665_), .B(_07670_), .Y(alu_out[13]));
NAND_g _28943_ (.A(_14029_), .B(_07656_), .Y(_07671_));
NAND_g _28944_ (.A(_14102_), .B(_07671_), .Y(_07672_));
AND_g _28945_ (.A(_14027_), .B(_14031_), .Y(_07673_));
AND_g _28946_ (.A(_07660_), .B(_07673_), .Y(_07674_));
NOR_g _28947_ (.A(_14026_), .B(_07674_), .Y(_07675_));
NOR_g _28948_ (.A(instr_sub), .B(_07675_), .Y(_07676_));
AND_g _28949_ (.A(instr_sub), .B(_07672_), .Y(_07677_));
NOR_g _28950_ (.A(_07676_), .B(_07677_), .Y(_07678_));
XNOR_g _28951_ (.A(_14042_), .B(_07678_), .Y(_07679_));
NAND_g _28952_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07679_), .Y(_07680_));
NAND_g _28953_ (.A(_10743_), .B(_14041_), .Y(_07681_));
NOR_g _28954_ (.A(_14040_), .B(_07497_), .Y(_07682_));
NOR_g _28955_ (.A(_14039_), .B(_07496_), .Y(_07683_));
NOR_g _28956_ (.A(_07682_), .B(_07683_), .Y(_07684_));
AND_g _28957_ (.A(_07681_), .B(_07684_), .Y(_07685_));
NAND_g _28958_ (.A(_07680_), .B(_07685_), .Y(alu_out[14]));
NAND_g _28959_ (.A(_14042_), .B(_07672_), .Y(_07686_));
NAND_g _28960_ (.A(_14120_), .B(_07686_), .Y(_07687_));
NAND_g _28961_ (.A(instr_sub), .B(_07687_), .Y(_07688_));
NAND_g _28962_ (.A(_14041_), .B(_07675_), .Y(_07689_));
AND_g _28963_ (.A(_08794_), .B(_14040_), .Y(_07690_));
NAND_g _28964_ (.A(_07689_), .B(_07690_), .Y(_07691_));
AND_g _28965_ (.A(_07688_), .B(_07691_), .Y(_07692_));
NAND_g _28966_ (.A(_07688_), .B(_07691_), .Y(_07693_));
NAND_g _28967_ (.A(_14037_), .B(_07692_), .Y(_07694_));
NAND_g _28968_ (.A(_14038_), .B(_07693_), .Y(_07695_));
AND_g _28969_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07695_), .Y(_07696_));
NAND_g _28970_ (.A(_07694_), .B(_07696_), .Y(_07697_));
NAND_g _28971_ (.A(_10743_), .B(_14037_), .Y(_07698_));
NOR_g _28972_ (.A(_14036_), .B(_07497_), .Y(_07699_));
NOR_g _28973_ (.A(_14035_), .B(_07496_), .Y(_07700_));
NOR_g _28974_ (.A(_07699_), .B(_07700_), .Y(_07701_));
AND_g _28975_ (.A(_07698_), .B(_07701_), .Y(_07702_));
NAND_g _28976_ (.A(_07697_), .B(_07702_), .Y(alu_out[15]));
AND_g _28977_ (.A(_14036_), .B(_14040_), .Y(_07703_));
AND_g _28978_ (.A(_07689_), .B(_07703_), .Y(_07704_));
NOR_g _28979_ (.A(_14035_), .B(_07704_), .Y(_07705_));
NOR_g _28980_ (.A(instr_sub), .B(_07705_), .Y(_07706_));
NOT_g _28981_ (.A(_07706_), .Y(_07707_));
NAND_g _28982_ (.A(instr_sub), .B(_14124_), .Y(_07708_));
NAND_g _28983_ (.A(_07707_), .B(_07708_), .Y(_07709_));
XNOR_g _28984_ (.A(_14128_), .B(_07709_), .Y(_07710_));
NAND_g _28985_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07710_), .Y(_07711_));
NAND_g _28986_ (.A(_10743_), .B(_14128_), .Y(_07712_));
NOR_g _28987_ (.A(_14127_), .B(_07497_), .Y(_07713_));
NOR_g _28988_ (.A(_14126_), .B(_07496_), .Y(_07714_));
NOR_g _28989_ (.A(_07713_), .B(_07714_), .Y(_07715_));
AND_g _28990_ (.A(_07712_), .B(_07715_), .Y(_07716_));
NAND_g _28991_ (.A(_07711_), .B(_07716_), .Y(alu_out[16]));
AND_g _28992_ (.A(instr_sub), .B(_13997_), .Y(_07717_));
NOR_g _28993_ (.A(_14128_), .B(_07708_), .Y(_07718_));
NOR_g _28994_ (.A(_07717_), .B(_07718_), .Y(_07719_));
NAND_g _28995_ (.A(_14128_), .B(_07705_), .Y(_07720_));
AND_g _28996_ (.A(_08794_), .B(_14127_), .Y(_07721_));
NAND_g _28997_ (.A(_07720_), .B(_07721_), .Y(_07722_));
AND_g _28998_ (.A(_07719_), .B(_07722_), .Y(_07723_));
XNOR_g _28999_ (.A(_13996_), .B(_07723_), .Y(_07724_));
NAND_g _29000_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07724_), .Y(_07725_));
NAND_g _29001_ (.A(_10743_), .B(_13995_), .Y(_07726_));
NOR_g _29002_ (.A(_13993_), .B(_07496_), .Y(_07727_));
NOR_g _29003_ (.A(_13994_), .B(_07497_), .Y(_07728_));
NOR_g _29004_ (.A(_07727_), .B(_07728_), .Y(_07729_));
AND_g _29005_ (.A(_07726_), .B(_07729_), .Y(_07730_));
NAND_g _29006_ (.A(_07725_), .B(_07730_), .Y(alu_out[17]));
AND_g _29007_ (.A(_13994_), .B(_14127_), .Y(_07731_));
AND_g _29008_ (.A(_07720_), .B(_07731_), .Y(_07732_));
NOR_g _29009_ (.A(_13993_), .B(_07732_), .Y(_07733_));
NOR_g _29010_ (.A(instr_sub), .B(_07733_), .Y(_07734_));
NAND_g _29011_ (.A(_13999_), .B(_14131_), .Y(_07735_));
AND_g _29012_ (.A(instr_sub), .B(_07735_), .Y(_07736_));
NOR_g _29013_ (.A(_07734_), .B(_07736_), .Y(_07737_));
XNOR_g _29014_ (.A(_13991_), .B(_07737_), .Y(_07738_));
NAND_g _29015_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07738_), .Y(_07739_));
NAND_g _29016_ (.A(_10743_), .B(_13990_), .Y(_07740_));
NOR_g _29017_ (.A(_13989_), .B(_07497_), .Y(_07741_));
NOR_g _29018_ (.A(_13987_), .B(_07496_), .Y(_07742_));
NOR_g _29019_ (.A(_07741_), .B(_07742_), .Y(_07743_));
AND_g _29020_ (.A(_07740_), .B(_07743_), .Y(_07744_));
NAND_g _29021_ (.A(_07739_), .B(_07744_), .Y(alu_out[18]));
NAND_g _29022_ (.A(_13991_), .B(_07735_), .Y(_07745_));
NAND_g _29023_ (.A(_13986_), .B(_07745_), .Y(_07746_));
NAND_g _29024_ (.A(instr_sub), .B(_07746_), .Y(_07747_));
NAND_g _29025_ (.A(_13988_), .B(_07733_), .Y(_07748_));
AND_g _29026_ (.A(_08794_), .B(_13989_), .Y(_07749_));
NAND_g _29027_ (.A(_07748_), .B(_07749_), .Y(_07750_));
AND_g _29028_ (.A(_07747_), .B(_07750_), .Y(_07751_));
XNOR_g _29029_ (.A(_13985_), .B(_07751_), .Y(_07752_));
NAND_g _29030_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07752_), .Y(_07753_));
NAND_g _29031_ (.A(_10743_), .B(_13984_), .Y(_07754_));
NOR_g _29032_ (.A(_13981_), .B(_07496_), .Y(_07755_));
NOR_g _29033_ (.A(_13983_), .B(_07497_), .Y(_07756_));
NOR_g _29034_ (.A(_07755_), .B(_07756_), .Y(_07757_));
AND_g _29035_ (.A(_07754_), .B(_07757_), .Y(_07758_));
NAND_g _29036_ (.A(_07753_), .B(_07758_), .Y(alu_out[19]));
NAND_g _29037_ (.A(instr_sub), .B(_14133_), .Y(_07759_));
AND_g _29038_ (.A(_13983_), .B(_13989_), .Y(_07760_));
NAND_g _29039_ (.A(_07748_), .B(_07760_), .Y(_07761_));
NAND_g _29040_ (.A(_13982_), .B(_07761_), .Y(_07762_));
NAND_g _29041_ (.A(_08794_), .B(_07762_), .Y(_07763_));
AND_g _29042_ (.A(_07759_), .B(_07763_), .Y(_07764_));
NAND_g _29043_ (.A(_07759_), .B(_07763_), .Y(_07765_));
NAND_g _29044_ (.A(_14136_), .B(_07764_), .Y(_07766_));
NAND_g _29045_ (.A(_14137_), .B(_07765_), .Y(_07767_));
AND_g _29046_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07767_), .Y(_07768_));
NAND_g _29047_ (.A(_07766_), .B(_07768_), .Y(_07769_));
NAND_g _29048_ (.A(_10743_), .B(_14136_), .Y(_07770_));
NOR_g _29049_ (.A(_14135_), .B(_07497_), .Y(_07771_));
NOR_g _29050_ (.A(_14134_), .B(_07496_), .Y(_07772_));
NOR_g _29051_ (.A(_07771_), .B(_07772_), .Y(_07773_));
AND_g _29052_ (.A(_07770_), .B(_07773_), .Y(_07774_));
NAND_g _29053_ (.A(_07769_), .B(_07774_), .Y(alu_out[20]));
AND_g _29054_ (.A(_14135_), .B(_07762_), .Y(_07775_));
NOR_g _29055_ (.A(_14134_), .B(_07775_), .Y(_07776_));
AND_g _29056_ (.A(_08794_), .B(_07776_), .Y(_07777_));
NAND_g _29057_ (.A(instr_sub), .B(_13969_), .Y(_07778_));
NOR_g _29058_ (.A(_14138_), .B(_07778_), .Y(_07779_));
NOR_g _29059_ (.A(_07777_), .B(_07779_), .Y(_07780_));
XNOR_g _29060_ (.A(_13966_), .B(_07780_), .Y(_07781_));
NAND_g _29061_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07781_), .Y(_07782_));
NAND_g _29062_ (.A(_10743_), .B(_13966_), .Y(_07783_));
NOR_g _29063_ (.A(_13963_), .B(_07496_), .Y(_07784_));
NOR_g _29064_ (.A(_13965_), .B(_07497_), .Y(_07785_));
NOR_g _29065_ (.A(_07784_), .B(_07785_), .Y(_07786_));
AND_g _29066_ (.A(_07783_), .B(_07786_), .Y(_07787_));
NAND_g _29067_ (.A(_07782_), .B(_07787_), .Y(alu_out[21]));
NAND_g _29068_ (.A(_13964_), .B(_07776_), .Y(_07788_));
NAND_g _29069_ (.A(_13965_), .B(_07788_), .Y(_07789_));
AND_g _29070_ (.A(_13965_), .B(_07788_), .Y(_07790_));
NAND_g _29071_ (.A(_08794_), .B(_07790_), .Y(_07791_));
NAND_g _29072_ (.A(_13971_), .B(_14139_), .Y(_07792_));
NAND_g _29073_ (.A(instr_sub), .B(_07792_), .Y(_07793_));
AND_g _29074_ (.A(_07791_), .B(_07793_), .Y(_07794_));
NAND_g _29075_ (.A(_07791_), .B(_07793_), .Y(_07795_));
NAND_g _29076_ (.A(_13959_), .B(_07794_), .Y(_07796_));
NAND_g _29077_ (.A(_13960_), .B(_07795_), .Y(_07797_));
AND_g _29078_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07797_), .Y(_07798_));
NAND_g _29079_ (.A(_07796_), .B(_07798_), .Y(_07799_));
NAND_g _29080_ (.A(_10743_), .B(_13959_), .Y(_07800_));
NOR_g _29081_ (.A(_13958_), .B(_07497_), .Y(_07801_));
NOR_g _29082_ (.A(_13956_), .B(_07496_), .Y(_07802_));
NOR_g _29083_ (.A(_07801_), .B(_07802_), .Y(_07803_));
AND_g _29084_ (.A(_07800_), .B(_07803_), .Y(_07804_));
NAND_g _29085_ (.A(_07799_), .B(_07804_), .Y(alu_out[22]));
NAND_g _29086_ (.A(_13960_), .B(_07792_), .Y(_07805_));
NAND_g _29087_ (.A(_13975_), .B(_07805_), .Y(_07806_));
NAND_g _29088_ (.A(instr_sub), .B(_07806_), .Y(_07807_));
NAND_g _29089_ (.A(_13957_), .B(_07789_), .Y(_07808_));
AND_g _29090_ (.A(_08794_), .B(_13958_), .Y(_07809_));
NAND_g _29091_ (.A(_07808_), .B(_07809_), .Y(_07810_));
AND_g _29092_ (.A(_07807_), .B(_07810_), .Y(_07811_));
NAND_g _29093_ (.A(_07807_), .B(_07810_), .Y(_07812_));
NAND_g _29094_ (.A(_13954_), .B(_07811_), .Y(_07813_));
NAND_g _29095_ (.A(_13955_), .B(_07812_), .Y(_07814_));
AND_g _29096_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07814_), .Y(_07815_));
NAND_g _29097_ (.A(_07813_), .B(_07815_), .Y(_07816_));
NAND_g _29098_ (.A(_10743_), .B(_13954_), .Y(_07817_));
NOR_g _29099_ (.A(_13953_), .B(_07497_), .Y(_07818_));
NOR_g _29100_ (.A(_13952_), .B(_07496_), .Y(_07819_));
NOR_g _29101_ (.A(_07818_), .B(_07819_), .Y(_07820_));
AND_g _29102_ (.A(_07817_), .B(_07820_), .Y(_07821_));
NAND_g _29103_ (.A(_07816_), .B(_07821_), .Y(alu_out[23]));
AND_g _29104_ (.A(_13953_), .B(_13958_), .Y(_07822_));
AND_g _29105_ (.A(_07808_), .B(_07822_), .Y(_07823_));
NOR_g _29106_ (.A(_13952_), .B(_07823_), .Y(_07824_));
NOR_g _29107_ (.A(instr_sub), .B(_07824_), .Y(_07825_));
AND_g _29108_ (.A(instr_sub), .B(_14143_), .Y(_07826_));
NOR_g _29109_ (.A(_07825_), .B(_07826_), .Y(_07827_));
XNOR_g _29110_ (.A(_14147_), .B(_07827_), .Y(_07828_));
NAND_g _29111_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07828_), .Y(_07829_));
NAND_g _29112_ (.A(_10743_), .B(_14146_), .Y(_07830_));
NOR_g _29113_ (.A(_14145_), .B(_07497_), .Y(_07831_));
NOR_g _29114_ (.A(_14144_), .B(_07496_), .Y(_07832_));
NOR_g _29115_ (.A(_07831_), .B(_07832_), .Y(_07833_));
AND_g _29116_ (.A(_07830_), .B(_07833_), .Y(_07834_));
NAND_g _29117_ (.A(_07829_), .B(_07834_), .Y(alu_out[24]));
NAND_g _29118_ (.A(_14146_), .B(_07824_), .Y(_07835_));
AND_g _29119_ (.A(_08794_), .B(_14145_), .Y(_07836_));
NAND_g _29120_ (.A(_07835_), .B(_07836_), .Y(_07837_));
NAND_g _29121_ (.A(instr_sub), .B(_13940_), .Y(_07838_));
NAND_g _29122_ (.A(_14147_), .B(_07826_), .Y(_07839_));
AND_g _29123_ (.A(_07838_), .B(_07839_), .Y(_07840_));
AND_g _29124_ (.A(_07837_), .B(_07840_), .Y(_07841_));
NAND_g _29125_ (.A(_07837_), .B(_07840_), .Y(_07842_));
NAND_g _29126_ (.A(_13938_), .B(_07841_), .Y(_07843_));
NAND_g _29127_ (.A(_13939_), .B(_07842_), .Y(_07844_));
AND_g _29128_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07844_), .Y(_07845_));
NAND_g _29129_ (.A(_07843_), .B(_07845_), .Y(_07846_));
NAND_g _29130_ (.A(_10743_), .B(_13938_), .Y(_07847_));
NOR_g _29131_ (.A(_13937_), .B(_07497_), .Y(_07848_));
NOR_g _29132_ (.A(_13936_), .B(_07496_), .Y(_07849_));
NOR_g _29133_ (.A(_07848_), .B(_07849_), .Y(_07850_));
AND_g _29134_ (.A(_07847_), .B(_07850_), .Y(_07851_));
NAND_g _29135_ (.A(_07846_), .B(_07851_), .Y(alu_out[25]));
AND_g _29136_ (.A(_13937_), .B(_14145_), .Y(_07852_));
AND_g _29137_ (.A(_07835_), .B(_07852_), .Y(_07853_));
NOR_g _29138_ (.A(_13936_), .B(_07853_), .Y(_07854_));
NOR_g _29139_ (.A(instr_sub), .B(_07854_), .Y(_07855_));
NAND_g _29140_ (.A(_13942_), .B(_14150_), .Y(_07856_));
AND_g _29141_ (.A(instr_sub), .B(_07856_), .Y(_07857_));
NOR_g _29142_ (.A(_07855_), .B(_07857_), .Y(_07858_));
XNOR_g _29143_ (.A(_13933_), .B(_07858_), .Y(_07859_));
NAND_g _29144_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07859_), .Y(_07860_));
NAND_g _29145_ (.A(_10743_), .B(_13932_), .Y(_07861_));
NOR_g _29146_ (.A(_13931_), .B(_07497_), .Y(_07862_));
NOR_g _29147_ (.A(_13930_), .B(_07496_), .Y(_07863_));
NOR_g _29148_ (.A(_07862_), .B(_07863_), .Y(_07864_));
AND_g _29149_ (.A(_07861_), .B(_07864_), .Y(_07865_));
NAND_g _29150_ (.A(_07860_), .B(_07865_), .Y(alu_out[26]));
NAND_g _29151_ (.A(_13933_), .B(_07856_), .Y(_07866_));
NAND_g _29152_ (.A(_13946_), .B(_07866_), .Y(_07867_));
NAND_g _29153_ (.A(instr_sub), .B(_07867_), .Y(_07868_));
NAND_g _29154_ (.A(_13932_), .B(_07854_), .Y(_07869_));
AND_g _29155_ (.A(_08794_), .B(_13931_), .Y(_07870_));
NAND_g _29156_ (.A(_07869_), .B(_07870_), .Y(_07871_));
AND_g _29157_ (.A(_07868_), .B(_07871_), .Y(_07872_));
XNOR_g _29158_ (.A(_13929_), .B(_07872_), .Y(_07873_));
NAND_g _29159_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07873_), .Y(_07874_));
NAND_g _29160_ (.A(_10743_), .B(_13928_), .Y(_07875_));
NOR_g _29161_ (.A(_13925_), .B(_07496_), .Y(_07876_));
NOR_g _29162_ (.A(_13927_), .B(_07497_), .Y(_07877_));
NOR_g _29163_ (.A(_07876_), .B(_07877_), .Y(_07878_));
AND_g _29164_ (.A(_07875_), .B(_07878_), .Y(_07879_));
NAND_g _29165_ (.A(_07874_), .B(_07879_), .Y(alu_out[27]));
AND_g _29166_ (.A(_13927_), .B(_13931_), .Y(_07880_));
NAND_g _29167_ (.A(_07869_), .B(_07880_), .Y(_07881_));
NAND_g _29168_ (.A(_13926_), .B(_07881_), .Y(_07882_));
NAND_g _29169_ (.A(_08794_), .B(_07882_), .Y(_07883_));
NAND_g _29170_ (.A(instr_sub), .B(_14152_), .Y(_07884_));
AND_g _29171_ (.A(_07883_), .B(_07884_), .Y(_07885_));
XNOR_g _29172_ (.A(_13924_), .B(_07885_), .Y(_07886_));
NAND_g _29173_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07886_), .Y(_07887_));
NAND_g _29174_ (.A(_10743_), .B(_13923_), .Y(_07888_));
NOR_g _29175_ (.A(_13921_), .B(_07496_), .Y(_07889_));
NOR_g _29176_ (.A(_13922_), .B(_07497_), .Y(_07890_));
NOR_g _29177_ (.A(_07889_), .B(_07890_), .Y(_07891_));
AND_g _29178_ (.A(_07888_), .B(_07891_), .Y(_07892_));
NAND_g _29179_ (.A(_07887_), .B(_07892_), .Y(alu_out[28]));
AND_g _29180_ (.A(_13922_), .B(_07882_), .Y(_07893_));
NOR_g _29181_ (.A(_13921_), .B(_07893_), .Y(_07894_));
NAND_g _29182_ (.A(_08794_), .B(_07894_), .Y(_07895_));
NOR_g _29183_ (.A(_08794_), .B(_13917_), .Y(_07896_));
NAND_g _29184_ (.A(_14154_), .B(_07896_), .Y(_07897_));
AND_g _29185_ (.A(_07895_), .B(_07897_), .Y(_07898_));
NAND_g _29186_ (.A(_13916_), .B(_07898_), .Y(_07899_));
NOR_g _29187_ (.A(_13916_), .B(_07898_), .Y(_07900_));
NOR_g _29188_ (.A(_09023_), .B(_07900_), .Y(_07901_));
NAND_g _29189_ (.A(_07899_), .B(_07901_), .Y(_07902_));
NAND_g _29190_ (.A(_10743_), .B(_13915_), .Y(_07903_));
NOR_g _29191_ (.A(_13914_), .B(_07497_), .Y(_07904_));
NOR_g _29192_ (.A(_13912_), .B(_07496_), .Y(_07905_));
NOR_g _29193_ (.A(_07904_), .B(_07905_), .Y(_07906_));
AND_g _29194_ (.A(_07903_), .B(_07906_), .Y(_07907_));
NAND_g _29195_ (.A(_07902_), .B(_07907_), .Y(alu_out[29]));
NAND_g _29196_ (.A(_13913_), .B(_07894_), .Y(_07908_));
AND_g _29197_ (.A(_13914_), .B(_07908_), .Y(_07909_));
NAND_g _29198_ (.A(_13914_), .B(_07908_), .Y(_07910_));
NAND_g _29199_ (.A(_08794_), .B(_07909_), .Y(_07911_));
NAND_g _29200_ (.A(instr_sub), .B(_14156_), .Y(_07912_));
AND_g _29201_ (.A(_07911_), .B(_07912_), .Y(_07913_));
NAND_g _29202_ (.A(_07911_), .B(_07912_), .Y(_07914_));
NAND_g _29203_ (.A(_13909_), .B(_07913_), .Y(_07915_));
NAND_g _29204_ (.A(_13910_), .B(_07914_), .Y(_07916_));
AND_g _29205_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07916_), .Y(_07917_));
NAND_g _29206_ (.A(_07915_), .B(_07917_), .Y(_07918_));
NAND_g _29207_ (.A(_10743_), .B(_13909_), .Y(_07919_));
NOR_g _29208_ (.A(_13908_), .B(_07497_), .Y(_07920_));
NOR_g _29209_ (.A(_13907_), .B(_07496_), .Y(_07921_));
NOR_g _29210_ (.A(_07920_), .B(_07921_), .Y(_07922_));
AND_g _29211_ (.A(_07919_), .B(_07922_), .Y(_07923_));
NAND_g _29212_ (.A(_07918_), .B(_07923_), .Y(alu_out[30]));
NAND_g _29213_ (.A(instr_sub), .B(_14159_), .Y(_07924_));
NAND_g _29214_ (.A(_13909_), .B(_07910_), .Y(_07925_));
AND_g _29215_ (.A(_08794_), .B(_13908_), .Y(_07926_));
NAND_g _29216_ (.A(_07925_), .B(_07926_), .Y(_07927_));
AND_g _29217_ (.A(_07924_), .B(_07927_), .Y(_07928_));
XNOR_g _29218_ (.A(_13904_), .B(_07928_), .Y(_07929_));
NAND_g _29219_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_07929_), .Y(_07930_));
NAND_g _29220_ (.A(_10743_), .B(_13903_), .Y(_07931_));
NOR_g _29221_ (.A(_13901_), .B(_07496_), .Y(_07932_));
NOR_g _29222_ (.A(_13902_), .B(_07497_), .Y(_07933_));
NOR_g _29223_ (.A(_07932_), .B(_07933_), .Y(_07934_));
AND_g _29224_ (.A(_07931_), .B(_07934_), .Y(_07935_));
NAND_g _29225_ (.A(_07930_), .B(_07935_), .Y(alu_out[31]));
NAND_g _29226_ (.A(_14212_), .B(_14221_), .Y(_07936_));
NAND_g _29227_ (.A(_14393_), .B(_07936_), .Y(_07937_));
NAND_g _29228_ (.A(_13861_), .B(_07937_), .Y(_00000_));
NAND_g _29229_ (.A(_08799_), .B(_08800_), .Y(_07938_));
NOR_g _29230_ (.A(latched_is_lb), .B(_07938_), .Y(_07939_));
NOT_g _29231_ (.A(_07939_), .Y(_07940_));
AND_g _29232_ (.A(_13849_), .B(_13854_), .Y(_07941_));
AND_g _29233_ (.A(_07940_), .B(_07941_), .Y(_07942_));
NAND_g _29234_ (.A(mem_rdata[16]), .B(_01791_), .Y(_07943_));
NAND_g _29235_ (.A(mem_rdata[0]), .B(mem_la_wstrb[0]), .Y(_07944_));
NOR_g _29236_ (.A(_08843_), .B(_01784_), .Y(_07945_));
NAND_g _29237_ (.A(mem_rdata[8]), .B(_07945_), .Y(_07946_));
NAND_g _29238_ (.A(mem_rdata[24]), .B(_01796_), .Y(_07947_));
AND_g _29239_ (.A(_07946_), .B(_07947_), .Y(_07948_));
AND_g _29240_ (.A(_07944_), .B(_07948_), .Y(_07949_));
NAND_g _29241_ (.A(_07943_), .B(_07949_), .Y(_07950_));
NAND_g _29242_ (.A(_07942_), .B(_07950_), .Y(_07951_));
NAND_g _29243_ (.A(pcpi_rs1[0]), .B(_13889_), .Y(_07952_));
NAND_g _29244_ (.A(count_instr[0]), .B(instr_rdinstr), .Y(_07953_));
NAND_g _29245_ (.A(instr_rdcycleh), .B(count_cycle[32]), .Y(_07954_));
AND_g _29246_ (.A(_07953_), .B(_07954_), .Y(_07955_));
NAND_g _29247_ (.A(instr_rdcycle), .B(count_cycle[0]), .Y(_07956_));
NAND_g _29248_ (.A(count_instr[32]), .B(instr_rdinstrh), .Y(_07957_));
AND_g _29249_ (.A(_07956_), .B(_07957_), .Y(_07958_));
NAND_g _29250_ (.A(_07955_), .B(_07958_), .Y(_07959_));
NAND_g _29251_ (.A(_10595_), .B(_07959_), .Y(_07960_));
AND_g _29252_ (.A(reg_next_pc[0]), .B(decoded_imm[0]), .Y(_07961_));
XOR_g _29253_ (.A(reg_next_pc[0]), .B(decoded_imm[0]), .Y(_07962_));
NAND_g _29254_ (.A(_14214_), .B(_07962_), .Y(_07963_));
AND_g _29255_ (.A(_07960_), .B(_07963_), .Y(_07964_));
AND_g _29256_ (.A(_07952_), .B(_07964_), .Y(_07965_));
NAND_g _29257_ (.A(_07951_), .B(_07965_), .Y(_07966_));
AND_g _29258_ (.A(resetn), .B(_07966_), .Y(_00005_[0]));
NAND_g _29259_ (.A(mem_rdata[17]), .B(_01791_), .Y(_07967_));
NAND_g _29260_ (.A(mem_rdata[9]), .B(_07945_), .Y(_07968_));
NAND_g _29261_ (.A(mem_rdata[1]), .B(mem_la_wstrb[0]), .Y(_07969_));
NAND_g _29262_ (.A(mem_rdata[25]), .B(_01796_), .Y(_07970_));
AND_g _29263_ (.A(_07969_), .B(_07970_), .Y(_07971_));
AND_g _29264_ (.A(_07968_), .B(_07971_), .Y(_07972_));
NAND_g _29265_ (.A(_07967_), .B(_07972_), .Y(_07973_));
NAND_g _29266_ (.A(_07942_), .B(_07973_), .Y(_07974_));
NAND_g _29267_ (.A(pcpi_rs1[1]), .B(_13889_), .Y(_07975_));
NAND_g _29268_ (.A(count_instr[33]), .B(instr_rdinstrh), .Y(_07976_));
NAND_g _29269_ (.A(instr_rdcycle), .B(count_cycle[1]), .Y(_07977_));
NAND_g _29270_ (.A(instr_rdcycleh), .B(count_cycle[33]), .Y(_07978_));
NAND_g _29271_ (.A(count_instr[1]), .B(instr_rdinstr), .Y(_07979_));
AND_g _29272_ (.A(_07977_), .B(_07979_), .Y(_07980_));
AND_g _29273_ (.A(_07976_), .B(_07978_), .Y(_07981_));
NAND_g _29274_ (.A(_07980_), .B(_07981_), .Y(_07982_));
NAND_g _29275_ (.A(_10595_), .B(_07982_), .Y(_07983_));
NAND_g _29276_ (.A(reg_pc[1]), .B(decoded_imm[1]), .Y(_07984_));
XOR_g _29277_ (.A(reg_pc[1]), .B(decoded_imm[1]), .Y(_07985_));
NAND_g _29278_ (.A(_07961_), .B(_07985_), .Y(_07986_));
XOR_g _29279_ (.A(_07961_), .B(_07985_), .Y(_07987_));
NAND_g _29280_ (.A(_14214_), .B(_07987_), .Y(_07988_));
AND_g _29281_ (.A(_07983_), .B(_07988_), .Y(_07989_));
AND_g _29282_ (.A(_07975_), .B(_07989_), .Y(_07990_));
NAND_g _29283_ (.A(_07974_), .B(_07990_), .Y(_07991_));
AND_g _29284_ (.A(resetn), .B(_07991_), .Y(_00005_[1]));
NAND_g _29285_ (.A(mem_rdata[18]), .B(_01791_), .Y(_07992_));
NAND_g _29286_ (.A(mem_rdata[10]), .B(_07945_), .Y(_07993_));
NAND_g _29287_ (.A(mem_rdata[2]), .B(mem_la_wstrb[0]), .Y(_07994_));
NAND_g _29288_ (.A(mem_rdata[26]), .B(_01796_), .Y(_07995_));
AND_g _29289_ (.A(_07994_), .B(_07995_), .Y(_07996_));
AND_g _29290_ (.A(_07993_), .B(_07996_), .Y(_07997_));
NAND_g _29291_ (.A(_07992_), .B(_07997_), .Y(_07998_));
NAND_g _29292_ (.A(_07942_), .B(_07998_), .Y(_07999_));
NAND_g _29293_ (.A(pcpi_rs1[2]), .B(_13889_), .Y(_08000_));
NAND_g _29294_ (.A(count_instr[2]), .B(instr_rdinstr), .Y(_08001_));
NAND_g _29295_ (.A(instr_rdcycleh), .B(count_cycle[34]), .Y(_08002_));
NAND_g _29296_ (.A(instr_rdcycle), .B(count_cycle[2]), .Y(_08003_));
NAND_g _29297_ (.A(count_instr[34]), .B(instr_rdinstrh), .Y(_08004_));
AND_g _29298_ (.A(_08002_), .B(_08004_), .Y(_08005_));
AND_g _29299_ (.A(_08001_), .B(_08003_), .Y(_08006_));
NAND_g _29300_ (.A(_08005_), .B(_08006_), .Y(_08007_));
NAND_g _29301_ (.A(_10595_), .B(_08007_), .Y(_08008_));
AND_g _29302_ (.A(_08000_), .B(_08008_), .Y(_08009_));
NAND_g _29303_ (.A(_07984_), .B(_07986_), .Y(_08010_));
NAND_g _29304_ (.A(reg_pc[2]), .B(decoded_imm[2]), .Y(_08011_));
XOR_g _29305_ (.A(reg_pc[2]), .B(decoded_imm[2]), .Y(_08012_));
NAND_g _29306_ (.A(_08010_), .B(_08012_), .Y(_08013_));
AND_g _29307_ (.A(_07999_), .B(_08009_), .Y(_08014_));
XOR_g _29308_ (.A(_08010_), .B(_08012_), .Y(_08015_));
NAND_g _29309_ (.A(_14217_), .B(_08015_), .Y(_08016_));
NAND_g _29310_ (.A(_08014_), .B(_08016_), .Y(_08017_));
AND_g _29311_ (.A(resetn), .B(_08017_), .Y(_00005_[2]));
AND_g _29312_ (.A(_08011_), .B(_08013_), .Y(_08018_));
NAND_g _29313_ (.A(_08011_), .B(_08013_), .Y(_08019_));
NAND_g _29314_ (.A(reg_pc[3]), .B(decoded_imm[3]), .Y(_08020_));
XOR_g _29315_ (.A(reg_pc[3]), .B(decoded_imm[3]), .Y(_08021_));
XNOR_g _29316_ (.A(reg_pc[3]), .B(decoded_imm[3]), .Y(_08022_));
NAND_g _29317_ (.A(_08018_), .B(_08022_), .Y(_08023_));
NAND_g _29318_ (.A(_08019_), .B(_08021_), .Y(_08024_));
NAND_g _29319_ (.A(mem_rdata[19]), .B(_01791_), .Y(_08025_));
NAND_g _29320_ (.A(mem_rdata[11]), .B(_07945_), .Y(_08026_));
NAND_g _29321_ (.A(mem_rdata[3]), .B(mem_la_wstrb[0]), .Y(_08027_));
NAND_g _29322_ (.A(mem_rdata[27]), .B(_01796_), .Y(_08028_));
AND_g _29323_ (.A(_08027_), .B(_08028_), .Y(_08029_));
AND_g _29324_ (.A(_08026_), .B(_08029_), .Y(_08030_));
NAND_g _29325_ (.A(_08025_), .B(_08030_), .Y(_08031_));
NAND_g _29326_ (.A(_07942_), .B(_08031_), .Y(_08032_));
NAND_g _29327_ (.A(pcpi_rs1[3]), .B(_13889_), .Y(_08033_));
NAND_g _29328_ (.A(instr_rdcycleh), .B(count_cycle[35]), .Y(_08034_));
NAND_g _29329_ (.A(count_instr[35]), .B(instr_rdinstrh), .Y(_08035_));
AND_g _29330_ (.A(_08034_), .B(_08035_), .Y(_08036_));
NAND_g _29331_ (.A(count_instr[3]), .B(instr_rdinstr), .Y(_08037_));
NAND_g _29332_ (.A(instr_rdcycle), .B(count_cycle[3]), .Y(_08038_));
AND_g _29333_ (.A(_08037_), .B(_08038_), .Y(_08039_));
NAND_g _29334_ (.A(_08036_), .B(_08039_), .Y(_08040_));
NAND_g _29335_ (.A(_10595_), .B(_08040_), .Y(_08041_));
AND_g _29336_ (.A(_08033_), .B(_08041_), .Y(_08042_));
AND_g _29337_ (.A(_14217_), .B(_08023_), .Y(_08043_));
NAND_g _29338_ (.A(_08024_), .B(_08043_), .Y(_08044_));
AND_g _29339_ (.A(_08042_), .B(_08044_), .Y(_08045_));
NAND_g _29340_ (.A(_08032_), .B(_08045_), .Y(_08046_));
AND_g _29341_ (.A(resetn), .B(_08046_), .Y(_00005_[3]));
NAND_g _29342_ (.A(mem_rdata[20]), .B(_01791_), .Y(_08047_));
NAND_g _29343_ (.A(mem_rdata[4]), .B(mem_la_wstrb[0]), .Y(_08048_));
NAND_g _29344_ (.A(mem_rdata[12]), .B(_07945_), .Y(_08049_));
NAND_g _29345_ (.A(mem_rdata[28]), .B(_01796_), .Y(_08050_));
AND_g _29346_ (.A(_08049_), .B(_08050_), .Y(_08051_));
AND_g _29347_ (.A(_08048_), .B(_08051_), .Y(_08052_));
NAND_g _29348_ (.A(_08047_), .B(_08052_), .Y(_08053_));
NAND_g _29349_ (.A(_07942_), .B(_08053_), .Y(_08054_));
NAND_g _29350_ (.A(count_instr[4]), .B(instr_rdinstr), .Y(_08055_));
NAND_g _29351_ (.A(instr_rdcycleh), .B(count_cycle[36]), .Y(_08056_));
AND_g _29352_ (.A(_08055_), .B(_08056_), .Y(_08057_));
NAND_g _29353_ (.A(count_instr[36]), .B(instr_rdinstrh), .Y(_08058_));
NAND_g _29354_ (.A(instr_rdcycle), .B(count_cycle[4]), .Y(_08059_));
AND_g _29355_ (.A(_08058_), .B(_08059_), .Y(_08060_));
NAND_g _29356_ (.A(_08057_), .B(_08060_), .Y(_08061_));
NAND_g _29357_ (.A(_10595_), .B(_08061_), .Y(_08062_));
NAND_g _29358_ (.A(pcpi_rs1[4]), .B(_13889_), .Y(_08063_));
AND_g _29359_ (.A(_08062_), .B(_08063_), .Y(_08064_));
AND_g _29360_ (.A(_08054_), .B(_08064_), .Y(_08065_));
NAND_g _29361_ (.A(_08020_), .B(_08024_), .Y(_08066_));
NAND_g _29362_ (.A(reg_pc[4]), .B(decoded_imm[4]), .Y(_08067_));
XOR_g _29363_ (.A(reg_pc[4]), .B(decoded_imm[4]), .Y(_08068_));
NAND_g _29364_ (.A(_08066_), .B(_08068_), .Y(_08069_));
XOR_g _29365_ (.A(_08066_), .B(_08068_), .Y(_08070_));
NAND_g _29366_ (.A(_14217_), .B(_08070_), .Y(_08071_));
NAND_g _29367_ (.A(_08065_), .B(_08071_), .Y(_08072_));
AND_g _29368_ (.A(resetn), .B(_08072_), .Y(_00005_[4]));
NAND_g _29369_ (.A(mem_rdata[21]), .B(_01791_), .Y(_08073_));
NAND_g _29370_ (.A(mem_rdata[13]), .B(_07945_), .Y(_08074_));
NAND_g _29371_ (.A(mem_rdata[5]), .B(mem_la_wstrb[0]), .Y(_08075_));
NAND_g _29372_ (.A(mem_rdata[29]), .B(_01796_), .Y(_08076_));
AND_g _29373_ (.A(_08075_), .B(_08076_), .Y(_08077_));
AND_g _29374_ (.A(_08074_), .B(_08077_), .Y(_08078_));
NAND_g _29375_ (.A(_08073_), .B(_08078_), .Y(_08079_));
NAND_g _29376_ (.A(_07942_), .B(_08079_), .Y(_08080_));
NAND_g _29377_ (.A(instr_rdcycleh), .B(count_cycle[37]), .Y(_08081_));
NAND_g _29378_ (.A(count_instr[37]), .B(instr_rdinstrh), .Y(_08082_));
AND_g _29379_ (.A(_08081_), .B(_08082_), .Y(_08083_));
NAND_g _29380_ (.A(count_instr[5]), .B(instr_rdinstr), .Y(_08084_));
NAND_g _29381_ (.A(instr_rdcycle), .B(count_cycle[5]), .Y(_08085_));
AND_g _29382_ (.A(_08084_), .B(_08085_), .Y(_08086_));
NAND_g _29383_ (.A(_08083_), .B(_08086_), .Y(_08087_));
NAND_g _29384_ (.A(_10595_), .B(_08087_), .Y(_08088_));
NAND_g _29385_ (.A(pcpi_rs1[5]), .B(_13889_), .Y(_08089_));
AND_g _29386_ (.A(_08088_), .B(_08089_), .Y(_08090_));
AND_g _29387_ (.A(_08080_), .B(_08090_), .Y(_08091_));
NAND_g _29388_ (.A(_08067_), .B(_08069_), .Y(_08092_));
NAND_g _29389_ (.A(reg_pc[5]), .B(decoded_imm[5]), .Y(_08093_));
XOR_g _29390_ (.A(reg_pc[5]), .B(decoded_imm[5]), .Y(_08094_));
NAND_g _29391_ (.A(_08092_), .B(_08094_), .Y(_08095_));
XOR_g _29392_ (.A(_08092_), .B(_08094_), .Y(_08096_));
NAND_g _29393_ (.A(_14217_), .B(_08096_), .Y(_08097_));
NAND_g _29394_ (.A(_08091_), .B(_08097_), .Y(_08098_));
AND_g _29395_ (.A(resetn), .B(_08098_), .Y(_00005_[5]));
NAND_g _29396_ (.A(mem_rdata[22]), .B(_01791_), .Y(_08099_));
NAND_g _29397_ (.A(mem_rdata[6]), .B(mem_la_wstrb[0]), .Y(_08100_));
NAND_g _29398_ (.A(mem_rdata[14]), .B(_07945_), .Y(_08101_));
NAND_g _29399_ (.A(mem_rdata[30]), .B(_01796_), .Y(_08102_));
AND_g _29400_ (.A(_08101_), .B(_08102_), .Y(_08103_));
AND_g _29401_ (.A(_08100_), .B(_08103_), .Y(_08104_));
NAND_g _29402_ (.A(_08099_), .B(_08104_), .Y(_08105_));
NAND_g _29403_ (.A(_07942_), .B(_08105_), .Y(_08106_));
NAND_g _29404_ (.A(instr_rdcycleh), .B(count_cycle[38]), .Y(_08107_));
NAND_g _29405_ (.A(count_instr[38]), .B(instr_rdinstrh), .Y(_08108_));
AND_g _29406_ (.A(_08107_), .B(_08108_), .Y(_08109_));
NAND_g _29407_ (.A(count_instr[6]), .B(instr_rdinstr), .Y(_08110_));
NAND_g _29408_ (.A(instr_rdcycle), .B(count_cycle[6]), .Y(_08111_));
AND_g _29409_ (.A(_08110_), .B(_08111_), .Y(_08112_));
NAND_g _29410_ (.A(_08109_), .B(_08112_), .Y(_08113_));
NAND_g _29411_ (.A(_10595_), .B(_08113_), .Y(_08114_));
NAND_g _29412_ (.A(pcpi_rs1[6]), .B(_13889_), .Y(_08115_));
AND_g _29413_ (.A(_08114_), .B(_08115_), .Y(_08116_));
AND_g _29414_ (.A(_08106_), .B(_08116_), .Y(_08117_));
NAND_g _29415_ (.A(_08093_), .B(_08095_), .Y(_08118_));
NAND_g _29416_ (.A(reg_pc[6]), .B(decoded_imm[6]), .Y(_08119_));
XOR_g _29417_ (.A(reg_pc[6]), .B(decoded_imm[6]), .Y(_08120_));
NAND_g _29418_ (.A(_08118_), .B(_08120_), .Y(_08121_));
XOR_g _29419_ (.A(_08118_), .B(_08120_), .Y(_08122_));
NAND_g _29420_ (.A(_14217_), .B(_08122_), .Y(_08123_));
NAND_g _29421_ (.A(_08117_), .B(_08123_), .Y(_08124_));
AND_g _29422_ (.A(resetn), .B(_08124_), .Y(_00005_[6]));
AND_g _29423_ (.A(_08119_), .B(_08121_), .Y(_08125_));
NAND_g _29424_ (.A(reg_pc[7]), .B(decoded_imm[7]), .Y(_08126_));
NOR_g _29425_ (.A(reg_pc[7]), .B(decoded_imm[7]), .Y(_08127_));
XOR_g _29426_ (.A(reg_pc[7]), .B(decoded_imm[7]), .Y(_08128_));
NAND_g _29427_ (.A(mem_rdata[23]), .B(_01791_), .Y(_08129_));
NAND_g _29428_ (.A(mem_rdata[31]), .B(_01796_), .Y(_08130_));
NAND_g _29429_ (.A(mem_rdata[15]), .B(_07945_), .Y(_08131_));
NAND_g _29430_ (.A(mem_rdata[7]), .B(mem_la_wstrb[0]), .Y(_08132_));
AND_g _29431_ (.A(_08131_), .B(_08132_), .Y(_08133_));
AND_g _29432_ (.A(_08130_), .B(_08133_), .Y(_08134_));
NAND_g _29433_ (.A(_08129_), .B(_08134_), .Y(_08135_));
NAND_g _29434_ (.A(_07942_), .B(_08135_), .Y(_08136_));
NAND_g _29435_ (.A(instr_rdcycleh), .B(count_cycle[39]), .Y(_08137_));
NAND_g _29436_ (.A(count_instr[39]), .B(instr_rdinstrh), .Y(_08138_));
AND_g _29437_ (.A(_08137_), .B(_08138_), .Y(_08139_));
NAND_g _29438_ (.A(count_instr[7]), .B(instr_rdinstr), .Y(_08140_));
NAND_g _29439_ (.A(instr_rdcycle), .B(count_cycle[7]), .Y(_08141_));
AND_g _29440_ (.A(_08140_), .B(_08141_), .Y(_08142_));
NAND_g _29441_ (.A(_08139_), .B(_08142_), .Y(_08143_));
NAND_g _29442_ (.A(_10595_), .B(_08143_), .Y(_08144_));
NAND_g _29443_ (.A(pcpi_rs1[7]), .B(_13889_), .Y(_08145_));
AND_g _29444_ (.A(_08144_), .B(_08145_), .Y(_08146_));
XNOR_g _29445_ (.A(_08125_), .B(_08128_), .Y(_08147_));
NAND_g _29446_ (.A(_14217_), .B(_08147_), .Y(_08148_));
AND_g _29447_ (.A(_08146_), .B(_08148_), .Y(_08149_));
NAND_g _29448_ (.A(_08136_), .B(_08149_), .Y(_08150_));
AND_g _29449_ (.A(resetn), .B(_08150_), .Y(_00005_[7]));
NAND_g _29450_ (.A(latched_is_lb), .B(_08135_), .Y(_08151_));
NAND_g _29451_ (.A(mem_rdata[24]), .B(_01789_), .Y(_08152_));
NAND_g _29452_ (.A(mem_rdata[8]), .B(_01780_), .Y(_08153_));
NAND_g _29453_ (.A(_08152_), .B(_08153_), .Y(_08154_));
NAND_g _29454_ (.A(_07938_), .B(_08154_), .Y(_08155_));
NAND_g _29455_ (.A(_08151_), .B(_08155_), .Y(_08156_));
NAND_g _29456_ (.A(_07941_), .B(_08156_), .Y(_08157_));
NAND_g _29457_ (.A(pcpi_rs1[8]), .B(_13889_), .Y(_08158_));
NAND_g _29458_ (.A(instr_rdcycleh), .B(count_cycle[40]), .Y(_08159_));
NAND_g _29459_ (.A(count_instr[40]), .B(instr_rdinstrh), .Y(_08160_));
AND_g _29460_ (.A(_08159_), .B(_08160_), .Y(_08161_));
NAND_g _29461_ (.A(count_instr[8]), .B(instr_rdinstr), .Y(_08162_));
NAND_g _29462_ (.A(instr_rdcycle), .B(count_cycle[8]), .Y(_08163_));
AND_g _29463_ (.A(_08162_), .B(_08163_), .Y(_08164_));
NAND_g _29464_ (.A(_08161_), .B(_08164_), .Y(_08165_));
NAND_g _29465_ (.A(_10595_), .B(_08165_), .Y(_08166_));
AND_g _29466_ (.A(_08158_), .B(_08166_), .Y(_08167_));
NAND_g _29467_ (.A(_08157_), .B(_08167_), .Y(_08168_));
NAND_g _29468_ (.A(reg_pc[8]), .B(decoded_imm[8]), .Y(_08169_));
XOR_g _29469_ (.A(reg_pc[8]), .B(decoded_imm[8]), .Y(_08170_));
AND_g _29470_ (.A(_08125_), .B(_08126_), .Y(_08171_));
NOR_g _29471_ (.A(_08127_), .B(_08171_), .Y(_08172_));
NAND_g _29472_ (.A(_08170_), .B(_08172_), .Y(_08173_));
NOR_g _29473_ (.A(_08170_), .B(_08172_), .Y(_08174_));
NAND_g _29474_ (.A(_14217_), .B(_08173_), .Y(_08175_));
NOR_g _29475_ (.A(_08174_), .B(_08175_), .Y(_08176_));
NOR_g _29476_ (.A(_08168_), .B(_08176_), .Y(_08177_));
NOR_g _29477_ (.A(_08811_), .B(_08177_), .Y(_00005_[8]));
NAND_g _29478_ (.A(mem_rdata[25]), .B(_01789_), .Y(_08178_));
NAND_g _29479_ (.A(mem_rdata[9]), .B(_01780_), .Y(_08179_));
NAND_g _29480_ (.A(_08178_), .B(_08179_), .Y(_08180_));
NAND_g _29481_ (.A(_07938_), .B(_08180_), .Y(_08181_));
NAND_g _29482_ (.A(_08151_), .B(_08181_), .Y(_08182_));
NAND_g _29483_ (.A(_07941_), .B(_08182_), .Y(_08183_));
NAND_g _29484_ (.A(instr_rdcycleh), .B(count_cycle[41]), .Y(_08184_));
NAND_g _29485_ (.A(count_instr[41]), .B(instr_rdinstrh), .Y(_08185_));
AND_g _29486_ (.A(_08184_), .B(_08185_), .Y(_08186_));
NAND_g _29487_ (.A(count_instr[9]), .B(instr_rdinstr), .Y(_08187_));
NAND_g _29488_ (.A(instr_rdcycle), .B(count_cycle[9]), .Y(_08188_));
AND_g _29489_ (.A(_08187_), .B(_08188_), .Y(_08189_));
NAND_g _29490_ (.A(_08186_), .B(_08189_), .Y(_08190_));
NAND_g _29491_ (.A(_10595_), .B(_08190_), .Y(_08191_));
NAND_g _29492_ (.A(pcpi_rs1[9]), .B(_13889_), .Y(_08192_));
AND_g _29493_ (.A(_08191_), .B(_08192_), .Y(_08193_));
AND_g _29494_ (.A(_08183_), .B(_08193_), .Y(_08194_));
AND_g _29495_ (.A(_08169_), .B(_08173_), .Y(_08195_));
NAND_g _29496_ (.A(reg_pc[9]), .B(decoded_imm[9]), .Y(_08196_));
NOR_g _29497_ (.A(reg_pc[9]), .B(decoded_imm[9]), .Y(_08197_));
XOR_g _29498_ (.A(reg_pc[9]), .B(decoded_imm[9]), .Y(_08198_));
XNOR_g _29499_ (.A(_08195_), .B(_08198_), .Y(_08199_));
NAND_g _29500_ (.A(_14217_), .B(_08199_), .Y(_08200_));
NAND_g _29501_ (.A(_08194_), .B(_08200_), .Y(_08201_));
AND_g _29502_ (.A(resetn), .B(_08201_), .Y(_00005_[9]));
NAND_g _29503_ (.A(mem_rdata[26]), .B(_01789_), .Y(_08202_));
NAND_g _29504_ (.A(mem_rdata[10]), .B(_01780_), .Y(_08203_));
NAND_g _29505_ (.A(_08202_), .B(_08203_), .Y(_08204_));
NAND_g _29506_ (.A(_07938_), .B(_08204_), .Y(_08205_));
NAND_g _29507_ (.A(_08151_), .B(_08205_), .Y(_08206_));
NAND_g _29508_ (.A(_07941_), .B(_08206_), .Y(_08207_));
NAND_g _29509_ (.A(instr_rdcycleh), .B(count_cycle[42]), .Y(_08208_));
NAND_g _29510_ (.A(count_instr[42]), .B(instr_rdinstrh), .Y(_08209_));
AND_g _29511_ (.A(_08208_), .B(_08209_), .Y(_08210_));
NAND_g _29512_ (.A(count_instr[10]), .B(instr_rdinstr), .Y(_08211_));
NAND_g _29513_ (.A(instr_rdcycle), .B(count_cycle[10]), .Y(_08212_));
AND_g _29514_ (.A(_08211_), .B(_08212_), .Y(_08213_));
NAND_g _29515_ (.A(_08210_), .B(_08213_), .Y(_08214_));
NAND_g _29516_ (.A(_10595_), .B(_08214_), .Y(_08215_));
NAND_g _29517_ (.A(pcpi_rs1[10]), .B(_13889_), .Y(_08216_));
NAND_g _29518_ (.A(_08215_), .B(_08216_), .Y(_08217_));
NAND_g _29519_ (.A(reg_pc[10]), .B(decoded_imm[10]), .Y(_08218_));
XOR_g _29520_ (.A(reg_pc[10]), .B(decoded_imm[10]), .Y(_08219_));
AND_g _29521_ (.A(_08195_), .B(_08196_), .Y(_08220_));
NOR_g _29522_ (.A(_08197_), .B(_08220_), .Y(_08221_));
NAND_g _29523_ (.A(_08219_), .B(_08221_), .Y(_08222_));
NOR_g _29524_ (.A(_08219_), .B(_08221_), .Y(_08223_));
NAND_g _29525_ (.A(_14217_), .B(_08222_), .Y(_08224_));
NOR_g _29526_ (.A(_08223_), .B(_08224_), .Y(_08225_));
NOR_g _29527_ (.A(_08217_), .B(_08225_), .Y(_08226_));
NAND_g _29528_ (.A(_08207_), .B(_08226_), .Y(_08227_));
AND_g _29529_ (.A(resetn), .B(_08227_), .Y(_00005_[10]));
AND_g _29530_ (.A(_08218_), .B(_08222_), .Y(_08228_));
NAND_g _29531_ (.A(reg_pc[11]), .B(decoded_imm[11]), .Y(_08229_));
NOR_g _29532_ (.A(reg_pc[11]), .B(decoded_imm[11]), .Y(_08230_));
XOR_g _29533_ (.A(reg_pc[11]), .B(decoded_imm[11]), .Y(_08231_));
NAND_g _29534_ (.A(mem_rdata[27]), .B(_01789_), .Y(_08232_));
NAND_g _29535_ (.A(mem_rdata[11]), .B(_01780_), .Y(_08233_));
NAND_g _29536_ (.A(_08232_), .B(_08233_), .Y(_08234_));
NAND_g _29537_ (.A(_07938_), .B(_08234_), .Y(_08235_));
NAND_g _29538_ (.A(_08151_), .B(_08235_), .Y(_08236_));
NAND_g _29539_ (.A(_07941_), .B(_08236_), .Y(_08237_));
NAND_g _29540_ (.A(instr_rdcycleh), .B(count_cycle[43]), .Y(_08238_));
NAND_g _29541_ (.A(count_instr[43]), .B(instr_rdinstrh), .Y(_08239_));
AND_g _29542_ (.A(_08238_), .B(_08239_), .Y(_08240_));
NAND_g _29543_ (.A(count_instr[11]), .B(instr_rdinstr), .Y(_08241_));
NAND_g _29544_ (.A(instr_rdcycle), .B(count_cycle[11]), .Y(_08242_));
AND_g _29545_ (.A(_08241_), .B(_08242_), .Y(_08243_));
NAND_g _29546_ (.A(_08240_), .B(_08243_), .Y(_08244_));
NAND_g _29547_ (.A(_10595_), .B(_08244_), .Y(_08245_));
NAND_g _29548_ (.A(pcpi_rs1[11]), .B(_13889_), .Y(_08246_));
AND_g _29549_ (.A(_08245_), .B(_08246_), .Y(_08247_));
XNOR_g _29550_ (.A(_08228_), .B(_08231_), .Y(_08248_));
NAND_g _29551_ (.A(_14217_), .B(_08248_), .Y(_08249_));
AND_g _29552_ (.A(_08247_), .B(_08249_), .Y(_08250_));
NAND_g _29553_ (.A(_08237_), .B(_08250_), .Y(_08251_));
AND_g _29554_ (.A(resetn), .B(_08251_), .Y(_00005_[11]));
NAND_g _29555_ (.A(mem_rdata[28]), .B(_01789_), .Y(_08252_));
NAND_g _29556_ (.A(mem_rdata[12]), .B(_01780_), .Y(_08253_));
NAND_g _29557_ (.A(_08252_), .B(_08253_), .Y(_08254_));
NAND_g _29558_ (.A(_07938_), .B(_08254_), .Y(_08255_));
NAND_g _29559_ (.A(_08151_), .B(_08255_), .Y(_08256_));
NAND_g _29560_ (.A(_07941_), .B(_08256_), .Y(_08257_));
NAND_g _29561_ (.A(instr_rdcycleh), .B(count_cycle[44]), .Y(_08258_));
NAND_g _29562_ (.A(count_instr[44]), .B(instr_rdinstrh), .Y(_08259_));
AND_g _29563_ (.A(_08258_), .B(_08259_), .Y(_08260_));
NAND_g _29564_ (.A(count_instr[12]), .B(instr_rdinstr), .Y(_08261_));
NAND_g _29565_ (.A(instr_rdcycle), .B(count_cycle[12]), .Y(_08262_));
AND_g _29566_ (.A(_08261_), .B(_08262_), .Y(_08263_));
NAND_g _29567_ (.A(_08260_), .B(_08263_), .Y(_08264_));
NAND_g _29568_ (.A(_10595_), .B(_08264_), .Y(_08265_));
NAND_g _29569_ (.A(pcpi_rs1[12]), .B(_13889_), .Y(_08266_));
AND_g _29570_ (.A(_08265_), .B(_08266_), .Y(_08267_));
NAND_g _29571_ (.A(_08257_), .B(_08267_), .Y(_08268_));
NAND_g _29572_ (.A(reg_pc[12]), .B(decoded_imm[12]), .Y(_08269_));
XOR_g _29573_ (.A(reg_pc[12]), .B(decoded_imm[12]), .Y(_08270_));
AND_g _29574_ (.A(_08228_), .B(_08229_), .Y(_08271_));
NOR_g _29575_ (.A(_08230_), .B(_08271_), .Y(_08272_));
NAND_g _29576_ (.A(_08270_), .B(_08272_), .Y(_08273_));
NOR_g _29577_ (.A(_08270_), .B(_08272_), .Y(_08274_));
NAND_g _29578_ (.A(_14217_), .B(_08273_), .Y(_08275_));
NOR_g _29579_ (.A(_08274_), .B(_08275_), .Y(_08276_));
NOR_g _29580_ (.A(_08268_), .B(_08276_), .Y(_08277_));
NOR_g _29581_ (.A(_08811_), .B(_08277_), .Y(_00005_[12]));
AND_g _29582_ (.A(_08269_), .B(_08273_), .Y(_08278_));
NAND_g _29583_ (.A(reg_pc[13]), .B(decoded_imm[13]), .Y(_08279_));
NOR_g _29584_ (.A(reg_pc[13]), .B(decoded_imm[13]), .Y(_08280_));
XNOR_g _29585_ (.A(reg_pc[13]), .B(decoded_imm[13]), .Y(_08281_));
NOR_g _29586_ (.A(_08278_), .B(_08281_), .Y(_08282_));
NAND_g _29587_ (.A(_08278_), .B(_08281_), .Y(_08283_));
NAND_g _29588_ (.A(mem_rdata[29]), .B(_01789_), .Y(_08284_));
NAND_g _29589_ (.A(mem_rdata[13]), .B(_01780_), .Y(_08285_));
NAND_g _29590_ (.A(_08284_), .B(_08285_), .Y(_08286_));
NAND_g _29591_ (.A(_07938_), .B(_08286_), .Y(_08287_));
NAND_g _29592_ (.A(_08151_), .B(_08287_), .Y(_08288_));
NAND_g _29593_ (.A(_07941_), .B(_08288_), .Y(_08289_));
NAND_g _29594_ (.A(instr_rdcycleh), .B(count_cycle[45]), .Y(_08290_));
NAND_g _29595_ (.A(count_instr[45]), .B(instr_rdinstrh), .Y(_08291_));
AND_g _29596_ (.A(_08290_), .B(_08291_), .Y(_08292_));
NAND_g _29597_ (.A(count_instr[13]), .B(instr_rdinstr), .Y(_08293_));
NAND_g _29598_ (.A(instr_rdcycle), .B(count_cycle[13]), .Y(_08294_));
AND_g _29599_ (.A(_08293_), .B(_08294_), .Y(_08295_));
NAND_g _29600_ (.A(_08292_), .B(_08295_), .Y(_08296_));
NAND_g _29601_ (.A(_10595_), .B(_08296_), .Y(_08297_));
NAND_g _29602_ (.A(pcpi_rs1[13]), .B(_13889_), .Y(_08298_));
AND_g _29603_ (.A(_08297_), .B(_08298_), .Y(_08299_));
NOR_g _29604_ (.A(_14218_), .B(_08282_), .Y(_08300_));
NAND_g _29605_ (.A(_08283_), .B(_08300_), .Y(_08301_));
AND_g _29606_ (.A(_08299_), .B(_08301_), .Y(_08302_));
NAND_g _29607_ (.A(_08289_), .B(_08302_), .Y(_08303_));
AND_g _29608_ (.A(resetn), .B(_08303_), .Y(_00005_[13]));
NAND_g _29609_ (.A(mem_rdata[30]), .B(_01789_), .Y(_08304_));
NAND_g _29610_ (.A(mem_rdata[14]), .B(_01780_), .Y(_08305_));
NAND_g _29611_ (.A(_08304_), .B(_08305_), .Y(_08306_));
NAND_g _29612_ (.A(_07938_), .B(_08306_), .Y(_08307_));
NAND_g _29613_ (.A(_08151_), .B(_08307_), .Y(_08308_));
NAND_g _29614_ (.A(_07941_), .B(_08308_), .Y(_08309_));
NAND_g _29615_ (.A(pcpi_rs1[14]), .B(_13889_), .Y(_08310_));
NAND_g _29616_ (.A(instr_rdcycleh), .B(count_cycle[46]), .Y(_08311_));
NAND_g _29617_ (.A(count_instr[46]), .B(instr_rdinstrh), .Y(_08312_));
AND_g _29618_ (.A(_08311_), .B(_08312_), .Y(_08313_));
NAND_g _29619_ (.A(count_instr[14]), .B(instr_rdinstr), .Y(_08314_));
NAND_g _29620_ (.A(instr_rdcycle), .B(count_cycle[14]), .Y(_08315_));
AND_g _29621_ (.A(_08314_), .B(_08315_), .Y(_08316_));
NAND_g _29622_ (.A(_08313_), .B(_08316_), .Y(_08317_));
NAND_g _29623_ (.A(_10595_), .B(_08317_), .Y(_08318_));
AND_g _29624_ (.A(_08310_), .B(_08318_), .Y(_08319_));
NAND_g _29625_ (.A(_08309_), .B(_08319_), .Y(_08320_));
NAND_g _29626_ (.A(reg_pc[14]), .B(decoded_imm[14]), .Y(_08321_));
XOR_g _29627_ (.A(reg_pc[14]), .B(decoded_imm[14]), .Y(_08322_));
AND_g _29628_ (.A(_08278_), .B(_08279_), .Y(_08323_));
NOR_g _29629_ (.A(_08280_), .B(_08323_), .Y(_08324_));
NAND_g _29630_ (.A(_08322_), .B(_08324_), .Y(_08325_));
NOR_g _29631_ (.A(_08322_), .B(_08324_), .Y(_08326_));
NAND_g _29632_ (.A(_14217_), .B(_08325_), .Y(_08327_));
NOR_g _29633_ (.A(_08326_), .B(_08327_), .Y(_08328_));
NOR_g _29634_ (.A(_08320_), .B(_08328_), .Y(_08329_));
NOR_g _29635_ (.A(_08811_), .B(_08329_), .Y(_00005_[14]));
AND_g _29636_ (.A(_08321_), .B(_08325_), .Y(_08330_));
NAND_g _29637_ (.A(reg_pc[15]), .B(decoded_imm[15]), .Y(_08331_));
NOR_g _29638_ (.A(reg_pc[15]), .B(decoded_imm[15]), .Y(_08332_));
XNOR_g _29639_ (.A(reg_pc[15]), .B(decoded_imm[15]), .Y(_08333_));
NOR_g _29640_ (.A(_08330_), .B(_08333_), .Y(_08334_));
NAND_g _29641_ (.A(_08330_), .B(_08333_), .Y(_08335_));
NAND_g _29642_ (.A(mem_rdata[31]), .B(_01789_), .Y(_08336_));
NAND_g _29643_ (.A(mem_rdata[15]), .B(_01780_), .Y(_08337_));
NAND_g _29644_ (.A(_08336_), .B(_08337_), .Y(_08338_));
NAND_g _29645_ (.A(_07938_), .B(_08338_), .Y(_08339_));
NAND_g _29646_ (.A(_08151_), .B(_08339_), .Y(_08340_));
NAND_g _29647_ (.A(_07941_), .B(_08340_), .Y(_08341_));
NAND_g _29648_ (.A(instr_rdcycleh), .B(count_cycle[47]), .Y(_08342_));
NAND_g _29649_ (.A(count_instr[47]), .B(instr_rdinstrh), .Y(_08343_));
AND_g _29650_ (.A(_08342_), .B(_08343_), .Y(_08344_));
NAND_g _29651_ (.A(count_instr[15]), .B(instr_rdinstr), .Y(_08345_));
NAND_g _29652_ (.A(instr_rdcycle), .B(count_cycle[15]), .Y(_08346_));
AND_g _29653_ (.A(_08345_), .B(_08346_), .Y(_08347_));
NAND_g _29654_ (.A(_08344_), .B(_08347_), .Y(_08348_));
NAND_g _29655_ (.A(_10595_), .B(_08348_), .Y(_08349_));
NAND_g _29656_ (.A(pcpi_rs1[15]), .B(_13889_), .Y(_08350_));
AND_g _29657_ (.A(_08349_), .B(_08350_), .Y(_08351_));
NOR_g _29658_ (.A(_14218_), .B(_08334_), .Y(_08352_));
NAND_g _29659_ (.A(_08335_), .B(_08352_), .Y(_08353_));
AND_g _29660_ (.A(_08351_), .B(_08353_), .Y(_08354_));
NAND_g _29661_ (.A(_08341_), .B(_08354_), .Y(_08355_));
AND_g _29662_ (.A(resetn), .B(_08355_), .Y(_00005_[15]));
NAND_g _29663_ (.A(reg_pc[16]), .B(decoded_imm[16]), .Y(_08356_));
XOR_g _29664_ (.A(reg_pc[16]), .B(decoded_imm[16]), .Y(_08357_));
AND_g _29665_ (.A(_08330_), .B(_08331_), .Y(_08358_));
NOR_g _29666_ (.A(_08332_), .B(_08358_), .Y(_08359_));
NAND_g _29667_ (.A(_08357_), .B(_08359_), .Y(_08360_));
NAND_g _29668_ (.A(latched_is_lh), .B(_08338_), .Y(_08361_));
AND_g _29669_ (.A(_08151_), .B(_08361_), .Y(_08362_));
AND_g _29670_ (.A(latched_is_lu), .B(mem_rdata[16]), .Y(_08363_));
NAND_g _29671_ (.A(_01700_), .B(_08363_), .Y(_08364_));
NAND_g _29672_ (.A(_08362_), .B(_08364_), .Y(_08365_));
NAND_g _29673_ (.A(_07941_), .B(_08365_), .Y(_08366_));
NAND_g _29674_ (.A(instr_rdcycleh), .B(count_cycle[48]), .Y(_08367_));
NAND_g _29675_ (.A(count_instr[48]), .B(instr_rdinstrh), .Y(_08368_));
AND_g _29676_ (.A(_08367_), .B(_08368_), .Y(_08369_));
NAND_g _29677_ (.A(count_instr[16]), .B(instr_rdinstr), .Y(_08370_));
NAND_g _29678_ (.A(instr_rdcycle), .B(count_cycle[16]), .Y(_08371_));
AND_g _29679_ (.A(_08370_), .B(_08371_), .Y(_08372_));
NAND_g _29680_ (.A(_08369_), .B(_08372_), .Y(_08373_));
NAND_g _29681_ (.A(_10595_), .B(_08373_), .Y(_08374_));
NAND_g _29682_ (.A(pcpi_rs1[16]), .B(_13889_), .Y(_08375_));
AND_g _29683_ (.A(_08374_), .B(_08375_), .Y(_08376_));
XOR_g _29684_ (.A(_08357_), .B(_08359_), .Y(_08377_));
NAND_g _29685_ (.A(_14217_), .B(_08377_), .Y(_08378_));
AND_g _29686_ (.A(_08376_), .B(_08378_), .Y(_08379_));
NAND_g _29687_ (.A(_08366_), .B(_08379_), .Y(_08380_));
AND_g _29688_ (.A(resetn), .B(_08380_), .Y(_00005_[16]));
AND_g _29689_ (.A(_08356_), .B(_08360_), .Y(_08381_));
NAND_g _29690_ (.A(reg_pc[17]), .B(decoded_imm[17]), .Y(_08382_));
NOR_g _29691_ (.A(reg_pc[17]), .B(decoded_imm[17]), .Y(_08383_));
XNOR_g _29692_ (.A(reg_pc[17]), .B(decoded_imm[17]), .Y(_08384_));
NOR_g _29693_ (.A(_08381_), .B(_08384_), .Y(_08385_));
NAND_g _29694_ (.A(_08381_), .B(_08384_), .Y(_08386_));
AND_g _29695_ (.A(latched_is_lu), .B(mem_rdata[17]), .Y(_08387_));
NAND_g _29696_ (.A(_01700_), .B(_08387_), .Y(_08388_));
NAND_g _29697_ (.A(_08362_), .B(_08388_), .Y(_08389_));
NAND_g _29698_ (.A(_07941_), .B(_08389_), .Y(_08390_));
NAND_g _29699_ (.A(instr_rdcycleh), .B(count_cycle[49]), .Y(_08391_));
NAND_g _29700_ (.A(count_instr[49]), .B(instr_rdinstrh), .Y(_08392_));
AND_g _29701_ (.A(_08391_), .B(_08392_), .Y(_08393_));
NAND_g _29702_ (.A(count_instr[17]), .B(instr_rdinstr), .Y(_08394_));
NAND_g _29703_ (.A(instr_rdcycle), .B(count_cycle[17]), .Y(_08395_));
AND_g _29704_ (.A(_08394_), .B(_08395_), .Y(_08396_));
NAND_g _29705_ (.A(_08393_), .B(_08396_), .Y(_08397_));
NAND_g _29706_ (.A(_10595_), .B(_08397_), .Y(_08398_));
NAND_g _29707_ (.A(pcpi_rs1[17]), .B(_13889_), .Y(_08399_));
AND_g _29708_ (.A(_08398_), .B(_08399_), .Y(_08400_));
NOR_g _29709_ (.A(_14218_), .B(_08385_), .Y(_08401_));
NAND_g _29710_ (.A(_08386_), .B(_08401_), .Y(_08402_));
AND_g _29711_ (.A(_08400_), .B(_08402_), .Y(_08403_));
NAND_g _29712_ (.A(_08390_), .B(_08403_), .Y(_08404_));
AND_g _29713_ (.A(resetn), .B(_08404_), .Y(_00005_[17]));
AND_g _29714_ (.A(latched_is_lu), .B(mem_rdata[18]), .Y(_08405_));
NAND_g _29715_ (.A(_01700_), .B(_08405_), .Y(_08406_));
NAND_g _29716_ (.A(_08362_), .B(_08406_), .Y(_08407_));
NAND_g _29717_ (.A(_07941_), .B(_08407_), .Y(_08408_));
NAND_g _29718_ (.A(instr_rdcycleh), .B(count_cycle[50]), .Y(_08409_));
NAND_g _29719_ (.A(count_instr[50]), .B(instr_rdinstrh), .Y(_08410_));
AND_g _29720_ (.A(_08409_), .B(_08410_), .Y(_08411_));
NAND_g _29721_ (.A(count_instr[18]), .B(instr_rdinstr), .Y(_08412_));
NAND_g _29722_ (.A(instr_rdcycle), .B(count_cycle[18]), .Y(_08413_));
AND_g _29723_ (.A(_08412_), .B(_08413_), .Y(_08414_));
NAND_g _29724_ (.A(_08411_), .B(_08414_), .Y(_08415_));
NAND_g _29725_ (.A(_10595_), .B(_08415_), .Y(_08416_));
NAND_g _29726_ (.A(pcpi_rs1[18]), .B(_13889_), .Y(_08417_));
AND_g _29727_ (.A(_08416_), .B(_08417_), .Y(_08418_));
NAND_g _29728_ (.A(_08408_), .B(_08418_), .Y(_08419_));
NAND_g _29729_ (.A(reg_pc[18]), .B(decoded_imm[18]), .Y(_08420_));
XOR_g _29730_ (.A(reg_pc[18]), .B(decoded_imm[18]), .Y(_08421_));
AND_g _29731_ (.A(_08381_), .B(_08382_), .Y(_08422_));
NOR_g _29732_ (.A(_08383_), .B(_08422_), .Y(_08423_));
NAND_g _29733_ (.A(_08421_), .B(_08423_), .Y(_08424_));
NOR_g _29734_ (.A(_08421_), .B(_08423_), .Y(_08425_));
NAND_g _29735_ (.A(_14217_), .B(_08424_), .Y(_08426_));
NOR_g _29736_ (.A(_08425_), .B(_08426_), .Y(_08427_));
NOR_g _29737_ (.A(_08419_), .B(_08427_), .Y(_08428_));
NOR_g _29738_ (.A(_08811_), .B(_08428_), .Y(_00005_[18]));
AND_g _29739_ (.A(_08420_), .B(_08424_), .Y(_08429_));
NAND_g _29740_ (.A(reg_pc[19]), .B(decoded_imm[19]), .Y(_08430_));
NOR_g _29741_ (.A(reg_pc[19]), .B(decoded_imm[19]), .Y(_08431_));
XNOR_g _29742_ (.A(reg_pc[19]), .B(decoded_imm[19]), .Y(_08432_));
NOR_g _29743_ (.A(_08429_), .B(_08432_), .Y(_08433_));
NAND_g _29744_ (.A(_08429_), .B(_08432_), .Y(_08434_));
AND_g _29745_ (.A(latched_is_lu), .B(mem_rdata[19]), .Y(_08435_));
NAND_g _29746_ (.A(_01700_), .B(_08435_), .Y(_08436_));
NAND_g _29747_ (.A(_08362_), .B(_08436_), .Y(_08437_));
NAND_g _29748_ (.A(_07941_), .B(_08437_), .Y(_08438_));
NAND_g _29749_ (.A(pcpi_rs1[19]), .B(_13889_), .Y(_08439_));
NAND_g _29750_ (.A(instr_rdcycleh), .B(count_cycle[51]), .Y(_08440_));
NAND_g _29751_ (.A(count_instr[51]), .B(instr_rdinstrh), .Y(_08441_));
AND_g _29752_ (.A(_08440_), .B(_08441_), .Y(_08442_));
NAND_g _29753_ (.A(count_instr[19]), .B(instr_rdinstr), .Y(_08443_));
NAND_g _29754_ (.A(instr_rdcycle), .B(count_cycle[19]), .Y(_08444_));
AND_g _29755_ (.A(_08443_), .B(_08444_), .Y(_08445_));
NAND_g _29756_ (.A(_08442_), .B(_08445_), .Y(_08446_));
NAND_g _29757_ (.A(_10595_), .B(_08446_), .Y(_08447_));
AND_g _29758_ (.A(_08439_), .B(_08447_), .Y(_08448_));
NOR_g _29759_ (.A(_14218_), .B(_08433_), .Y(_08449_));
NAND_g _29760_ (.A(_08434_), .B(_08449_), .Y(_08450_));
AND_g _29761_ (.A(_08448_), .B(_08450_), .Y(_08451_));
NAND_g _29762_ (.A(_08438_), .B(_08451_), .Y(_08452_));
AND_g _29763_ (.A(resetn), .B(_08452_), .Y(_00005_[19]));
NAND_g _29764_ (.A(reg_pc[20]), .B(decoded_imm[20]), .Y(_08453_));
XOR_g _29765_ (.A(reg_pc[20]), .B(decoded_imm[20]), .Y(_08454_));
AND_g _29766_ (.A(_08429_), .B(_08430_), .Y(_08455_));
NOR_g _29767_ (.A(_08431_), .B(_08455_), .Y(_08456_));
NAND_g _29768_ (.A(_08454_), .B(_08456_), .Y(_08457_));
AND_g _29769_ (.A(latched_is_lu), .B(mem_rdata[20]), .Y(_08458_));
NAND_g _29770_ (.A(_01700_), .B(_08458_), .Y(_08459_));
NAND_g _29771_ (.A(_08362_), .B(_08459_), .Y(_08460_));
NAND_g _29772_ (.A(_07941_), .B(_08460_), .Y(_08461_));
NAND_g _29773_ (.A(instr_rdcycleh), .B(count_cycle[52]), .Y(_08462_));
NAND_g _29774_ (.A(count_instr[52]), .B(instr_rdinstrh), .Y(_08463_));
AND_g _29775_ (.A(_08462_), .B(_08463_), .Y(_08464_));
NAND_g _29776_ (.A(count_instr[20]), .B(instr_rdinstr), .Y(_08465_));
NAND_g _29777_ (.A(instr_rdcycle), .B(count_cycle[20]), .Y(_08466_));
AND_g _29778_ (.A(_08465_), .B(_08466_), .Y(_08467_));
NAND_g _29779_ (.A(_08464_), .B(_08467_), .Y(_08468_));
NAND_g _29780_ (.A(_10595_), .B(_08468_), .Y(_08469_));
NAND_g _29781_ (.A(pcpi_rs1[20]), .B(_13889_), .Y(_08470_));
AND_g _29782_ (.A(_08469_), .B(_08470_), .Y(_08471_));
XOR_g _29783_ (.A(_08454_), .B(_08456_), .Y(_08472_));
NAND_g _29784_ (.A(_14217_), .B(_08472_), .Y(_08473_));
AND_g _29785_ (.A(_08471_), .B(_08473_), .Y(_08474_));
NAND_g _29786_ (.A(_08461_), .B(_08474_), .Y(_08475_));
AND_g _29787_ (.A(resetn), .B(_08475_), .Y(_00005_[20]));
AND_g _29788_ (.A(_08453_), .B(_08457_), .Y(_08476_));
NAND_g _29789_ (.A(reg_pc[21]), .B(decoded_imm[21]), .Y(_08477_));
NOR_g _29790_ (.A(reg_pc[21]), .B(decoded_imm[21]), .Y(_08478_));
XNOR_g _29791_ (.A(reg_pc[21]), .B(decoded_imm[21]), .Y(_08479_));
NOR_g _29792_ (.A(_08476_), .B(_08479_), .Y(_08480_));
NAND_g _29793_ (.A(_08476_), .B(_08479_), .Y(_08481_));
AND_g _29794_ (.A(latched_is_lu), .B(mem_rdata[21]), .Y(_08482_));
NAND_g _29795_ (.A(_01700_), .B(_08482_), .Y(_08483_));
NAND_g _29796_ (.A(_08362_), .B(_08483_), .Y(_08484_));
NAND_g _29797_ (.A(_07941_), .B(_08484_), .Y(_08485_));
NAND_g _29798_ (.A(instr_rdcycleh), .B(count_cycle[53]), .Y(_08486_));
NAND_g _29799_ (.A(count_instr[53]), .B(instr_rdinstrh), .Y(_08487_));
AND_g _29800_ (.A(_08486_), .B(_08487_), .Y(_08488_));
NAND_g _29801_ (.A(count_instr[21]), .B(instr_rdinstr), .Y(_08489_));
NAND_g _29802_ (.A(instr_rdcycle), .B(count_cycle[21]), .Y(_08490_));
AND_g _29803_ (.A(_08489_), .B(_08490_), .Y(_08491_));
NAND_g _29804_ (.A(_08488_), .B(_08491_), .Y(_08492_));
NAND_g _29805_ (.A(_10595_), .B(_08492_), .Y(_08493_));
NAND_g _29806_ (.A(pcpi_rs1[21]), .B(_13889_), .Y(_08494_));
AND_g _29807_ (.A(_08493_), .B(_08494_), .Y(_08495_));
NOR_g _29808_ (.A(_14218_), .B(_08480_), .Y(_08496_));
NAND_g _29809_ (.A(_08481_), .B(_08496_), .Y(_08497_));
AND_g _29810_ (.A(_08495_), .B(_08497_), .Y(_08498_));
NAND_g _29811_ (.A(_08485_), .B(_08498_), .Y(_08499_));
AND_g _29812_ (.A(resetn), .B(_08499_), .Y(_00005_[21]));
NAND_g _29813_ (.A(reg_pc[22]), .B(decoded_imm[22]), .Y(_08500_));
XOR_g _29814_ (.A(reg_pc[22]), .B(decoded_imm[22]), .Y(_08501_));
AND_g _29815_ (.A(_08476_), .B(_08477_), .Y(_08502_));
NOR_g _29816_ (.A(_08478_), .B(_08502_), .Y(_08503_));
NAND_g _29817_ (.A(_08501_), .B(_08503_), .Y(_08504_));
NOR_g _29818_ (.A(_08501_), .B(_08503_), .Y(_08505_));
NOR_g _29819_ (.A(_14215_), .B(_08505_), .Y(_08506_));
NAND_g _29820_ (.A(_08504_), .B(_08506_), .Y(_08507_));
AND_g _29821_ (.A(latched_is_lu), .B(mem_rdata[22]), .Y(_08508_));
NAND_g _29822_ (.A(_01700_), .B(_08508_), .Y(_08509_));
NAND_g _29823_ (.A(_08362_), .B(_08509_), .Y(_08510_));
NAND_g _29824_ (.A(_07941_), .B(_08510_), .Y(_08511_));
NAND_g _29825_ (.A(instr_rdcycleh), .B(count_cycle[54]), .Y(_08512_));
NAND_g _29826_ (.A(count_instr[54]), .B(instr_rdinstrh), .Y(_08513_));
AND_g _29827_ (.A(_08512_), .B(_08513_), .Y(_08514_));
NAND_g _29828_ (.A(count_instr[22]), .B(instr_rdinstr), .Y(_08515_));
NAND_g _29829_ (.A(instr_rdcycle), .B(count_cycle[22]), .Y(_08516_));
AND_g _29830_ (.A(_08515_), .B(_08516_), .Y(_08517_));
NAND_g _29831_ (.A(_08514_), .B(_08517_), .Y(_08518_));
NAND_g _29832_ (.A(_10595_), .B(_08518_), .Y(_08519_));
NAND_g _29833_ (.A(pcpi_rs1[22]), .B(_13889_), .Y(_08520_));
AND_g _29834_ (.A(_08519_), .B(_08520_), .Y(_08521_));
AND_g _29835_ (.A(_08511_), .B(_08521_), .Y(_08522_));
NAND_g _29836_ (.A(_08507_), .B(_08522_), .Y(_08523_));
AND_g _29837_ (.A(resetn), .B(_08523_), .Y(_00005_[22]));
AND_g _29838_ (.A(_08500_), .B(_08504_), .Y(_08524_));
NAND_g _29839_ (.A(reg_pc[23]), .B(decoded_imm[23]), .Y(_08525_));
NOR_g _29840_ (.A(reg_pc[23]), .B(decoded_imm[23]), .Y(_08526_));
XNOR_g _29841_ (.A(reg_pc[23]), .B(decoded_imm[23]), .Y(_08527_));
NOR_g _29842_ (.A(_08524_), .B(_08527_), .Y(_08528_));
NAND_g _29843_ (.A(_08524_), .B(_08527_), .Y(_08529_));
AND_g _29844_ (.A(latched_is_lu), .B(mem_rdata[23]), .Y(_08530_));
NAND_g _29845_ (.A(_01700_), .B(_08530_), .Y(_08531_));
NAND_g _29846_ (.A(_08362_), .B(_08531_), .Y(_08532_));
NAND_g _29847_ (.A(_07941_), .B(_08532_), .Y(_08533_));
NAND_g _29848_ (.A(pcpi_rs1[23]), .B(_13889_), .Y(_08534_));
NAND_g _29849_ (.A(instr_rdcycleh), .B(count_cycle[55]), .Y(_08535_));
NAND_g _29850_ (.A(count_instr[55]), .B(instr_rdinstrh), .Y(_08536_));
AND_g _29851_ (.A(_08535_), .B(_08536_), .Y(_08537_));
NAND_g _29852_ (.A(count_instr[23]), .B(instr_rdinstr), .Y(_08538_));
NAND_g _29853_ (.A(instr_rdcycle), .B(count_cycle[23]), .Y(_08539_));
AND_g _29854_ (.A(_08538_), .B(_08539_), .Y(_08540_));
NAND_g _29855_ (.A(_08537_), .B(_08540_), .Y(_08541_));
NAND_g _29856_ (.A(_10595_), .B(_08541_), .Y(_08542_));
AND_g _29857_ (.A(_08534_), .B(_08542_), .Y(_08543_));
NOR_g _29858_ (.A(_14218_), .B(_08528_), .Y(_08544_));
NAND_g _29859_ (.A(_08529_), .B(_08544_), .Y(_08545_));
AND_g _29860_ (.A(_08543_), .B(_08545_), .Y(_08546_));
NAND_g _29861_ (.A(_08533_), .B(_08546_), .Y(_08547_));
AND_g _29862_ (.A(resetn), .B(_08547_), .Y(_00005_[23]));
AND_g _29863_ (.A(latched_is_lu), .B(mem_rdata[24]), .Y(_08548_));
NAND_g _29864_ (.A(_01700_), .B(_08548_), .Y(_08549_));
NAND_g _29865_ (.A(_08362_), .B(_08549_), .Y(_08550_));
NAND_g _29866_ (.A(_07941_), .B(_08550_), .Y(_08551_));
NAND_g _29867_ (.A(instr_rdcycleh), .B(count_cycle[56]), .Y(_08552_));
NAND_g _29868_ (.A(count_instr[56]), .B(instr_rdinstrh), .Y(_08553_));
AND_g _29869_ (.A(_08552_), .B(_08553_), .Y(_08554_));
NAND_g _29870_ (.A(count_instr[24]), .B(instr_rdinstr), .Y(_08555_));
NAND_g _29871_ (.A(instr_rdcycle), .B(count_cycle[24]), .Y(_08556_));
AND_g _29872_ (.A(_08555_), .B(_08556_), .Y(_08557_));
NAND_g _29873_ (.A(_08554_), .B(_08557_), .Y(_08558_));
NAND_g _29874_ (.A(_10595_), .B(_08558_), .Y(_08559_));
NAND_g _29875_ (.A(pcpi_rs1[24]), .B(_13889_), .Y(_08560_));
AND_g _29876_ (.A(_08559_), .B(_08560_), .Y(_08561_));
NAND_g _29877_ (.A(_08551_), .B(_08561_), .Y(_08562_));
NAND_g _29878_ (.A(reg_pc[24]), .B(decoded_imm[24]), .Y(_08563_));
XOR_g _29879_ (.A(reg_pc[24]), .B(decoded_imm[24]), .Y(_08564_));
AND_g _29880_ (.A(_08524_), .B(_08525_), .Y(_08565_));
NOR_g _29881_ (.A(_08526_), .B(_08565_), .Y(_08566_));
NAND_g _29882_ (.A(_08564_), .B(_08566_), .Y(_08567_));
NOR_g _29883_ (.A(_08564_), .B(_08566_), .Y(_08568_));
NAND_g _29884_ (.A(_14217_), .B(_08567_), .Y(_08569_));
NOR_g _29885_ (.A(_08568_), .B(_08569_), .Y(_08570_));
NOR_g _29886_ (.A(_08562_), .B(_08570_), .Y(_08571_));
NOR_g _29887_ (.A(_08811_), .B(_08571_), .Y(_00005_[24]));
AND_g _29888_ (.A(latched_is_lu), .B(mem_rdata[25]), .Y(_08572_));
NAND_g _29889_ (.A(_01700_), .B(_08572_), .Y(_08573_));
NAND_g _29890_ (.A(_08362_), .B(_08573_), .Y(_08574_));
NAND_g _29891_ (.A(_07941_), .B(_08574_), .Y(_08575_));
NAND_g _29892_ (.A(instr_rdcycleh), .B(count_cycle[57]), .Y(_08576_));
NAND_g _29893_ (.A(count_instr[57]), .B(instr_rdinstrh), .Y(_08577_));
AND_g _29894_ (.A(_08576_), .B(_08577_), .Y(_08578_));
NAND_g _29895_ (.A(count_instr[25]), .B(instr_rdinstr), .Y(_08579_));
NAND_g _29896_ (.A(instr_rdcycle), .B(count_cycle[25]), .Y(_08580_));
AND_g _29897_ (.A(_08579_), .B(_08580_), .Y(_08581_));
NAND_g _29898_ (.A(_08578_), .B(_08581_), .Y(_08582_));
NAND_g _29899_ (.A(_10595_), .B(_08582_), .Y(_08583_));
NAND_g _29900_ (.A(pcpi_rs1[25]), .B(_13889_), .Y(_08584_));
AND_g _29901_ (.A(_08583_), .B(_08584_), .Y(_08585_));
AND_g _29902_ (.A(_08575_), .B(_08585_), .Y(_08586_));
AND_g _29903_ (.A(_08563_), .B(_08567_), .Y(_08587_));
NAND_g _29904_ (.A(reg_pc[25]), .B(decoded_imm[25]), .Y(_08588_));
NOR_g _29905_ (.A(reg_pc[25]), .B(decoded_imm[25]), .Y(_08589_));
XOR_g _29906_ (.A(reg_pc[25]), .B(decoded_imm[25]), .Y(_08590_));
XNOR_g _29907_ (.A(_08587_), .B(_08590_), .Y(_08591_));
NAND_g _29908_ (.A(_14217_), .B(_08591_), .Y(_08592_));
NAND_g _29909_ (.A(_08586_), .B(_08592_), .Y(_08593_));
AND_g _29910_ (.A(resetn), .B(_08593_), .Y(_00005_[25]));
NAND_g _29911_ (.A(reg_pc[26]), .B(decoded_imm[26]), .Y(_08594_));
XOR_g _29912_ (.A(reg_pc[26]), .B(decoded_imm[26]), .Y(_08595_));
AND_g _29913_ (.A(_08587_), .B(_08588_), .Y(_08596_));
NOR_g _29914_ (.A(_08589_), .B(_08596_), .Y(_08597_));
NAND_g _29915_ (.A(_08595_), .B(_08597_), .Y(_08598_));
AND_g _29916_ (.A(latched_is_lu), .B(mem_rdata[26]), .Y(_08599_));
NAND_g _29917_ (.A(_01700_), .B(_08599_), .Y(_08600_));
NAND_g _29918_ (.A(_08362_), .B(_08600_), .Y(_08601_));
NAND_g _29919_ (.A(_07941_), .B(_08601_), .Y(_08602_));
NAND_g _29920_ (.A(instr_rdcycleh), .B(count_cycle[58]), .Y(_08603_));
NAND_g _29921_ (.A(count_instr[58]), .B(instr_rdinstrh), .Y(_08604_));
AND_g _29922_ (.A(_08603_), .B(_08604_), .Y(_08605_));
NAND_g _29923_ (.A(count_instr[26]), .B(instr_rdinstr), .Y(_08606_));
NAND_g _29924_ (.A(instr_rdcycle), .B(count_cycle[26]), .Y(_08607_));
AND_g _29925_ (.A(_08606_), .B(_08607_), .Y(_08608_));
NAND_g _29926_ (.A(_08605_), .B(_08608_), .Y(_08609_));
NAND_g _29927_ (.A(_10595_), .B(_08609_), .Y(_08610_));
NAND_g _29928_ (.A(pcpi_rs1[26]), .B(_13889_), .Y(_08611_));
AND_g _29929_ (.A(_08610_), .B(_08611_), .Y(_08612_));
XOR_g _29930_ (.A(_08595_), .B(_08597_), .Y(_08613_));
NAND_g _29931_ (.A(_14217_), .B(_08613_), .Y(_08614_));
AND_g _29932_ (.A(_08612_), .B(_08614_), .Y(_08615_));
NAND_g _29933_ (.A(_08602_), .B(_08615_), .Y(_08616_));
AND_g _29934_ (.A(resetn), .B(_08616_), .Y(_00005_[26]));
AND_g _29935_ (.A(_08594_), .B(_08598_), .Y(_08617_));
NAND_g _29936_ (.A(reg_pc[27]), .B(decoded_imm[27]), .Y(_08618_));
NOR_g _29937_ (.A(reg_pc[27]), .B(decoded_imm[27]), .Y(_08619_));
XNOR_g _29938_ (.A(reg_pc[27]), .B(decoded_imm[27]), .Y(_08620_));
NOR_g _29939_ (.A(_08617_), .B(_08620_), .Y(_08621_));
NAND_g _29940_ (.A(_08617_), .B(_08620_), .Y(_08622_));
AND_g _29941_ (.A(latched_is_lu), .B(mem_rdata[27]), .Y(_08623_));
NAND_g _29942_ (.A(_01700_), .B(_08623_), .Y(_08624_));
NAND_g _29943_ (.A(_08362_), .B(_08624_), .Y(_08625_));
NAND_g _29944_ (.A(_07941_), .B(_08625_), .Y(_08626_));
NAND_g _29945_ (.A(instr_rdcycleh), .B(count_cycle[59]), .Y(_08627_));
NAND_g _29946_ (.A(count_instr[59]), .B(instr_rdinstrh), .Y(_08628_));
AND_g _29947_ (.A(_08627_), .B(_08628_), .Y(_08629_));
NAND_g _29948_ (.A(count_instr[27]), .B(instr_rdinstr), .Y(_08630_));
NAND_g _29949_ (.A(instr_rdcycle), .B(count_cycle[27]), .Y(_08631_));
AND_g _29950_ (.A(_08630_), .B(_08631_), .Y(_08632_));
NAND_g _29951_ (.A(_08629_), .B(_08632_), .Y(_08633_));
NAND_g _29952_ (.A(_10595_), .B(_08633_), .Y(_08634_));
NAND_g _29953_ (.A(pcpi_rs1[27]), .B(_13889_), .Y(_08635_));
AND_g _29954_ (.A(_08634_), .B(_08635_), .Y(_08636_));
NOR_g _29955_ (.A(_14218_), .B(_08621_), .Y(_08637_));
NAND_g _29956_ (.A(_08622_), .B(_08637_), .Y(_08638_));
AND_g _29957_ (.A(_08636_), .B(_08638_), .Y(_08639_));
NAND_g _29958_ (.A(_08626_), .B(_08639_), .Y(_08640_));
AND_g _29959_ (.A(resetn), .B(_08640_), .Y(_00005_[27]));
NAND_g _29960_ (.A(reg_pc[28]), .B(decoded_imm[28]), .Y(_08641_));
XOR_g _29961_ (.A(reg_pc[28]), .B(decoded_imm[28]), .Y(_08642_));
AND_g _29962_ (.A(_08617_), .B(_08618_), .Y(_08643_));
NOR_g _29963_ (.A(_08619_), .B(_08643_), .Y(_08644_));
NAND_g _29964_ (.A(_08642_), .B(_08644_), .Y(_08645_));
NOR_g _29965_ (.A(_08642_), .B(_08644_), .Y(_08646_));
NOR_g _29966_ (.A(_14215_), .B(_08646_), .Y(_08647_));
NAND_g _29967_ (.A(_08645_), .B(_08647_), .Y(_08648_));
AND_g _29968_ (.A(latched_is_lu), .B(mem_rdata[28]), .Y(_08649_));
NAND_g _29969_ (.A(_01700_), .B(_08649_), .Y(_08650_));
NAND_g _29970_ (.A(_08362_), .B(_08650_), .Y(_08651_));
NAND_g _29971_ (.A(_07941_), .B(_08651_), .Y(_08652_));
NAND_g _29972_ (.A(instr_rdcycleh), .B(count_cycle[60]), .Y(_08653_));
NAND_g _29973_ (.A(count_instr[60]), .B(instr_rdinstrh), .Y(_08654_));
AND_g _29974_ (.A(_08653_), .B(_08654_), .Y(_08655_));
NAND_g _29975_ (.A(count_instr[28]), .B(instr_rdinstr), .Y(_08656_));
NAND_g _29976_ (.A(instr_rdcycle), .B(count_cycle[28]), .Y(_08657_));
AND_g _29977_ (.A(_08656_), .B(_08657_), .Y(_08658_));
NAND_g _29978_ (.A(_08655_), .B(_08658_), .Y(_08659_));
NAND_g _29979_ (.A(_10595_), .B(_08659_), .Y(_08660_));
NAND_g _29980_ (.A(pcpi_rs1[28]), .B(_13889_), .Y(_08661_));
AND_g _29981_ (.A(_08660_), .B(_08661_), .Y(_08662_));
AND_g _29982_ (.A(_08652_), .B(_08662_), .Y(_08663_));
NAND_g _29983_ (.A(_08648_), .B(_08663_), .Y(_08664_));
AND_g _29984_ (.A(resetn), .B(_08664_), .Y(_00005_[28]));
AND_g _29985_ (.A(latched_is_lu), .B(mem_rdata[29]), .Y(_08665_));
NAND_g _29986_ (.A(_01700_), .B(_08665_), .Y(_08666_));
NAND_g _29987_ (.A(_08362_), .B(_08666_), .Y(_08667_));
NAND_g _29988_ (.A(_07941_), .B(_08667_), .Y(_08668_));
NAND_g _29989_ (.A(instr_rdcycleh), .B(count_cycle[61]), .Y(_08669_));
NAND_g _29990_ (.A(count_instr[61]), .B(instr_rdinstrh), .Y(_08670_));
AND_g _29991_ (.A(_08669_), .B(_08670_), .Y(_08671_));
NAND_g _29992_ (.A(count_instr[29]), .B(instr_rdinstr), .Y(_08672_));
NAND_g _29993_ (.A(instr_rdcycle), .B(count_cycle[29]), .Y(_08673_));
AND_g _29994_ (.A(_08672_), .B(_08673_), .Y(_08674_));
NAND_g _29995_ (.A(_08671_), .B(_08674_), .Y(_08675_));
NAND_g _29996_ (.A(_10595_), .B(_08675_), .Y(_08676_));
NAND_g _29997_ (.A(pcpi_rs1[29]), .B(_13889_), .Y(_08677_));
AND_g _29998_ (.A(_08676_), .B(_08677_), .Y(_08678_));
AND_g _29999_ (.A(_08668_), .B(_08678_), .Y(_08679_));
NAND_g _30000_ (.A(_08641_), .B(_08645_), .Y(_08680_));
NAND_g _30001_ (.A(reg_pc[29]), .B(decoded_imm[29]), .Y(_08681_));
XOR_g _30002_ (.A(reg_pc[29]), .B(decoded_imm[29]), .Y(_08682_));
NAND_g _30003_ (.A(_08680_), .B(_08682_), .Y(_08683_));
XOR_g _30004_ (.A(_08680_), .B(_08682_), .Y(_08684_));
NAND_g _30005_ (.A(_14217_), .B(_08684_), .Y(_08685_));
NAND_g _30006_ (.A(_08679_), .B(_08685_), .Y(_08686_));
AND_g _30007_ (.A(resetn), .B(_08686_), .Y(_00005_[29]));
NAND_g _30008_ (.A(_08681_), .B(_08683_), .Y(_08687_));
NAND_g _30009_ (.A(reg_pc[30]), .B(decoded_imm[30]), .Y(_08688_));
XOR_g _30010_ (.A(reg_pc[30]), .B(decoded_imm[30]), .Y(_08689_));
NAND_g _30011_ (.A(_08687_), .B(_08689_), .Y(_08690_));
AND_g _30012_ (.A(latched_is_lu), .B(mem_rdata[30]), .Y(_08691_));
NAND_g _30013_ (.A(_01700_), .B(_08691_), .Y(_08692_));
NAND_g _30014_ (.A(_08362_), .B(_08692_), .Y(_08693_));
NAND_g _30015_ (.A(_07941_), .B(_08693_), .Y(_08694_));
NAND_g _30016_ (.A(instr_rdcycleh), .B(count_cycle[62]), .Y(_08695_));
NAND_g _30017_ (.A(count_instr[62]), .B(instr_rdinstrh), .Y(_08696_));
AND_g _30018_ (.A(_08695_), .B(_08696_), .Y(_08697_));
NAND_g _30019_ (.A(count_instr[30]), .B(instr_rdinstr), .Y(_08698_));
NAND_g _30020_ (.A(instr_rdcycle), .B(count_cycle[30]), .Y(_08699_));
AND_g _30021_ (.A(_08698_), .B(_08699_), .Y(_08700_));
NAND_g _30022_ (.A(_08697_), .B(_08700_), .Y(_08701_));
NAND_g _30023_ (.A(_10595_), .B(_08701_), .Y(_08702_));
NAND_g _30024_ (.A(pcpi_rs1[30]), .B(_13889_), .Y(_08703_));
AND_g _30025_ (.A(_08702_), .B(_08703_), .Y(_08704_));
XOR_g _30026_ (.A(_08687_), .B(_08689_), .Y(_08705_));
NAND_g _30027_ (.A(_14217_), .B(_08705_), .Y(_08706_));
AND_g _30028_ (.A(_08704_), .B(_08706_), .Y(_08707_));
NAND_g _30029_ (.A(_08694_), .B(_08707_), .Y(_08708_));
AND_g _30030_ (.A(resetn), .B(_08708_), .Y(_00005_[30]));
AND_g _30031_ (.A(_08688_), .B(_08690_), .Y(_08709_));
NAND_g _30032_ (.A(_08688_), .B(_08690_), .Y(_08710_));
XNOR_g _30033_ (.A(reg_pc[31]), .B(decoded_imm[31]), .Y(_08711_));
XOR_g _30034_ (.A(reg_pc[31]), .B(decoded_imm[31]), .Y(_08712_));
NAND_g _30035_ (.A(_08710_), .B(_08712_), .Y(_08713_));
NAND_g _30036_ (.A(_08709_), .B(_08711_), .Y(_08714_));
AND_g _30037_ (.A(_14214_), .B(_08714_), .Y(_08715_));
NAND_g _30038_ (.A(_08713_), .B(_08715_), .Y(_08716_));
AND_g _30039_ (.A(latched_is_lu), .B(mem_rdata[31]), .Y(_08717_));
NAND_g _30040_ (.A(_01700_), .B(_08717_), .Y(_08718_));
NAND_g _30041_ (.A(_08362_), .B(_08718_), .Y(_08719_));
NAND_g _30042_ (.A(_07941_), .B(_08719_), .Y(_08720_));
NAND_g _30043_ (.A(instr_rdcycleh), .B(count_cycle[63]), .Y(_08721_));
NAND_g _30044_ (.A(count_instr[63]), .B(instr_rdinstrh), .Y(_08722_));
AND_g _30045_ (.A(_08721_), .B(_08722_), .Y(_08723_));
NAND_g _30046_ (.A(count_instr[31]), .B(instr_rdinstr), .Y(_08724_));
NAND_g _30047_ (.A(instr_rdcycle), .B(count_cycle[31]), .Y(_08725_));
AND_g _30048_ (.A(_08724_), .B(_08725_), .Y(_08726_));
NAND_g _30049_ (.A(_08723_), .B(_08726_), .Y(_08727_));
NAND_g _30050_ (.A(_10595_), .B(_08727_), .Y(_08728_));
NAND_g _30051_ (.A(pcpi_rs1[31]), .B(_13889_), .Y(_08729_));
AND_g _30052_ (.A(_08728_), .B(_08729_), .Y(_08730_));
AND_g _30053_ (.A(_08720_), .B(_08730_), .Y(_08731_));
NAND_g _30054_ (.A(_08716_), .B(_08731_), .Y(_08732_));
AND_g _30055_ (.A(resetn), .B(_08732_), .Y(_00005_[31]));
XNOR_g _30056_ (.A(_09021_), .B(_13879_), .Y(_08733_));
NAND_g _30057_ (.A(_13883_), .B(_08733_), .Y(_08734_));
NAND_g _30058_ (.A(decoded_imm_j[11]), .B(_02997_), .Y(_08735_));
AND_g _30059_ (.A(_08734_), .B(_08735_), .Y(_08736_));
NAND_g _30060_ (.A(_10757_), .B(_08736_), .Y(_08737_));
AND_g _30061_ (.A(resetn), .B(_08737_), .Y(_00006_[0]));
NAND_g _30062_ (.A(decoded_imm_j[1]), .B(_02997_), .Y(_08738_));
AND_g _30063_ (.A(reg_sh[1]), .B(_13881_), .Y(_08739_));
NAND_g _30064_ (.A(_13876_), .B(_08739_), .Y(_08740_));
AND_g _30065_ (.A(_08738_), .B(_08740_), .Y(_08741_));
NAND_g _30066_ (.A(_10858_), .B(_08741_), .Y(_08742_));
AND_g _30067_ (.A(resetn), .B(_08742_), .Y(_00006_[1]));
NAND_g _30068_ (.A(decoded_imm_j[2]), .B(_02997_), .Y(_08743_));
NOR_g _30069_ (.A(reg_sh[2]), .B(_13879_), .Y(_08744_));
NAND_g _30070_ (.A(_13876_), .B(_08744_), .Y(_08745_));
AND_g _30071_ (.A(_08743_), .B(_08745_), .Y(_08746_));
NAND_g _30072_ (.A(_10960_), .B(_08746_), .Y(_08747_));
AND_g _30073_ (.A(resetn), .B(_08747_), .Y(_00006_[2]));
NAND_g _30074_ (.A(reg_sh[3]), .B(reg_sh[2]), .Y(_08748_));
NAND_g _30075_ (.A(reg_sh[4]), .B(_13878_), .Y(_08749_));
NAND_g _30076_ (.A(_08748_), .B(_08749_), .Y(_08750_));
NAND_g _30077_ (.A(_13876_), .B(_08750_), .Y(_08751_));
NAND_g _30078_ (.A(decoded_imm_j[3]), .B(_02997_), .Y(_08752_));
AND_g _30079_ (.A(_08751_), .B(_08752_), .Y(_08753_));
AND_g _30080_ (.A(_11060_), .B(_08753_), .Y(_08754_));
NAND_g _30081_ (.A(_11059_), .B(_08754_), .Y(_08755_));
AND_g _30082_ (.A(resetn), .B(_08755_), .Y(_00006_[3]));
NAND_g _30083_ (.A(decoded_imm_j[4]), .B(_02997_), .Y(_08756_));
NOR_g _30084_ (.A(_09022_), .B(_13878_), .Y(_08757_));
NAND_g _30085_ (.A(_13876_), .B(_08757_), .Y(_08758_));
AND_g _30086_ (.A(_08756_), .B(_08758_), .Y(_08759_));
NAND_g _30087_ (.A(_11164_), .B(_08759_), .Y(_08760_));
AND_g _30088_ (.A(resetn), .B(_08760_), .Y(_00006_[4]));
BUF_g _30089_ (.A(cpuregs[0][0]), .Y(_01113_));
BUF_g _30090_ (.A(cpuregs[0][1]), .Y(_01114_));
BUF_g _30091_ (.A(cpuregs[0][2]), .Y(_01115_));
BUF_g _30092_ (.A(cpuregs[0][3]), .Y(_01116_));
BUF_g _30093_ (.A(cpuregs[0][4]), .Y(_01117_));
BUF_g _30094_ (.A(cpuregs[0][5]), .Y(_01118_));
BUF_g _30095_ (.A(cpuregs[0][6]), .Y(_01119_));
BUF_g _30096_ (.A(cpuregs[0][7]), .Y(_01120_));
BUF_g _30097_ (.A(cpuregs[0][8]), .Y(_01121_));
BUF_g _30098_ (.A(cpuregs[0][9]), .Y(_01122_));
BUF_g _30099_ (.A(cpuregs[0][10]), .Y(_01123_));
BUF_g _30100_ (.A(cpuregs[0][11]), .Y(_01124_));
BUF_g _30101_ (.A(cpuregs[0][12]), .Y(_01125_));
BUF_g _30102_ (.A(cpuregs[0][13]), .Y(_01126_));
BUF_g _30103_ (.A(cpuregs[0][14]), .Y(_01127_));
BUF_g _30104_ (.A(cpuregs[0][15]), .Y(_01128_));
BUF_g _30105_ (.A(cpuregs[0][16]), .Y(_01129_));
BUF_g _30106_ (.A(cpuregs[0][17]), .Y(_01130_));
BUF_g _30107_ (.A(cpuregs[0][18]), .Y(_01131_));
BUF_g _30108_ (.A(cpuregs[0][19]), .Y(_01132_));
BUF_g _30109_ (.A(cpuregs[0][20]), .Y(_01133_));
BUF_g _30110_ (.A(cpuregs[0][21]), .Y(_01134_));
BUF_g _30111_ (.A(cpuregs[0][22]), .Y(_01135_));
BUF_g _30112_ (.A(cpuregs[0][23]), .Y(_01136_));
BUF_g _30113_ (.A(cpuregs[0][24]), .Y(_01137_));
BUF_g _30114_ (.A(cpuregs[0][25]), .Y(_01138_));
BUF_g _30115_ (.A(cpuregs[0][26]), .Y(_01139_));
BUF_g _30116_ (.A(cpuregs[0][27]), .Y(_01140_));
BUF_g _30117_ (.A(cpuregs[0][28]), .Y(_01141_));
BUF_g _30118_ (.A(cpuregs[0][29]), .Y(_01142_));
BUF_g _30119_ (.A(cpuregs[0][30]), .Y(_01143_));
BUF_g _30120_ (.A(cpuregs[0][31]), .Y(_01144_));
NAND_g _30121_ (.A(_14848_), .B(_14849_), .Y(_00009_));
NAND_g _30122_ (.A(_14852_), .B(_14853_), .Y(_00010_));
NAND_g _30123_ (.A(_14856_), .B(_14857_), .Y(_00011_));
NAND_g _30124_ (.A(_14860_), .B(_14861_), .Y(_00012_));
NAND_g _30125_ (.A(_02030_), .B(_02031_), .Y(_00013_));
NAND_g _30126_ (.A(_02964_), .B(_02965_), .Y(_00014_));
NAND_g _30127_ (.A(_02966_), .B(_02967_), .Y(_00015_));
NAND_g _30128_ (.A(_02968_), .B(_02969_), .Y(_00016_));
NAND_g _30129_ (.A(_02970_), .B(_02971_), .Y(_00017_));
NAND_g _30130_ (.A(_02972_), .B(_02973_), .Y(_00018_));
DFFcell _30131_ (.C(clk), .D(_00019_), .Q(cpuregs[15][0]));
DFFcell _30132_ (.C(clk), .D(_00020_), .Q(cpuregs[15][1]));
DFFcell _30133_ (.C(clk), .D(_00021_), .Q(cpuregs[15][2]));
DFFcell _30134_ (.C(clk), .D(_00022_), .Q(cpuregs[15][3]));
DFFcell _30135_ (.C(clk), .D(_00023_), .Q(cpuregs[15][4]));
DFFcell _30136_ (.C(clk), .D(_00024_), .Q(cpuregs[15][5]));
DFFcell _30137_ (.C(clk), .D(_00025_), .Q(cpuregs[15][6]));
DFFcell _30138_ (.C(clk), .D(_00026_), .Q(cpuregs[15][7]));
DFFcell _30139_ (.C(clk), .D(_00027_), .Q(cpuregs[15][8]));
DFFcell _30140_ (.C(clk), .D(_00028_), .Q(cpuregs[15][9]));
DFFcell _30141_ (.C(clk), .D(_00029_), .Q(cpuregs[15][10]));
DFFcell _30142_ (.C(clk), .D(_00030_), .Q(cpuregs[15][11]));
DFFcell _30143_ (.C(clk), .D(_00031_), .Q(cpuregs[15][12]));
DFFcell _30144_ (.C(clk), .D(_00032_), .Q(cpuregs[15][13]));
DFFcell _30145_ (.C(clk), .D(_00033_), .Q(cpuregs[15][14]));
DFFcell _30146_ (.C(clk), .D(_00034_), .Q(cpuregs[15][15]));
DFFcell _30147_ (.C(clk), .D(_00035_), .Q(cpuregs[15][16]));
DFFcell _30148_ (.C(clk), .D(_00036_), .Q(cpuregs[15][17]));
DFFcell _30149_ (.C(clk), .D(_00037_), .Q(cpuregs[15][18]));
DFFcell _30150_ (.C(clk), .D(_00038_), .Q(cpuregs[15][19]));
DFFcell _30151_ (.C(clk), .D(_00039_), .Q(cpuregs[15][20]));
DFFcell _30152_ (.C(clk), .D(_00040_), .Q(cpuregs[15][21]));
DFFcell _30153_ (.C(clk), .D(_00041_), .Q(cpuregs[15][22]));
DFFcell _30154_ (.C(clk), .D(_00042_), .Q(cpuregs[15][23]));
DFFcell _30155_ (.C(clk), .D(_00043_), .Q(cpuregs[15][24]));
DFFcell _30156_ (.C(clk), .D(_00044_), .Q(cpuregs[15][25]));
DFFcell _30157_ (.C(clk), .D(_00045_), .Q(cpuregs[15][26]));
DFFcell _30158_ (.C(clk), .D(_00046_), .Q(cpuregs[15][27]));
DFFcell _30159_ (.C(clk), .D(_00047_), .Q(cpuregs[15][28]));
DFFcell _30160_ (.C(clk), .D(_00048_), .Q(cpuregs[15][29]));
DFFcell _30161_ (.C(clk), .D(_00049_), .Q(cpuregs[15][30]));
DFFcell _30162_ (.C(clk), .D(_00050_), .Q(cpuregs[15][31]));
DFFcell _30163_ (.C(clk), .D(_00009_), .Q(_00007_[0]));
DFFcell _30164_ (.C(clk), .D(_00010_), .Q(_00007_[1]));
DFFcell _30165_ (.C(clk), .D(_00011_), .Q(_00007_[2]));
DFFcell _30166_ (.C(clk), .D(_00012_), .Q(_00007_[3]));
DFFcell _30167_ (.C(clk), .D(_00013_), .Q(_00007_[4]));
DFFcell _30168_ (.C(clk), .D(_00051_), .Q(cpuregs[30][0]));
DFFcell _30169_ (.C(clk), .D(_00052_), .Q(cpuregs[30][1]));
DFFcell _30170_ (.C(clk), .D(_00053_), .Q(cpuregs[30][2]));
DFFcell _30171_ (.C(clk), .D(_00054_), .Q(cpuregs[30][3]));
DFFcell _30172_ (.C(clk), .D(_00055_), .Q(cpuregs[30][4]));
DFFcell _30173_ (.C(clk), .D(_00056_), .Q(cpuregs[30][5]));
DFFcell _30174_ (.C(clk), .D(_00057_), .Q(cpuregs[30][6]));
DFFcell _30175_ (.C(clk), .D(_00058_), .Q(cpuregs[30][7]));
DFFcell _30176_ (.C(clk), .D(_00059_), .Q(cpuregs[30][8]));
DFFcell _30177_ (.C(clk), .D(_00060_), .Q(cpuregs[30][9]));
DFFcell _30178_ (.C(clk), .D(_00061_), .Q(cpuregs[30][10]));
DFFcell _30179_ (.C(clk), .D(_00062_), .Q(cpuregs[30][11]));
DFFcell _30180_ (.C(clk), .D(_00063_), .Q(cpuregs[30][12]));
DFFcell _30181_ (.C(clk), .D(_00064_), .Q(cpuregs[30][13]));
DFFcell _30182_ (.C(clk), .D(_00065_), .Q(cpuregs[30][14]));
DFFcell _30183_ (.C(clk), .D(_00066_), .Q(cpuregs[30][15]));
DFFcell _30184_ (.C(clk), .D(_00067_), .Q(cpuregs[30][16]));
DFFcell _30185_ (.C(clk), .D(_00068_), .Q(cpuregs[30][17]));
DFFcell _30186_ (.C(clk), .D(_00069_), .Q(cpuregs[30][18]));
DFFcell _30187_ (.C(clk), .D(_00070_), .Q(cpuregs[30][19]));
DFFcell _30188_ (.C(clk), .D(_00071_), .Q(cpuregs[30][20]));
DFFcell _30189_ (.C(clk), .D(_00072_), .Q(cpuregs[30][21]));
DFFcell _30190_ (.C(clk), .D(_00073_), .Q(cpuregs[30][22]));
DFFcell _30191_ (.C(clk), .D(_00074_), .Q(cpuregs[30][23]));
DFFcell _30192_ (.C(clk), .D(_00075_), .Q(cpuregs[30][24]));
DFFcell _30193_ (.C(clk), .D(_00076_), .Q(cpuregs[30][25]));
DFFcell _30194_ (.C(clk), .D(_00077_), .Q(cpuregs[30][26]));
DFFcell _30195_ (.C(clk), .D(_00078_), .Q(cpuregs[30][27]));
DFFcell _30196_ (.C(clk), .D(_00079_), .Q(cpuregs[30][28]));
DFFcell _30197_ (.C(clk), .D(_00080_), .Q(cpuregs[30][29]));
DFFcell _30198_ (.C(clk), .D(_00081_), .Q(cpuregs[30][30]));
DFFcell _30199_ (.C(clk), .D(_00082_), .Q(cpuregs[30][31]));
DFFcell _30200_ (.C(clk), .D(_00083_), .Q(cpuregs[2][0]));
DFFcell _30201_ (.C(clk), .D(_00084_), .Q(cpuregs[2][1]));
DFFcell _30202_ (.C(clk), .D(_00085_), .Q(cpuregs[2][2]));
DFFcell _30203_ (.C(clk), .D(_00086_), .Q(cpuregs[2][3]));
DFFcell _30204_ (.C(clk), .D(_00087_), .Q(cpuregs[2][4]));
DFFcell _30205_ (.C(clk), .D(_00088_), .Q(cpuregs[2][5]));
DFFcell _30206_ (.C(clk), .D(_00089_), .Q(cpuregs[2][6]));
DFFcell _30207_ (.C(clk), .D(_00090_), .Q(cpuregs[2][7]));
DFFcell _30208_ (.C(clk), .D(_00091_), .Q(cpuregs[2][8]));
DFFcell _30209_ (.C(clk), .D(_00092_), .Q(cpuregs[2][9]));
DFFcell _30210_ (.C(clk), .D(_00093_), .Q(cpuregs[2][10]));
DFFcell _30211_ (.C(clk), .D(_00094_), .Q(cpuregs[2][11]));
DFFcell _30212_ (.C(clk), .D(_00095_), .Q(cpuregs[2][12]));
DFFcell _30213_ (.C(clk), .D(_00096_), .Q(cpuregs[2][13]));
DFFcell _30214_ (.C(clk), .D(_00097_), .Q(cpuregs[2][14]));
DFFcell _30215_ (.C(clk), .D(_00098_), .Q(cpuregs[2][15]));
DFFcell _30216_ (.C(clk), .D(_00099_), .Q(cpuregs[2][16]));
DFFcell _30217_ (.C(clk), .D(_00100_), .Q(cpuregs[2][17]));
DFFcell _30218_ (.C(clk), .D(_00101_), .Q(cpuregs[2][18]));
DFFcell _30219_ (.C(clk), .D(_00102_), .Q(cpuregs[2][19]));
DFFcell _30220_ (.C(clk), .D(_00103_), .Q(cpuregs[2][20]));
DFFcell _30221_ (.C(clk), .D(_00104_), .Q(cpuregs[2][21]));
DFFcell _30222_ (.C(clk), .D(_00105_), .Q(cpuregs[2][22]));
DFFcell _30223_ (.C(clk), .D(_00106_), .Q(cpuregs[2][23]));
DFFcell _30224_ (.C(clk), .D(_00107_), .Q(cpuregs[2][24]));
DFFcell _30225_ (.C(clk), .D(_00108_), .Q(cpuregs[2][25]));
DFFcell _30226_ (.C(clk), .D(_00109_), .Q(cpuregs[2][26]));
DFFcell _30227_ (.C(clk), .D(_00110_), .Q(cpuregs[2][27]));
DFFcell _30228_ (.C(clk), .D(_00111_), .Q(cpuregs[2][28]));
DFFcell _30229_ (.C(clk), .D(_00112_), .Q(cpuregs[2][29]));
DFFcell _30230_ (.C(clk), .D(_00113_), .Q(cpuregs[2][30]));
DFFcell _30231_ (.C(clk), .D(_00114_), .Q(cpuregs[2][31]));
DFFcell _30232_ (.C(clk), .D(_00115_), .Q(count_cycle[0]));
DFFcell _30233_ (.C(clk), .D(_00116_), .Q(count_cycle[1]));
DFFcell _30234_ (.C(clk), .D(_00117_), .Q(count_cycle[2]));
DFFcell _30235_ (.C(clk), .D(_00118_), .Q(count_cycle[3]));
DFFcell _30236_ (.C(clk), .D(_00119_), .Q(count_cycle[4]));
DFFcell _30237_ (.C(clk), .D(_00120_), .Q(count_cycle[5]));
DFFcell _30238_ (.C(clk), .D(_00121_), .Q(count_cycle[6]));
DFFcell _30239_ (.C(clk), .D(_00122_), .Q(count_cycle[7]));
DFFcell _30240_ (.C(clk), .D(_00123_), .Q(count_cycle[8]));
DFFcell _30241_ (.C(clk), .D(_00124_), .Q(count_cycle[9]));
DFFcell _30242_ (.C(clk), .D(_00125_), .Q(count_cycle[10]));
DFFcell _30243_ (.C(clk), .D(_00126_), .Q(count_cycle[11]));
DFFcell _30244_ (.C(clk), .D(_00127_), .Q(count_cycle[12]));
DFFcell _30245_ (.C(clk), .D(_00128_), .Q(count_cycle[13]));
DFFcell _30246_ (.C(clk), .D(_00129_), .Q(count_cycle[14]));
DFFcell _30247_ (.C(clk), .D(_00130_), .Q(count_cycle[15]));
DFFcell _30248_ (.C(clk), .D(_00131_), .Q(count_cycle[16]));
DFFcell _30249_ (.C(clk), .D(_00132_), .Q(count_cycle[17]));
DFFcell _30250_ (.C(clk), .D(_00133_), .Q(count_cycle[18]));
DFFcell _30251_ (.C(clk), .D(_00134_), .Q(count_cycle[19]));
DFFcell _30252_ (.C(clk), .D(_00135_), .Q(count_cycle[20]));
DFFcell _30253_ (.C(clk), .D(_00136_), .Q(count_cycle[21]));
DFFcell _30254_ (.C(clk), .D(_00137_), .Q(count_cycle[22]));
DFFcell _30255_ (.C(clk), .D(_00138_), .Q(count_cycle[23]));
DFFcell _30256_ (.C(clk), .D(_00139_), .Q(count_cycle[24]));
DFFcell _30257_ (.C(clk), .D(_00140_), .Q(count_cycle[25]));
DFFcell _30258_ (.C(clk), .D(_00141_), .Q(count_cycle[26]));
DFFcell _30259_ (.C(clk), .D(_00142_), .Q(count_cycle[27]));
DFFcell _30260_ (.C(clk), .D(_00143_), .Q(count_cycle[28]));
DFFcell _30261_ (.C(clk), .D(_00144_), .Q(count_cycle[29]));
DFFcell _30262_ (.C(clk), .D(_00145_), .Q(count_cycle[30]));
DFFcell _30263_ (.C(clk), .D(_00146_), .Q(count_cycle[31]));
DFFcell _30264_ (.C(clk), .D(_00147_), .Q(count_cycle[32]));
DFFcell _30265_ (.C(clk), .D(_00148_), .Q(count_cycle[33]));
DFFcell _30266_ (.C(clk), .D(_00149_), .Q(count_cycle[34]));
DFFcell _30267_ (.C(clk), .D(_00150_), .Q(count_cycle[35]));
DFFcell _30268_ (.C(clk), .D(_00151_), .Q(count_cycle[36]));
DFFcell _30269_ (.C(clk), .D(_00152_), .Q(count_cycle[37]));
DFFcell _30270_ (.C(clk), .D(_00153_), .Q(count_cycle[38]));
DFFcell _30271_ (.C(clk), .D(_00154_), .Q(count_cycle[39]));
DFFcell _30272_ (.C(clk), .D(_00155_), .Q(count_cycle[40]));
DFFcell _30273_ (.C(clk), .D(_00156_), .Q(count_cycle[41]));
DFFcell _30274_ (.C(clk), .D(_00157_), .Q(count_cycle[42]));
DFFcell _30275_ (.C(clk), .D(_00158_), .Q(count_cycle[43]));
DFFcell _30276_ (.C(clk), .D(_00159_), .Q(count_cycle[44]));
DFFcell _30277_ (.C(clk), .D(_00160_), .Q(count_cycle[45]));
DFFcell _30278_ (.C(clk), .D(_00161_), .Q(count_cycle[46]));
DFFcell _30279_ (.C(clk), .D(_00162_), .Q(count_cycle[47]));
DFFcell _30280_ (.C(clk), .D(_00163_), .Q(count_cycle[48]));
DFFcell _30281_ (.C(clk), .D(_00164_), .Q(count_cycle[49]));
DFFcell _30282_ (.C(clk), .D(_00165_), .Q(count_cycle[50]));
DFFcell _30283_ (.C(clk), .D(_00166_), .Q(count_cycle[51]));
DFFcell _30284_ (.C(clk), .D(_00167_), .Q(count_cycle[52]));
DFFcell _30285_ (.C(clk), .D(_00168_), .Q(count_cycle[53]));
DFFcell _30286_ (.C(clk), .D(_00169_), .Q(count_cycle[54]));
DFFcell _30287_ (.C(clk), .D(_00170_), .Q(count_cycle[55]));
DFFcell _30288_ (.C(clk), .D(_00171_), .Q(count_cycle[56]));
DFFcell _30289_ (.C(clk), .D(_00172_), .Q(count_cycle[57]));
DFFcell _30290_ (.C(clk), .D(_00173_), .Q(count_cycle[58]));
DFFcell _30291_ (.C(clk), .D(_00174_), .Q(count_cycle[59]));
DFFcell _30292_ (.C(clk), .D(_00175_), .Q(count_cycle[60]));
DFFcell _30293_ (.C(clk), .D(_00176_), .Q(count_cycle[61]));
DFFcell _30294_ (.C(clk), .D(_00177_), .Q(count_cycle[62]));
DFFcell _30295_ (.C(clk), .D(_00178_), .Q(count_cycle[63]));
DFFcell _30296_ (.C(clk), .D(_00179_), .Q(trap));
DFFcell _30297_ (.C(clk), .D(_00180_), .Q(cpuregs[1][0]));
DFFcell _30298_ (.C(clk), .D(_00181_), .Q(cpuregs[1][1]));
DFFcell _30299_ (.C(clk), .D(_00182_), .Q(cpuregs[1][2]));
DFFcell _30300_ (.C(clk), .D(_00183_), .Q(cpuregs[1][3]));
DFFcell _30301_ (.C(clk), .D(_00184_), .Q(cpuregs[1][4]));
DFFcell _30302_ (.C(clk), .D(_00185_), .Q(cpuregs[1][5]));
DFFcell _30303_ (.C(clk), .D(_00186_), .Q(cpuregs[1][6]));
DFFcell _30304_ (.C(clk), .D(_00187_), .Q(cpuregs[1][7]));
DFFcell _30305_ (.C(clk), .D(_00188_), .Q(cpuregs[1][8]));
DFFcell _30306_ (.C(clk), .D(_00189_), .Q(cpuregs[1][9]));
DFFcell _30307_ (.C(clk), .D(_00190_), .Q(cpuregs[1][10]));
DFFcell _30308_ (.C(clk), .D(_00191_), .Q(cpuregs[1][11]));
DFFcell _30309_ (.C(clk), .D(_00192_), .Q(cpuregs[1][12]));
DFFcell _30310_ (.C(clk), .D(_00193_), .Q(cpuregs[1][13]));
DFFcell _30311_ (.C(clk), .D(_00194_), .Q(cpuregs[1][14]));
DFFcell _30312_ (.C(clk), .D(_00195_), .Q(cpuregs[1][15]));
DFFcell _30313_ (.C(clk), .D(_00196_), .Q(cpuregs[1][16]));
DFFcell _30314_ (.C(clk), .D(_00197_), .Q(cpuregs[1][17]));
DFFcell _30315_ (.C(clk), .D(_00198_), .Q(cpuregs[1][18]));
DFFcell _30316_ (.C(clk), .D(_00199_), .Q(cpuregs[1][19]));
DFFcell _30317_ (.C(clk), .D(_00200_), .Q(cpuregs[1][20]));
DFFcell _30318_ (.C(clk), .D(_00201_), .Q(cpuregs[1][21]));
DFFcell _30319_ (.C(clk), .D(_00202_), .Q(cpuregs[1][22]));
DFFcell _30320_ (.C(clk), .D(_00203_), .Q(cpuregs[1][23]));
DFFcell _30321_ (.C(clk), .D(_00204_), .Q(cpuregs[1][24]));
DFFcell _30322_ (.C(clk), .D(_00205_), .Q(cpuregs[1][25]));
DFFcell _30323_ (.C(clk), .D(_00206_), .Q(cpuregs[1][26]));
DFFcell _30324_ (.C(clk), .D(_00207_), .Q(cpuregs[1][27]));
DFFcell _30325_ (.C(clk), .D(_00208_), .Q(cpuregs[1][28]));
DFFcell _30326_ (.C(clk), .D(_00209_), .Q(cpuregs[1][29]));
DFFcell _30327_ (.C(clk), .D(_00210_), .Q(cpuregs[1][30]));
DFFcell _30328_ (.C(clk), .D(_00211_), .Q(cpuregs[1][31]));
DFFcell _30329_ (.C(clk), .D(_00212_), .Q(mem_do_prefetch));
DFFcell _30330_ (.C(clk), .D(_00213_), .Q(reg_pc[1]));
DFFcell _30331_ (.C(clk), .D(_00214_), .Q(reg_pc[2]));
DFFcell _30332_ (.C(clk), .D(_00215_), .Q(reg_pc[3]));
DFFcell _30333_ (.C(clk), .D(_00216_), .Q(reg_pc[4]));
DFFcell _30334_ (.C(clk), .D(_00217_), .Q(reg_pc[5]));
DFFcell _30335_ (.C(clk), .D(_00218_), .Q(reg_pc[6]));
DFFcell _30336_ (.C(clk), .D(_00219_), .Q(reg_pc[7]));
DFFcell _30337_ (.C(clk), .D(_00220_), .Q(reg_pc[8]));
DFFcell _30338_ (.C(clk), .D(_00221_), .Q(reg_pc[9]));
DFFcell _30339_ (.C(clk), .D(_00222_), .Q(reg_pc[10]));
DFFcell _30340_ (.C(clk), .D(_00223_), .Q(reg_pc[11]));
DFFcell _30341_ (.C(clk), .D(_00224_), .Q(reg_pc[12]));
DFFcell _30342_ (.C(clk), .D(_00225_), .Q(reg_pc[13]));
DFFcell _30343_ (.C(clk), .D(_00226_), .Q(reg_pc[14]));
DFFcell _30344_ (.C(clk), .D(_00227_), .Q(reg_pc[15]));
DFFcell _30345_ (.C(clk), .D(_00228_), .Q(reg_pc[16]));
DFFcell _30346_ (.C(clk), .D(_00229_), .Q(reg_pc[17]));
DFFcell _30347_ (.C(clk), .D(_00230_), .Q(reg_pc[18]));
DFFcell _30348_ (.C(clk), .D(_00231_), .Q(reg_pc[19]));
DFFcell _30349_ (.C(clk), .D(_00232_), .Q(reg_pc[20]));
DFFcell _30350_ (.C(clk), .D(_00233_), .Q(reg_pc[21]));
DFFcell _30351_ (.C(clk), .D(_00234_), .Q(reg_pc[22]));
DFFcell _30352_ (.C(clk), .D(_00235_), .Q(reg_pc[23]));
DFFcell _30353_ (.C(clk), .D(_00236_), .Q(reg_pc[24]));
DFFcell _30354_ (.C(clk), .D(_00237_), .Q(reg_pc[25]));
DFFcell _30355_ (.C(clk), .D(_00238_), .Q(reg_pc[26]));
DFFcell _30356_ (.C(clk), .D(_00239_), .Q(reg_pc[27]));
DFFcell _30357_ (.C(clk), .D(_00240_), .Q(reg_pc[28]));
DFFcell _30358_ (.C(clk), .D(_00241_), .Q(reg_pc[29]));
DFFcell _30359_ (.C(clk), .D(_00242_), .Q(reg_pc[30]));
DFFcell _30360_ (.C(clk), .D(_00243_), .Q(reg_pc[31]));
DFFcell _30361_ (.C(clk), .D(_00244_), .Q(reg_next_pc[1]));
DFFcell _30362_ (.C(clk), .D(_00245_), .Q(reg_next_pc[2]));
DFFcell _30363_ (.C(clk), .D(_00246_), .Q(reg_next_pc[3]));
DFFcell _30364_ (.C(clk), .D(_00247_), .Q(reg_next_pc[4]));
DFFcell _30365_ (.C(clk), .D(_00248_), .Q(reg_next_pc[5]));
DFFcell _30366_ (.C(clk), .D(_00249_), .Q(reg_next_pc[6]));
DFFcell _30367_ (.C(clk), .D(_00250_), .Q(reg_next_pc[7]));
DFFcell _30368_ (.C(clk), .D(_00251_), .Q(reg_next_pc[8]));
DFFcell _30369_ (.C(clk), .D(_00252_), .Q(reg_next_pc[9]));
DFFcell _30370_ (.C(clk), .D(_00253_), .Q(reg_next_pc[10]));
DFFcell _30371_ (.C(clk), .D(_00254_), .Q(reg_next_pc[11]));
DFFcell _30372_ (.C(clk), .D(_00255_), .Q(reg_next_pc[12]));
DFFcell _30373_ (.C(clk), .D(_00256_), .Q(reg_next_pc[13]));
DFFcell _30374_ (.C(clk), .D(_00257_), .Q(reg_next_pc[14]));
DFFcell _30375_ (.C(clk), .D(_00258_), .Q(reg_next_pc[15]));
DFFcell _30376_ (.C(clk), .D(_00259_), .Q(reg_next_pc[16]));
DFFcell _30377_ (.C(clk), .D(_00260_), .Q(reg_next_pc[17]));
DFFcell _30378_ (.C(clk), .D(_00261_), .Q(reg_next_pc[18]));
DFFcell _30379_ (.C(clk), .D(_00262_), .Q(reg_next_pc[19]));
DFFcell _30380_ (.C(clk), .D(_00263_), .Q(reg_next_pc[20]));
DFFcell _30381_ (.C(clk), .D(_00264_), .Q(reg_next_pc[21]));
DFFcell _30382_ (.C(clk), .D(_00265_), .Q(reg_next_pc[22]));
DFFcell _30383_ (.C(clk), .D(_00266_), .Q(reg_next_pc[23]));
DFFcell _30384_ (.C(clk), .D(_00267_), .Q(reg_next_pc[24]));
DFFcell _30385_ (.C(clk), .D(_00268_), .Q(reg_next_pc[25]));
DFFcell _30386_ (.C(clk), .D(_00269_), .Q(reg_next_pc[26]));
DFFcell _30387_ (.C(clk), .D(_00270_), .Q(reg_next_pc[27]));
DFFcell _30388_ (.C(clk), .D(_00271_), .Q(reg_next_pc[28]));
DFFcell _30389_ (.C(clk), .D(_00272_), .Q(reg_next_pc[29]));
DFFcell _30390_ (.C(clk), .D(_00273_), .Q(reg_next_pc[30]));
DFFcell _30391_ (.C(clk), .D(_00274_), .Q(reg_next_pc[31]));
DFFcell _30392_ (.C(clk), .D(_00275_), .Q(pcpi_rs2[0]));
DFFcell _30393_ (.C(clk), .D(_00276_), .Q(pcpi_rs2[1]));
DFFcell _30394_ (.C(clk), .D(_00277_), .Q(pcpi_rs2[2]));
DFFcell _30395_ (.C(clk), .D(_00278_), .Q(pcpi_rs2[3]));
DFFcell _30396_ (.C(clk), .D(_00279_), .Q(pcpi_rs2[4]));
DFFcell _30397_ (.C(clk), .D(_00280_), .Q(pcpi_rs2[5]));
DFFcell _30398_ (.C(clk), .D(_00281_), .Q(pcpi_rs2[6]));
DFFcell _30399_ (.C(clk), .D(_00282_), .Q(pcpi_rs2[7]));
DFFcell _30400_ (.C(clk), .D(_00283_), .Q(pcpi_rs2[8]));
DFFcell _30401_ (.C(clk), .D(_00284_), .Q(pcpi_rs2[9]));
DFFcell _30402_ (.C(clk), .D(_00285_), .Q(pcpi_rs2[10]));
DFFcell _30403_ (.C(clk), .D(_00286_), .Q(pcpi_rs2[11]));
DFFcell _30404_ (.C(clk), .D(_00287_), .Q(pcpi_rs2[12]));
DFFcell _30405_ (.C(clk), .D(_00288_), .Q(pcpi_rs2[13]));
DFFcell _30406_ (.C(clk), .D(_00289_), .Q(pcpi_rs2[14]));
DFFcell _30407_ (.C(clk), .D(_00290_), .Q(pcpi_rs2[15]));
DFFcell _30408_ (.C(clk), .D(_00291_), .Q(pcpi_rs2[16]));
DFFcell _30409_ (.C(clk), .D(_00292_), .Q(pcpi_rs2[17]));
DFFcell _30410_ (.C(clk), .D(_00293_), .Q(pcpi_rs2[18]));
DFFcell _30411_ (.C(clk), .D(_00294_), .Q(pcpi_rs2[19]));
DFFcell _30412_ (.C(clk), .D(_00295_), .Q(pcpi_rs2[20]));
DFFcell _30413_ (.C(clk), .D(_00296_), .Q(pcpi_rs2[21]));
DFFcell _30414_ (.C(clk), .D(_00297_), .Q(pcpi_rs2[22]));
DFFcell _30415_ (.C(clk), .D(_00298_), .Q(pcpi_rs2[23]));
DFFcell _30416_ (.C(clk), .D(_00299_), .Q(pcpi_rs2[24]));
DFFcell _30417_ (.C(clk), .D(_00300_), .Q(pcpi_rs2[25]));
DFFcell _30418_ (.C(clk), .D(_00301_), .Q(pcpi_rs2[26]));
DFFcell _30419_ (.C(clk), .D(_00302_), .Q(pcpi_rs2[27]));
DFFcell _30420_ (.C(clk), .D(_00303_), .Q(pcpi_rs2[28]));
DFFcell _30421_ (.C(clk), .D(_00304_), .Q(pcpi_rs2[29]));
DFFcell _30422_ (.C(clk), .D(_00305_), .Q(pcpi_rs2[30]));
DFFcell _30423_ (.C(clk), .D(_00306_), .Q(pcpi_rs2[31]));
DFFcell _30424_ (.C(clk), .D(_00005_[0]), .Q(reg_out[0]));
DFFcell _30425_ (.C(clk), .D(_00005_[1]), .Q(reg_out[1]));
DFFcell _30426_ (.C(clk), .D(_00005_[2]), .Q(reg_out[2]));
DFFcell _30427_ (.C(clk), .D(_00005_[3]), .Q(reg_out[3]));
DFFcell _30428_ (.C(clk), .D(_00005_[4]), .Q(reg_out[4]));
DFFcell _30429_ (.C(clk), .D(_00005_[5]), .Q(reg_out[5]));
DFFcell _30430_ (.C(clk), .D(_00005_[6]), .Q(reg_out[6]));
DFFcell _30431_ (.C(clk), .D(_00005_[7]), .Q(reg_out[7]));
DFFcell _30432_ (.C(clk), .D(_00005_[8]), .Q(reg_out[8]));
DFFcell _30433_ (.C(clk), .D(_00005_[9]), .Q(reg_out[9]));
DFFcell _30434_ (.C(clk), .D(_00005_[10]), .Q(reg_out[10]));
DFFcell _30435_ (.C(clk), .D(_00005_[11]), .Q(reg_out[11]));
DFFcell _30436_ (.C(clk), .D(_00005_[12]), .Q(reg_out[12]));
DFFcell _30437_ (.C(clk), .D(_00005_[13]), .Q(reg_out[13]));
DFFcell _30438_ (.C(clk), .D(_00005_[14]), .Q(reg_out[14]));
DFFcell _30439_ (.C(clk), .D(_00005_[15]), .Q(reg_out[15]));
DFFcell _30440_ (.C(clk), .D(_00005_[16]), .Q(reg_out[16]));
DFFcell _30441_ (.C(clk), .D(_00005_[17]), .Q(reg_out[17]));
DFFcell _30442_ (.C(clk), .D(_00005_[18]), .Q(reg_out[18]));
DFFcell _30443_ (.C(clk), .D(_00005_[19]), .Q(reg_out[19]));
DFFcell _30444_ (.C(clk), .D(_00005_[20]), .Q(reg_out[20]));
DFFcell _30445_ (.C(clk), .D(_00005_[21]), .Q(reg_out[21]));
DFFcell _30446_ (.C(clk), .D(_00005_[22]), .Q(reg_out[22]));
DFFcell _30447_ (.C(clk), .D(_00005_[23]), .Q(reg_out[23]));
DFFcell _30448_ (.C(clk), .D(_00005_[24]), .Q(reg_out[24]));
DFFcell _30449_ (.C(clk), .D(_00005_[25]), .Q(reg_out[25]));
DFFcell _30450_ (.C(clk), .D(_00005_[26]), .Q(reg_out[26]));
DFFcell _30451_ (.C(clk), .D(_00005_[27]), .Q(reg_out[27]));
DFFcell _30452_ (.C(clk), .D(_00005_[28]), .Q(reg_out[28]));
DFFcell _30453_ (.C(clk), .D(_00005_[29]), .Q(reg_out[29]));
DFFcell _30454_ (.C(clk), .D(_00005_[30]), .Q(reg_out[30]));
DFFcell _30455_ (.C(clk), .D(_00005_[31]), .Q(reg_out[31]));
DFFcell _30456_ (.C(clk), .D(_00006_[0]), .Q(reg_sh[0]));
DFFcell _30457_ (.C(clk), .D(_00006_[1]), .Q(reg_sh[1]));
DFFcell _30458_ (.C(clk), .D(_00006_[2]), .Q(reg_sh[2]));
DFFcell _30459_ (.C(clk), .D(_00006_[3]), .Q(reg_sh[3]));
DFFcell _30460_ (.C(clk), .D(_00006_[4]), .Q(reg_sh[4]));
DFFcell _30461_ (.C(clk), .D(_00307_), .Q(instr_sw));
DFFcell _30462_ (.C(clk), .D(_00308_), .Q(decoder_pseudo_trigger));
DFFcell _30463_ (.C(clk), .D(_00309_), .Q(mem_do_rinst));
DFFcell _30464_ (.C(clk), .D(_00310_), .Q(mem_do_rdata));
DFFcell _30465_ (.C(clk), .D(_00311_), .Q(mem_do_wdata));
DFFcell _30466_ (.C(clk), .D(_00000_), .Q(decoder_trigger));
DFFcell _30467_ (.C(clk), .D(_00312_), .Q(mem_wordsize[0]));
DFFcell _30468_ (.C(clk), .D(_00313_), .Q(mem_wordsize[1]));
DFFcell _30469_ (.C(clk), .D(_00314_), .Q(mem_valid));
DFFcell _30470_ (.C(clk), .D(_00315_), .Q(cpuregs[20][0]));
DFFcell _30471_ (.C(clk), .D(_00316_), .Q(cpuregs[20][1]));
DFFcell _30472_ (.C(clk), .D(_00317_), .Q(cpuregs[20][2]));
DFFcell _30473_ (.C(clk), .D(_00318_), .Q(cpuregs[20][3]));
DFFcell _30474_ (.C(clk), .D(_00319_), .Q(cpuregs[20][4]));
DFFcell _30475_ (.C(clk), .D(_00320_), .Q(cpuregs[20][5]));
DFFcell _30476_ (.C(clk), .D(_00321_), .Q(cpuregs[20][6]));
DFFcell _30477_ (.C(clk), .D(_00322_), .Q(cpuregs[20][7]));
DFFcell _30478_ (.C(clk), .D(_00323_), .Q(cpuregs[20][8]));
DFFcell _30479_ (.C(clk), .D(_00324_), .Q(cpuregs[20][9]));
DFFcell _30480_ (.C(clk), .D(_00325_), .Q(cpuregs[20][10]));
DFFcell _30481_ (.C(clk), .D(_00326_), .Q(cpuregs[20][11]));
DFFcell _30482_ (.C(clk), .D(_00327_), .Q(cpuregs[20][12]));
DFFcell _30483_ (.C(clk), .D(_00328_), .Q(cpuregs[20][13]));
DFFcell _30484_ (.C(clk), .D(_00329_), .Q(cpuregs[20][14]));
DFFcell _30485_ (.C(clk), .D(_00330_), .Q(cpuregs[20][15]));
DFFcell _30486_ (.C(clk), .D(_00331_), .Q(cpuregs[20][16]));
DFFcell _30487_ (.C(clk), .D(_00332_), .Q(cpuregs[20][17]));
DFFcell _30488_ (.C(clk), .D(_00333_), .Q(cpuregs[20][18]));
DFFcell _30489_ (.C(clk), .D(_00334_), .Q(cpuregs[20][19]));
DFFcell _30490_ (.C(clk), .D(_00335_), .Q(cpuregs[20][20]));
DFFcell _30491_ (.C(clk), .D(_00336_), .Q(cpuregs[20][21]));
DFFcell _30492_ (.C(clk), .D(_00337_), .Q(cpuregs[20][22]));
DFFcell _30493_ (.C(clk), .D(_00338_), .Q(cpuregs[20][23]));
DFFcell _30494_ (.C(clk), .D(_00339_), .Q(cpuregs[20][24]));
DFFcell _30495_ (.C(clk), .D(_00340_), .Q(cpuregs[20][25]));
DFFcell _30496_ (.C(clk), .D(_00341_), .Q(cpuregs[20][26]));
DFFcell _30497_ (.C(clk), .D(_00342_), .Q(cpuregs[20][27]));
DFFcell _30498_ (.C(clk), .D(_00343_), .Q(cpuregs[20][28]));
DFFcell _30499_ (.C(clk), .D(_00344_), .Q(cpuregs[20][29]));
DFFcell _30500_ (.C(clk), .D(_00345_), .Q(cpuregs[20][30]));
DFFcell _30501_ (.C(clk), .D(_00346_), .Q(cpuregs[20][31]));
DFFcell _30502_ (.C(clk), .D(_00347_), .Q(latched_store));
DFFcell _30503_ (.C(clk), .D(_00348_), .Q(latched_stalu));
DFFcell _30504_ (.C(clk), .D(_00349_), .Q(latched_branch));
DFFcell _30505_ (.C(clk), .D(_00350_), .Q(latched_is_lu));
DFFcell _30506_ (.C(clk), .D(_00351_), .Q(latched_is_lh));
DFFcell _30507_ (.C(clk), .D(_00352_), .Q(latched_is_lb));
DFFcell _30508_ (.C(clk), .D(_00353_), .Q(latched_rd[0]));
DFFcell _30509_ (.C(clk), .D(_00354_), .Q(latched_rd[1]));
DFFcell _30510_ (.C(clk), .D(_00355_), .Q(latched_rd[2]));
DFFcell _30511_ (.C(clk), .D(_00356_), .Q(latched_rd[3]));
DFFcell _30512_ (.C(clk), .D(_00357_), .Q(latched_rd[4]));
DFFcell _30513_ (.C(clk), .D(alu_out[0]), .Q(alu_out_q[0]));
DFFcell _30514_ (.C(clk), .D(alu_out[1]), .Q(alu_out_q[1]));
DFFcell _30515_ (.C(clk), .D(alu_out[2]), .Q(alu_out_q[2]));
DFFcell _30516_ (.C(clk), .D(alu_out[3]), .Q(alu_out_q[3]));
DFFcell _30517_ (.C(clk), .D(alu_out[4]), .Q(alu_out_q[4]));
DFFcell _30518_ (.C(clk), .D(alu_out[5]), .Q(alu_out_q[5]));
DFFcell _30519_ (.C(clk), .D(alu_out[6]), .Q(alu_out_q[6]));
DFFcell _30520_ (.C(clk), .D(alu_out[7]), .Q(alu_out_q[7]));
DFFcell _30521_ (.C(clk), .D(alu_out[8]), .Q(alu_out_q[8]));
DFFcell _30522_ (.C(clk), .D(alu_out[9]), .Q(alu_out_q[9]));
DFFcell _30523_ (.C(clk), .D(alu_out[10]), .Q(alu_out_q[10]));
DFFcell _30524_ (.C(clk), .D(alu_out[11]), .Q(alu_out_q[11]));
DFFcell _30525_ (.C(clk), .D(alu_out[12]), .Q(alu_out_q[12]));
DFFcell _30526_ (.C(clk), .D(alu_out[13]), .Q(alu_out_q[13]));
DFFcell _30527_ (.C(clk), .D(alu_out[14]), .Q(alu_out_q[14]));
DFFcell _30528_ (.C(clk), .D(alu_out[15]), .Q(alu_out_q[15]));
DFFcell _30529_ (.C(clk), .D(alu_out[16]), .Q(alu_out_q[16]));
DFFcell _30530_ (.C(clk), .D(alu_out[17]), .Q(alu_out_q[17]));
DFFcell _30531_ (.C(clk), .D(alu_out[18]), .Q(alu_out_q[18]));
DFFcell _30532_ (.C(clk), .D(alu_out[19]), .Q(alu_out_q[19]));
DFFcell _30533_ (.C(clk), .D(alu_out[20]), .Q(alu_out_q[20]));
DFFcell _30534_ (.C(clk), .D(alu_out[21]), .Q(alu_out_q[21]));
DFFcell _30535_ (.C(clk), .D(alu_out[22]), .Q(alu_out_q[22]));
DFFcell _30536_ (.C(clk), .D(alu_out[23]), .Q(alu_out_q[23]));
DFFcell _30537_ (.C(clk), .D(alu_out[24]), .Q(alu_out_q[24]));
DFFcell _30538_ (.C(clk), .D(alu_out[25]), .Q(alu_out_q[25]));
DFFcell _30539_ (.C(clk), .D(alu_out[26]), .Q(alu_out_q[26]));
DFFcell _30540_ (.C(clk), .D(alu_out[27]), .Q(alu_out_q[27]));
DFFcell _30541_ (.C(clk), .D(alu_out[28]), .Q(alu_out_q[28]));
DFFcell _30542_ (.C(clk), .D(alu_out[29]), .Q(alu_out_q[29]));
DFFcell _30543_ (.C(clk), .D(alu_out[30]), .Q(alu_out_q[30]));
DFFcell _30544_ (.C(clk), .D(alu_out[31]), .Q(alu_out_q[31]));
DFFcell _30545_ (.C(clk), .D(_00358_), .Q(instr_lui));
DFFcell _30546_ (.C(clk), .D(_00359_), .Q(instr_auipc));
DFFcell _30547_ (.C(clk), .D(_00360_), .Q(instr_jal));
DFFcell _30548_ (.C(clk), .D(_00361_), .Q(instr_beq));
DFFcell _30549_ (.C(clk), .D(_00362_), .Q(instr_bne));
DFFcell _30550_ (.C(clk), .D(_00363_), .Q(instr_blt));
DFFcell _30551_ (.C(clk), .D(_00364_), .Q(instr_bge));
DFFcell _30552_ (.C(clk), .D(_00365_), .Q(instr_bltu));
DFFcell _30553_ (.C(clk), .D(_00366_), .Q(instr_bgeu));
DFFcell _30554_ (.C(clk), .D(_00367_), .Q(instr_jalr));
DFFcell _30555_ (.C(clk), .D(_00368_), .Q(instr_lb));
DFFcell _30556_ (.C(clk), .D(_00369_), .Q(instr_lh));
DFFcell _30557_ (.C(clk), .D(_00370_), .Q(instr_lw));
DFFcell _30558_ (.C(clk), .D(_00371_), .Q(instr_lbu));
DFFcell _30559_ (.C(clk), .D(_00372_), .Q(instr_lhu));
DFFcell _30560_ (.C(clk), .D(_00373_), .Q(pcpi_rs1[31]));
DFFcell _30561_ (.C(clk), .D(_00374_), .Q(instr_sh));
DFFcell _30562_ (.C(clk), .D(_00375_), .Q(instr_addi));
DFFcell _30563_ (.C(clk), .D(_00376_), .Q(instr_slti));
DFFcell _30564_ (.C(clk), .D(_00377_), .Q(instr_sltiu));
DFFcell _30565_ (.C(clk), .D(_00378_), .Q(instr_xori));
DFFcell _30566_ (.C(clk), .D(_00379_), .Q(instr_ori));
DFFcell _30567_ (.C(clk), .D(_00380_), .Q(instr_andi));
DFFcell _30568_ (.C(clk), .D(_00381_), .Q(instr_sb));
DFFcell _30569_ (.C(clk), .D(_00382_), .Q(instr_slli));
DFFcell _30570_ (.C(clk), .D(_00383_), .Q(instr_srli));
DFFcell _30571_ (.C(clk), .D(_00384_), .Q(instr_add));
DFFcell _30572_ (.C(clk), .D(_00385_), .Q(instr_sub));
DFFcell _30573_ (.C(clk), .D(_00386_), .Q(instr_sll));
DFFcell _30574_ (.C(clk), .D(_00387_), .Q(instr_slt));
DFFcell _30575_ (.C(clk), .D(_00388_), .Q(instr_sltu));
DFFcell _30576_ (.C(clk), .D(_00389_), .Q(instr_xor));
DFFcell _30577_ (.C(clk), .D(_00390_), .Q(instr_srl));
DFFcell _30578_ (.C(clk), .D(_00391_), .Q(instr_sra));
DFFcell _30579_ (.C(clk), .D(_00392_), .Q(instr_or));
DFFcell _30580_ (.C(clk), .D(_00393_), .Q(instr_and));
DFFcell _30581_ (.C(clk), .D(_00394_), .Q(instr_srai));
DFFcell _30582_ (.C(clk), .D(_00395_), .Q(instr_rdcycle));
DFFcell _30583_ (.C(clk), .D(_00396_), .Q(instr_rdcycleh));
DFFcell _30584_ (.C(clk), .D(_00397_), .Q(instr_rdinstr));
DFFcell _30585_ (.C(clk), .D(_00398_), .Q(instr_rdinstrh));
DFFcell _30586_ (.C(clk), .D(_00399_), .Q(decoded_rd[0]));
DFFcell _30587_ (.C(clk), .D(_00400_), .Q(decoded_rd[1]));
DFFcell _30588_ (.C(clk), .D(_00401_), .Q(decoded_rd[2]));
DFFcell _30589_ (.C(clk), .D(_00402_), .Q(decoded_rd[3]));
DFFcell _30590_ (.C(clk), .D(_00403_), .Q(decoded_rd[4]));
DFFcell _30591_ (.C(clk), .D(_00404_), .Q(decoded_imm_j[11]));
DFFcell _30592_ (.C(clk), .D(_00405_), .Q(decoded_imm_j[1]));
DFFcell _30593_ (.C(clk), .D(_00406_), .Q(decoded_imm_j[2]));
DFFcell _30594_ (.C(clk), .D(_00407_), .Q(decoded_imm_j[3]));
DFFcell _30595_ (.C(clk), .D(_00408_), .Q(decoded_imm[0]));
DFFcell _30596_ (.C(clk), .D(_00409_), .Q(decoded_imm_j[10]));
DFFcell _30597_ (.C(clk), .D(_00002_), .Q(is_lui_auipc_jal));
DFFcell _30598_ (.C(clk), .D(_00410_), .Q(is_lb_lh_lw_lbu_lhu));
DFFcell _30599_ (.C(clk), .D(_00411_), .Q(is_slli_srli_srai));
DFFcell _30600_ (.C(clk), .D(_00412_), .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
DFFcell _30601_ (.C(clk), .D(_00413_), .Q(is_sll_srl_sra));
DFFcell _30602_ (.C(clk), .D(_00003_), .Q(is_slti_blt_slt));
DFFcell _30603_ (.C(clk), .D(_00004_), .Q(is_sltiu_bltu_sltu));
DFFcell _30604_ (.C(clk), .D(_00414_), .Q(is_beq_bne_blt_bge_bltu_bgeu));
DFFcell _30605_ (.C(clk), .D(_00001_), .Q(is_lbu_lhu_lw));
DFFcell _30606_ (.C(clk), .D(_00415_), .Q(is_lui_auipc_jal_jalr_addi_add_sub));
DFFcell _30607_ (.C(clk), .D(_00416_), .Q(is_alu_reg_imm));
DFFcell _30608_ (.C(clk), .D(_00417_), .Q(is_alu_reg_reg));
DFFcell _30609_ (.C(clk), .D(_00418_), .Q(is_sb_sh_sw));
DFFcell _30610_ (.C(clk), .D(_00419_), .Q(is_compare));
DFFcell _30611_ (.C(clk), .D(_00420_), .Q(mem_instr));
DFFcell _30612_ (.C(clk), .D(_00421_), .Q(mem_rdata_q[7]));
DFFcell _30613_ (.C(clk), .D(_00422_), .Q(mem_rdata_q[8]));
DFFcell _30614_ (.C(clk), .D(_00423_), .Q(mem_rdata_q[9]));
DFFcell _30615_ (.C(clk), .D(_00424_), .Q(mem_rdata_q[10]));
DFFcell _30616_ (.C(clk), .D(_00425_), .Q(mem_rdata_q[11]));
DFFcell _30617_ (.C(clk), .D(_00426_), .Q(mem_rdata_q[12]));
DFFcell _30618_ (.C(clk), .D(_00427_), .Q(mem_rdata_q[13]));
DFFcell _30619_ (.C(clk), .D(_00428_), .Q(mem_rdata_q[14]));
DFFcell _30620_ (.C(clk), .D(_00429_), .Q(mem_rdata_q[15]));
DFFcell _30621_ (.C(clk), .D(_00430_), .Q(mem_rdata_q[16]));
DFFcell _30622_ (.C(clk), .D(_00431_), .Q(mem_rdata_q[17]));
DFFcell _30623_ (.C(clk), .D(_00432_), .Q(mem_rdata_q[18]));
DFFcell _30624_ (.C(clk), .D(_00433_), .Q(mem_rdata_q[19]));
DFFcell _30625_ (.C(clk), .D(_00434_), .Q(mem_rdata_q[20]));
DFFcell _30626_ (.C(clk), .D(_00435_), .Q(mem_rdata_q[21]));
DFFcell _30627_ (.C(clk), .D(_00436_), .Q(mem_rdata_q[22]));
DFFcell _30628_ (.C(clk), .D(_00437_), .Q(mem_rdata_q[23]));
DFFcell _30629_ (.C(clk), .D(_00438_), .Q(mem_rdata_q[24]));
DFFcell _30630_ (.C(clk), .D(_00439_), .Q(mem_rdata_q[25]));
DFFcell _30631_ (.C(clk), .D(_00440_), .Q(mem_rdata_q[26]));
DFFcell _30632_ (.C(clk), .D(_00441_), .Q(mem_rdata_q[27]));
DFFcell _30633_ (.C(clk), .D(_00442_), .Q(mem_rdata_q[28]));
DFFcell _30634_ (.C(clk), .D(_00443_), .Q(mem_rdata_q[29]));
DFFcell _30635_ (.C(clk), .D(_00444_), .Q(mem_rdata_q[30]));
DFFcell _30636_ (.C(clk), .D(_00445_), .Q(mem_rdata_q[31]));
DFFcell _30637_ (.C(clk), .D(_00446_), .Q(mem_addr[2]));
DFFcell _30638_ (.C(clk), .D(_00447_), .Q(mem_addr[3]));
DFFcell _30639_ (.C(clk), .D(_00448_), .Q(mem_addr[4]));
DFFcell _30640_ (.C(clk), .D(_00449_), .Q(mem_addr[5]));
DFFcell _30641_ (.C(clk), .D(_00450_), .Q(mem_addr[6]));
DFFcell _30642_ (.C(clk), .D(_00451_), .Q(mem_addr[7]));
DFFcell _30643_ (.C(clk), .D(_00452_), .Q(mem_addr[8]));
DFFcell _30644_ (.C(clk), .D(_00453_), .Q(mem_addr[9]));
DFFcell _30645_ (.C(clk), .D(_00454_), .Q(mem_addr[10]));
DFFcell _30646_ (.C(clk), .D(_00455_), .Q(mem_addr[11]));
DFFcell _30647_ (.C(clk), .D(_00456_), .Q(mem_addr[12]));
DFFcell _30648_ (.C(clk), .D(_00457_), .Q(mem_addr[13]));
DFFcell _30649_ (.C(clk), .D(_00458_), .Q(mem_addr[14]));
DFFcell _30650_ (.C(clk), .D(_00459_), .Q(mem_addr[15]));
DFFcell _30651_ (.C(clk), .D(_00460_), .Q(mem_addr[16]));
DFFcell _30652_ (.C(clk), .D(_00461_), .Q(mem_addr[17]));
DFFcell _30653_ (.C(clk), .D(_00462_), .Q(mem_addr[18]));
DFFcell _30654_ (.C(clk), .D(_00463_), .Q(mem_addr[19]));
DFFcell _30655_ (.C(clk), .D(_00464_), .Q(mem_addr[20]));
DFFcell _30656_ (.C(clk), .D(_00465_), .Q(mem_addr[21]));
DFFcell _30657_ (.C(clk), .D(_00466_), .Q(mem_addr[22]));
DFFcell _30658_ (.C(clk), .D(_00467_), .Q(mem_addr[23]));
DFFcell _30659_ (.C(clk), .D(_00468_), .Q(mem_addr[24]));
DFFcell _30660_ (.C(clk), .D(_00469_), .Q(mem_addr[25]));
DFFcell _30661_ (.C(clk), .D(_00470_), .Q(mem_addr[26]));
DFFcell _30662_ (.C(clk), .D(_00471_), .Q(mem_addr[27]));
DFFcell _30663_ (.C(clk), .D(_00472_), .Q(mem_addr[28]));
DFFcell _30664_ (.C(clk), .D(_00473_), .Q(mem_addr[29]));
DFFcell _30665_ (.C(clk), .D(_00474_), .Q(mem_addr[30]));
DFFcell _30666_ (.C(clk), .D(_00475_), .Q(mem_addr[31]));
DFFcell _30667_ (.C(clk), .D(_00476_), .Q(mem_wdata[0]));
DFFcell _30668_ (.C(clk), .D(_00477_), .Q(mem_wdata[1]));
DFFcell _30669_ (.C(clk), .D(_00478_), .Q(mem_wdata[2]));
DFFcell _30670_ (.C(clk), .D(_00479_), .Q(mem_wdata[3]));
DFFcell _30671_ (.C(clk), .D(_00480_), .Q(mem_wdata[4]));
DFFcell _30672_ (.C(clk), .D(_00481_), .Q(mem_wdata[5]));
DFFcell _30673_ (.C(clk), .D(_00482_), .Q(mem_wdata[6]));
DFFcell _30674_ (.C(clk), .D(_00483_), .Q(mem_wdata[7]));
DFFcell _30675_ (.C(clk), .D(_00484_), .Q(mem_wdata[8]));
DFFcell _30676_ (.C(clk), .D(_00485_), .Q(mem_wdata[9]));
DFFcell _30677_ (.C(clk), .D(_00486_), .Q(mem_wdata[10]));
DFFcell _30678_ (.C(clk), .D(_00487_), .Q(mem_wdata[11]));
DFFcell _30679_ (.C(clk), .D(_00488_), .Q(mem_wdata[12]));
DFFcell _30680_ (.C(clk), .D(_00489_), .Q(mem_wdata[13]));
DFFcell _30681_ (.C(clk), .D(_00490_), .Q(mem_wdata[14]));
DFFcell _30682_ (.C(clk), .D(_00491_), .Q(mem_wdata[15]));
DFFcell _30683_ (.C(clk), .D(_00492_), .Q(mem_wdata[16]));
DFFcell _30684_ (.C(clk), .D(_00493_), .Q(mem_wdata[17]));
DFFcell _30685_ (.C(clk), .D(_00494_), .Q(mem_wdata[18]));
DFFcell _30686_ (.C(clk), .D(_00495_), .Q(mem_wdata[19]));
DFFcell _30687_ (.C(clk), .D(_00496_), .Q(mem_wdata[20]));
DFFcell _30688_ (.C(clk), .D(_00497_), .Q(mem_wdata[21]));
DFFcell _30689_ (.C(clk), .D(_00498_), .Q(mem_wdata[22]));
DFFcell _30690_ (.C(clk), .D(_00499_), .Q(mem_wdata[23]));
DFFcell _30691_ (.C(clk), .D(_00500_), .Q(mem_wdata[24]));
DFFcell _30692_ (.C(clk), .D(_00501_), .Q(mem_wdata[25]));
DFFcell _30693_ (.C(clk), .D(_00502_), .Q(mem_wdata[26]));
DFFcell _30694_ (.C(clk), .D(_00503_), .Q(mem_wdata[27]));
DFFcell _30695_ (.C(clk), .D(_00504_), .Q(mem_wdata[28]));
DFFcell _30696_ (.C(clk), .D(_00505_), .Q(mem_wdata[29]));
DFFcell _30697_ (.C(clk), .D(_00506_), .Q(mem_wdata[30]));
DFFcell _30698_ (.C(clk), .D(_00507_), .Q(mem_wdata[31]));
DFFcell _30699_ (.C(clk), .D(_00508_), .Q(mem_wstrb[0]));
DFFcell _30700_ (.C(clk), .D(_00509_), .Q(mem_wstrb[1]));
DFFcell _30701_ (.C(clk), .D(_00510_), .Q(mem_wstrb[2]));
DFFcell _30702_ (.C(clk), .D(_00511_), .Q(mem_wstrb[3]));
DFFcell _30703_ (.C(clk), .D(_00512_), .Q(mem_state[0]));
DFFcell _30704_ (.C(clk), .D(_00513_), .Q(mem_state[1]));
DFFcell _30705_ (.C(clk), .D(_00514_), .Q(mem_rdata_q[0]));
DFFcell _30706_ (.C(clk), .D(_00515_), .Q(mem_rdata_q[1]));
DFFcell _30707_ (.C(clk), .D(_00516_), .Q(mem_rdata_q[2]));
DFFcell _30708_ (.C(clk), .D(_00517_), .Q(mem_rdata_q[3]));
DFFcell _30709_ (.C(clk), .D(_00518_), .Q(mem_rdata_q[4]));
DFFcell _30710_ (.C(clk), .D(_00519_), .Q(mem_rdata_q[5]));
DFFcell _30711_ (.C(clk), .D(_00520_), .Q(mem_rdata_q[6]));
DFFcell _30712_ (.C(clk), .D(_00521_), .Q(decoded_imm[31]));
DFFcell _30713_ (.C(clk), .D(_00522_), .Q(decoded_imm[30]));
DFFcell _30714_ (.C(clk), .D(_00523_), .Q(decoded_imm[29]));
DFFcell _30715_ (.C(clk), .D(_00524_), .Q(decoded_imm[28]));
DFFcell _30716_ (.C(clk), .D(_00525_), .Q(decoded_imm[27]));
DFFcell _30717_ (.C(clk), .D(_00526_), .Q(decoded_imm[26]));
DFFcell _30718_ (.C(clk), .D(_00527_), .Q(decoded_imm[25]));
DFFcell _30719_ (.C(clk), .D(_00528_), .Q(decoded_imm[24]));
DFFcell _30720_ (.C(clk), .D(_00529_), .Q(decoded_imm[23]));
DFFcell _30721_ (.C(clk), .D(_00530_), .Q(decoded_imm[22]));
DFFcell _30722_ (.C(clk), .D(_00531_), .Q(decoded_imm[21]));
DFFcell _30723_ (.C(clk), .D(_00532_), .Q(decoded_imm[20]));
DFFcell _30724_ (.C(clk), .D(_00533_), .Q(decoded_imm[19]));
DFFcell _30725_ (.C(clk), .D(_00534_), .Q(decoded_imm[18]));
DFFcell _30726_ (.C(clk), .D(_00535_), .Q(decoded_imm[17]));
DFFcell _30727_ (.C(clk), .D(_00536_), .Q(decoded_imm[16]));
DFFcell _30728_ (.C(clk), .D(_00537_), .Q(decoded_imm[15]));
DFFcell _30729_ (.C(clk), .D(_00538_), .Q(decoded_imm[14]));
DFFcell _30730_ (.C(clk), .D(_00539_), .Q(decoded_imm[13]));
DFFcell _30731_ (.C(clk), .D(_00540_), .Q(decoded_imm[12]));
DFFcell _30732_ (.C(clk), .D(_00541_), .Q(decoded_imm[11]));
DFFcell _30733_ (.C(clk), .D(_00542_), .Q(decoded_imm[10]));
DFFcell _30734_ (.C(clk), .D(_00543_), .Q(decoded_imm[9]));
DFFcell _30735_ (.C(clk), .D(_00544_), .Q(decoded_imm[8]));
DFFcell _30736_ (.C(clk), .D(_00545_), .Q(decoded_imm[7]));
DFFcell _30737_ (.C(clk), .D(_00546_), .Q(decoded_imm[6]));
DFFcell _30738_ (.C(clk), .D(_00547_), .Q(decoded_imm[5]));
DFFcell _30739_ (.C(clk), .D(_00548_), .Q(decoded_imm[4]));
DFFcell _30740_ (.C(clk), .D(_00549_), .Q(decoded_imm[3]));
DFFcell _30741_ (.C(clk), .D(_00550_), .Q(decoded_imm[2]));
DFFcell _30742_ (.C(clk), .D(_00551_), .Q(decoded_imm[1]));
DFFcell _30743_ (.C(clk), .D(_00552_), .Q(reg_next_pc[0]));
DFFcell _30744_ (.C(clk), .D(_00553_), .Q(cpuregs[29][0]));
DFFcell _30745_ (.C(clk), .D(_00554_), .Q(cpuregs[29][1]));
DFFcell _30746_ (.C(clk), .D(_00555_), .Q(cpuregs[29][2]));
DFFcell _30747_ (.C(clk), .D(_00556_), .Q(cpuregs[29][3]));
DFFcell _30748_ (.C(clk), .D(_00557_), .Q(cpuregs[29][4]));
DFFcell _30749_ (.C(clk), .D(_00558_), .Q(cpuregs[29][5]));
DFFcell _30750_ (.C(clk), .D(_00559_), .Q(cpuregs[29][6]));
DFFcell _30751_ (.C(clk), .D(_00560_), .Q(cpuregs[29][7]));
DFFcell _30752_ (.C(clk), .D(_00561_), .Q(cpuregs[29][8]));
DFFcell _30753_ (.C(clk), .D(_00562_), .Q(cpuregs[29][9]));
DFFcell _30754_ (.C(clk), .D(_00563_), .Q(cpuregs[29][10]));
DFFcell _30755_ (.C(clk), .D(_00564_), .Q(cpuregs[29][11]));
DFFcell _30756_ (.C(clk), .D(_00565_), .Q(cpuregs[29][12]));
DFFcell _30757_ (.C(clk), .D(_00566_), .Q(cpuregs[29][13]));
DFFcell _30758_ (.C(clk), .D(_00567_), .Q(cpuregs[29][14]));
DFFcell _30759_ (.C(clk), .D(_00568_), .Q(cpuregs[29][15]));
DFFcell _30760_ (.C(clk), .D(_00569_), .Q(cpuregs[29][16]));
DFFcell _30761_ (.C(clk), .D(_00570_), .Q(cpuregs[29][17]));
DFFcell _30762_ (.C(clk), .D(_00571_), .Q(cpuregs[29][18]));
DFFcell _30763_ (.C(clk), .D(_00572_), .Q(cpuregs[29][19]));
DFFcell _30764_ (.C(clk), .D(_00573_), .Q(cpuregs[29][20]));
DFFcell _30765_ (.C(clk), .D(_00574_), .Q(cpuregs[29][21]));
DFFcell _30766_ (.C(clk), .D(_00575_), .Q(cpuregs[29][22]));
DFFcell _30767_ (.C(clk), .D(_00576_), .Q(cpuregs[29][23]));
DFFcell _30768_ (.C(clk), .D(_00577_), .Q(cpuregs[29][24]));
DFFcell _30769_ (.C(clk), .D(_00578_), .Q(cpuregs[29][25]));
DFFcell _30770_ (.C(clk), .D(_00579_), .Q(cpuregs[29][26]));
DFFcell _30771_ (.C(clk), .D(_00580_), .Q(cpuregs[29][27]));
DFFcell _30772_ (.C(clk), .D(_00581_), .Q(cpuregs[29][28]));
DFFcell _30773_ (.C(clk), .D(_00582_), .Q(cpuregs[29][29]));
DFFcell _30774_ (.C(clk), .D(_00583_), .Q(cpuregs[29][30]));
DFFcell _30775_ (.C(clk), .D(_00584_), .Q(cpuregs[29][31]));
DFFcell _30776_ (.C(clk), .D(_00585_), .Q(decoded_imm_j[4]));
DFFcell _30777_ (.C(clk), .D(_00586_), .Q(count_instr[0]));
DFFcell _30778_ (.C(clk), .D(_00587_), .Q(count_instr[1]));
DFFcell _30779_ (.C(clk), .D(_00588_), .Q(count_instr[2]));
DFFcell _30780_ (.C(clk), .D(_00589_), .Q(count_instr[3]));
DFFcell _30781_ (.C(clk), .D(_00590_), .Q(count_instr[4]));
DFFcell _30782_ (.C(clk), .D(_00591_), .Q(count_instr[5]));
DFFcell _30783_ (.C(clk), .D(_00592_), .Q(count_instr[6]));
DFFcell _30784_ (.C(clk), .D(_00593_), .Q(count_instr[7]));
DFFcell _30785_ (.C(clk), .D(_00594_), .Q(count_instr[8]));
DFFcell _30786_ (.C(clk), .D(_00595_), .Q(count_instr[9]));
DFFcell _30787_ (.C(clk), .D(_00596_), .Q(count_instr[10]));
DFFcell _30788_ (.C(clk), .D(_00597_), .Q(count_instr[11]));
DFFcell _30789_ (.C(clk), .D(_00598_), .Q(count_instr[12]));
DFFcell _30790_ (.C(clk), .D(_00599_), .Q(count_instr[13]));
DFFcell _30791_ (.C(clk), .D(_00600_), .Q(count_instr[14]));
DFFcell _30792_ (.C(clk), .D(_00601_), .Q(count_instr[15]));
DFFcell _30793_ (.C(clk), .D(_00602_), .Q(count_instr[16]));
DFFcell _30794_ (.C(clk), .D(_00603_), .Q(count_instr[17]));
DFFcell _30795_ (.C(clk), .D(_00604_), .Q(count_instr[18]));
DFFcell _30796_ (.C(clk), .D(_00605_), .Q(count_instr[19]));
DFFcell _30797_ (.C(clk), .D(_00606_), .Q(count_instr[20]));
DFFcell _30798_ (.C(clk), .D(_00607_), .Q(count_instr[21]));
DFFcell _30799_ (.C(clk), .D(_00608_), .Q(count_instr[22]));
DFFcell _30800_ (.C(clk), .D(_00609_), .Q(count_instr[23]));
DFFcell _30801_ (.C(clk), .D(_00610_), .Q(count_instr[24]));
DFFcell _30802_ (.C(clk), .D(_00611_), .Q(count_instr[25]));
DFFcell _30803_ (.C(clk), .D(_00612_), .Q(count_instr[26]));
DFFcell _30804_ (.C(clk), .D(_00613_), .Q(count_instr[27]));
DFFcell _30805_ (.C(clk), .D(_00614_), .Q(count_instr[28]));
DFFcell _30806_ (.C(clk), .D(_00615_), .Q(count_instr[29]));
DFFcell _30807_ (.C(clk), .D(_00616_), .Q(count_instr[30]));
DFFcell _30808_ (.C(clk), .D(_00617_), .Q(count_instr[31]));
DFFcell _30809_ (.C(clk), .D(_00618_), .Q(count_instr[32]));
DFFcell _30810_ (.C(clk), .D(_00619_), .Q(count_instr[33]));
DFFcell _30811_ (.C(clk), .D(_00620_), .Q(count_instr[34]));
DFFcell _30812_ (.C(clk), .D(_00621_), .Q(count_instr[35]));
DFFcell _30813_ (.C(clk), .D(_00622_), .Q(count_instr[36]));
DFFcell _30814_ (.C(clk), .D(_00623_), .Q(count_instr[37]));
DFFcell _30815_ (.C(clk), .D(_00624_), .Q(count_instr[38]));
DFFcell _30816_ (.C(clk), .D(_00625_), .Q(count_instr[39]));
DFFcell _30817_ (.C(clk), .D(_00626_), .Q(count_instr[40]));
DFFcell _30818_ (.C(clk), .D(_00627_), .Q(count_instr[41]));
DFFcell _30819_ (.C(clk), .D(_00628_), .Q(count_instr[42]));
DFFcell _30820_ (.C(clk), .D(_00629_), .Q(count_instr[43]));
DFFcell _30821_ (.C(clk), .D(_00630_), .Q(count_instr[44]));
DFFcell _30822_ (.C(clk), .D(_00631_), .Q(count_instr[45]));
DFFcell _30823_ (.C(clk), .D(_00632_), .Q(count_instr[46]));
DFFcell _30824_ (.C(clk), .D(_00633_), .Q(count_instr[47]));
DFFcell _30825_ (.C(clk), .D(_00634_), .Q(count_instr[48]));
DFFcell _30826_ (.C(clk), .D(_00635_), .Q(count_instr[49]));
DFFcell _30827_ (.C(clk), .D(_00636_), .Q(count_instr[50]));
DFFcell _30828_ (.C(clk), .D(_00637_), .Q(count_instr[51]));
DFFcell _30829_ (.C(clk), .D(_00638_), .Q(count_instr[52]));
DFFcell _30830_ (.C(clk), .D(_00639_), .Q(count_instr[53]));
DFFcell _30831_ (.C(clk), .D(_00640_), .Q(count_instr[54]));
DFFcell _30832_ (.C(clk), .D(_00641_), .Q(count_instr[55]));
DFFcell _30833_ (.C(clk), .D(_00642_), .Q(count_instr[56]));
DFFcell _30834_ (.C(clk), .D(_00643_), .Q(count_instr[57]));
DFFcell _30835_ (.C(clk), .D(_00644_), .Q(count_instr[58]));
DFFcell _30836_ (.C(clk), .D(_00645_), .Q(count_instr[59]));
DFFcell _30837_ (.C(clk), .D(_00646_), .Q(count_instr[60]));
DFFcell _30838_ (.C(clk), .D(_00647_), .Q(count_instr[61]));
DFFcell _30839_ (.C(clk), .D(_00648_), .Q(count_instr[62]));
DFFcell _30840_ (.C(clk), .D(_00649_), .Q(count_instr[63]));
DFFcell _30841_ (.C(clk), .D(_00650_), .Q(cpuregs[12][0]));
DFFcell _30842_ (.C(clk), .D(_00651_), .Q(cpuregs[12][1]));
DFFcell _30843_ (.C(clk), .D(_00652_), .Q(cpuregs[12][2]));
DFFcell _30844_ (.C(clk), .D(_00653_), .Q(cpuregs[12][3]));
DFFcell _30845_ (.C(clk), .D(_00654_), .Q(cpuregs[12][4]));
DFFcell _30846_ (.C(clk), .D(_00655_), .Q(cpuregs[12][5]));
DFFcell _30847_ (.C(clk), .D(_00656_), .Q(cpuregs[12][6]));
DFFcell _30848_ (.C(clk), .D(_00657_), .Q(cpuregs[12][7]));
DFFcell _30849_ (.C(clk), .D(_00658_), .Q(cpuregs[12][8]));
DFFcell _30850_ (.C(clk), .D(_00659_), .Q(cpuregs[12][9]));
DFFcell _30851_ (.C(clk), .D(_00660_), .Q(cpuregs[12][10]));
DFFcell _30852_ (.C(clk), .D(_00661_), .Q(cpuregs[12][11]));
DFFcell _30853_ (.C(clk), .D(_00662_), .Q(cpuregs[12][12]));
DFFcell _30854_ (.C(clk), .D(_00663_), .Q(cpuregs[12][13]));
DFFcell _30855_ (.C(clk), .D(_00664_), .Q(cpuregs[12][14]));
DFFcell _30856_ (.C(clk), .D(_00665_), .Q(cpuregs[12][15]));
DFFcell _30857_ (.C(clk), .D(_00666_), .Q(cpuregs[12][16]));
DFFcell _30858_ (.C(clk), .D(_00667_), .Q(cpuregs[12][17]));
DFFcell _30859_ (.C(clk), .D(_00668_), .Q(cpuregs[12][18]));
DFFcell _30860_ (.C(clk), .D(_00669_), .Q(cpuregs[12][19]));
DFFcell _30861_ (.C(clk), .D(_00670_), .Q(cpuregs[12][20]));
DFFcell _30862_ (.C(clk), .D(_00671_), .Q(cpuregs[12][21]));
DFFcell _30863_ (.C(clk), .D(_00672_), .Q(cpuregs[12][22]));
DFFcell _30864_ (.C(clk), .D(_00673_), .Q(cpuregs[12][23]));
DFFcell _30865_ (.C(clk), .D(_00674_), .Q(cpuregs[12][24]));
DFFcell _30866_ (.C(clk), .D(_00675_), .Q(cpuregs[12][25]));
DFFcell _30867_ (.C(clk), .D(_00676_), .Q(cpuregs[12][26]));
DFFcell _30868_ (.C(clk), .D(_00677_), .Q(cpuregs[12][27]));
DFFcell _30869_ (.C(clk), .D(_00678_), .Q(cpuregs[12][28]));
DFFcell _30870_ (.C(clk), .D(_00679_), .Q(cpuregs[12][29]));
DFFcell _30871_ (.C(clk), .D(_00680_), .Q(cpuregs[12][30]));
DFFcell _30872_ (.C(clk), .D(_00681_), .Q(cpuregs[12][31]));
DFFcell _30873_ (.C(clk), .D(_00682_), .Q(cpuregs[3][0]));
DFFcell _30874_ (.C(clk), .D(_00683_), .Q(cpuregs[3][1]));
DFFcell _30875_ (.C(clk), .D(_00684_), .Q(cpuregs[3][2]));
DFFcell _30876_ (.C(clk), .D(_00685_), .Q(cpuregs[3][3]));
DFFcell _30877_ (.C(clk), .D(_00686_), .Q(cpuregs[3][4]));
DFFcell _30878_ (.C(clk), .D(_00687_), .Q(cpuregs[3][5]));
DFFcell _30879_ (.C(clk), .D(_00688_), .Q(cpuregs[3][6]));
DFFcell _30880_ (.C(clk), .D(_00689_), .Q(cpuregs[3][7]));
DFFcell _30881_ (.C(clk), .D(_00690_), .Q(cpuregs[3][8]));
DFFcell _30882_ (.C(clk), .D(_00691_), .Q(cpuregs[3][9]));
DFFcell _30883_ (.C(clk), .D(_00692_), .Q(cpuregs[3][10]));
DFFcell _30884_ (.C(clk), .D(_00693_), .Q(cpuregs[3][11]));
DFFcell _30885_ (.C(clk), .D(_00694_), .Q(cpuregs[3][12]));
DFFcell _30886_ (.C(clk), .D(_00695_), .Q(cpuregs[3][13]));
DFFcell _30887_ (.C(clk), .D(_00696_), .Q(cpuregs[3][14]));
DFFcell _30888_ (.C(clk), .D(_00697_), .Q(cpuregs[3][15]));
DFFcell _30889_ (.C(clk), .D(_00698_), .Q(cpuregs[3][16]));
DFFcell _30890_ (.C(clk), .D(_00699_), .Q(cpuregs[3][17]));
DFFcell _30891_ (.C(clk), .D(_00700_), .Q(cpuregs[3][18]));
DFFcell _30892_ (.C(clk), .D(_00701_), .Q(cpuregs[3][19]));
DFFcell _30893_ (.C(clk), .D(_00702_), .Q(cpuregs[3][20]));
DFFcell _30894_ (.C(clk), .D(_00703_), .Q(cpuregs[3][21]));
DFFcell _30895_ (.C(clk), .D(_00704_), .Q(cpuregs[3][22]));
DFFcell _30896_ (.C(clk), .D(_00705_), .Q(cpuregs[3][23]));
DFFcell _30897_ (.C(clk), .D(_00706_), .Q(cpuregs[3][24]));
DFFcell _30898_ (.C(clk), .D(_00707_), .Q(cpuregs[3][25]));
DFFcell _30899_ (.C(clk), .D(_00708_), .Q(cpuregs[3][26]));
DFFcell _30900_ (.C(clk), .D(_00709_), .Q(cpuregs[3][27]));
DFFcell _30901_ (.C(clk), .D(_00710_), .Q(cpuregs[3][28]));
DFFcell _30902_ (.C(clk), .D(_00711_), .Q(cpuregs[3][29]));
DFFcell _30903_ (.C(clk), .D(_00712_), .Q(cpuregs[3][30]));
DFFcell _30904_ (.C(clk), .D(_00713_), .Q(cpuregs[3][31]));
DFFcell _30905_ (.C(clk), .D(_00714_), .Q(cpuregs[23][0]));
DFFcell _30906_ (.C(clk), .D(_00715_), .Q(cpuregs[23][1]));
DFFcell _30907_ (.C(clk), .D(_00716_), .Q(cpuregs[23][2]));
DFFcell _30908_ (.C(clk), .D(_00717_), .Q(cpuregs[23][3]));
DFFcell _30909_ (.C(clk), .D(_00718_), .Q(cpuregs[23][4]));
DFFcell _30910_ (.C(clk), .D(_00719_), .Q(cpuregs[23][5]));
DFFcell _30911_ (.C(clk), .D(_00720_), .Q(cpuregs[23][6]));
DFFcell _30912_ (.C(clk), .D(_00721_), .Q(cpuregs[23][7]));
DFFcell _30913_ (.C(clk), .D(_00722_), .Q(cpuregs[23][8]));
DFFcell _30914_ (.C(clk), .D(_00723_), .Q(cpuregs[23][9]));
DFFcell _30915_ (.C(clk), .D(_00724_), .Q(cpuregs[23][10]));
DFFcell _30916_ (.C(clk), .D(_00725_), .Q(cpuregs[23][11]));
DFFcell _30917_ (.C(clk), .D(_00726_), .Q(cpuregs[23][12]));
DFFcell _30918_ (.C(clk), .D(_00727_), .Q(cpuregs[23][13]));
DFFcell _30919_ (.C(clk), .D(_00728_), .Q(cpuregs[23][14]));
DFFcell _30920_ (.C(clk), .D(_00729_), .Q(cpuregs[23][15]));
DFFcell _30921_ (.C(clk), .D(_00730_), .Q(cpuregs[23][16]));
DFFcell _30922_ (.C(clk), .D(_00731_), .Q(cpuregs[23][17]));
DFFcell _30923_ (.C(clk), .D(_00732_), .Q(cpuregs[23][18]));
DFFcell _30924_ (.C(clk), .D(_00733_), .Q(cpuregs[23][19]));
DFFcell _30925_ (.C(clk), .D(_00734_), .Q(cpuregs[23][20]));
DFFcell _30926_ (.C(clk), .D(_00735_), .Q(cpuregs[23][21]));
DFFcell _30927_ (.C(clk), .D(_00736_), .Q(cpuregs[23][22]));
DFFcell _30928_ (.C(clk), .D(_00737_), .Q(cpuregs[23][23]));
DFFcell _30929_ (.C(clk), .D(_00738_), .Q(cpuregs[23][24]));
DFFcell _30930_ (.C(clk), .D(_00739_), .Q(cpuregs[23][25]));
DFFcell _30931_ (.C(clk), .D(_00740_), .Q(cpuregs[23][26]));
DFFcell _30932_ (.C(clk), .D(_00741_), .Q(cpuregs[23][27]));
DFFcell _30933_ (.C(clk), .D(_00742_), .Q(cpuregs[23][28]));
DFFcell _30934_ (.C(clk), .D(_00743_), .Q(cpuregs[23][29]));
DFFcell _30935_ (.C(clk), .D(_00744_), .Q(cpuregs[23][30]));
DFFcell _30936_ (.C(clk), .D(_00745_), .Q(cpuregs[23][31]));
DFFcell _30937_ (.C(clk), .D(_00746_), .Q(cpuregs[4][0]));
DFFcell _30938_ (.C(clk), .D(_00747_), .Q(cpuregs[4][1]));
DFFcell _30939_ (.C(clk), .D(_00748_), .Q(cpuregs[4][2]));
DFFcell _30940_ (.C(clk), .D(_00749_), .Q(cpuregs[4][3]));
DFFcell _30941_ (.C(clk), .D(_00750_), .Q(cpuregs[4][4]));
DFFcell _30942_ (.C(clk), .D(_00751_), .Q(cpuregs[4][5]));
DFFcell _30943_ (.C(clk), .D(_00752_), .Q(cpuregs[4][6]));
DFFcell _30944_ (.C(clk), .D(_00753_), .Q(cpuregs[4][7]));
DFFcell _30945_ (.C(clk), .D(_00754_), .Q(cpuregs[4][8]));
DFFcell _30946_ (.C(clk), .D(_00755_), .Q(cpuregs[4][9]));
DFFcell _30947_ (.C(clk), .D(_00756_), .Q(cpuregs[4][10]));
DFFcell _30948_ (.C(clk), .D(_00757_), .Q(cpuregs[4][11]));
DFFcell _30949_ (.C(clk), .D(_00758_), .Q(cpuregs[4][12]));
DFFcell _30950_ (.C(clk), .D(_00759_), .Q(cpuregs[4][13]));
DFFcell _30951_ (.C(clk), .D(_00760_), .Q(cpuregs[4][14]));
DFFcell _30952_ (.C(clk), .D(_00761_), .Q(cpuregs[4][15]));
DFFcell _30953_ (.C(clk), .D(_00762_), .Q(cpuregs[4][16]));
DFFcell _30954_ (.C(clk), .D(_00763_), .Q(cpuregs[4][17]));
DFFcell _30955_ (.C(clk), .D(_00764_), .Q(cpuregs[4][18]));
DFFcell _30956_ (.C(clk), .D(_00765_), .Q(cpuregs[4][19]));
DFFcell _30957_ (.C(clk), .D(_00766_), .Q(cpuregs[4][20]));
DFFcell _30958_ (.C(clk), .D(_00767_), .Q(cpuregs[4][21]));
DFFcell _30959_ (.C(clk), .D(_00768_), .Q(cpuregs[4][22]));
DFFcell _30960_ (.C(clk), .D(_00769_), .Q(cpuregs[4][23]));
DFFcell _30961_ (.C(clk), .D(_00770_), .Q(cpuregs[4][24]));
DFFcell _30962_ (.C(clk), .D(_00771_), .Q(cpuregs[4][25]));
DFFcell _30963_ (.C(clk), .D(_00772_), .Q(cpuregs[4][26]));
DFFcell _30964_ (.C(clk), .D(_00773_), .Q(cpuregs[4][27]));
DFFcell _30965_ (.C(clk), .D(_00774_), .Q(cpuregs[4][28]));
DFFcell _30966_ (.C(clk), .D(_00775_), .Q(cpuregs[4][29]));
DFFcell _30967_ (.C(clk), .D(_00776_), .Q(cpuregs[4][30]));
DFFcell _30968_ (.C(clk), .D(_00777_), .Q(cpuregs[4][31]));
DFFcell _30969_ (.C(clk), .D(_00778_), .Q(cpuregs[22][0]));
DFFcell _30970_ (.C(clk), .D(_00779_), .Q(cpuregs[22][1]));
DFFcell _30971_ (.C(clk), .D(_00780_), .Q(cpuregs[22][2]));
DFFcell _30972_ (.C(clk), .D(_00781_), .Q(cpuregs[22][3]));
DFFcell _30973_ (.C(clk), .D(_00782_), .Q(cpuregs[22][4]));
DFFcell _30974_ (.C(clk), .D(_00783_), .Q(cpuregs[22][5]));
DFFcell _30975_ (.C(clk), .D(_00784_), .Q(cpuregs[22][6]));
DFFcell _30976_ (.C(clk), .D(_00785_), .Q(cpuregs[22][7]));
DFFcell _30977_ (.C(clk), .D(_00786_), .Q(cpuregs[22][8]));
DFFcell _30978_ (.C(clk), .D(_00787_), .Q(cpuregs[22][9]));
DFFcell _30979_ (.C(clk), .D(_00788_), .Q(cpuregs[22][10]));
DFFcell _30980_ (.C(clk), .D(_00789_), .Q(cpuregs[22][11]));
DFFcell _30981_ (.C(clk), .D(_00790_), .Q(cpuregs[22][12]));
DFFcell _30982_ (.C(clk), .D(_00791_), .Q(cpuregs[22][13]));
DFFcell _30983_ (.C(clk), .D(_00792_), .Q(cpuregs[22][14]));
DFFcell _30984_ (.C(clk), .D(_00793_), .Q(cpuregs[22][15]));
DFFcell _30985_ (.C(clk), .D(_00794_), .Q(cpuregs[22][16]));
DFFcell _30986_ (.C(clk), .D(_00795_), .Q(cpuregs[22][17]));
DFFcell _30987_ (.C(clk), .D(_00796_), .Q(cpuregs[22][18]));
DFFcell _30988_ (.C(clk), .D(_00797_), .Q(cpuregs[22][19]));
DFFcell _30989_ (.C(clk), .D(_00798_), .Q(cpuregs[22][20]));
DFFcell _30990_ (.C(clk), .D(_00799_), .Q(cpuregs[22][21]));
DFFcell _30991_ (.C(clk), .D(_00800_), .Q(cpuregs[22][22]));
DFFcell _30992_ (.C(clk), .D(_00801_), .Q(cpuregs[22][23]));
DFFcell _30993_ (.C(clk), .D(_00802_), .Q(cpuregs[22][24]));
DFFcell _30994_ (.C(clk), .D(_00803_), .Q(cpuregs[22][25]));
DFFcell _30995_ (.C(clk), .D(_00804_), .Q(cpuregs[22][26]));
DFFcell _30996_ (.C(clk), .D(_00805_), .Q(cpuregs[22][27]));
DFFcell _30997_ (.C(clk), .D(_00806_), .Q(cpuregs[22][28]));
DFFcell _30998_ (.C(clk), .D(_00807_), .Q(cpuregs[22][29]));
DFFcell _30999_ (.C(clk), .D(_00808_), .Q(cpuregs[22][30]));
DFFcell _31000_ (.C(clk), .D(_00809_), .Q(cpuregs[22][31]));
DFFcell _31001_ (.C(clk), .D(_00810_), .Q(cpuregs[13][0]));
DFFcell _31002_ (.C(clk), .D(_00811_), .Q(cpuregs[13][1]));
DFFcell _31003_ (.C(clk), .D(_00812_), .Q(cpuregs[13][2]));
DFFcell _31004_ (.C(clk), .D(_00813_), .Q(cpuregs[13][3]));
DFFcell _31005_ (.C(clk), .D(_00814_), .Q(cpuregs[13][4]));
DFFcell _31006_ (.C(clk), .D(_00815_), .Q(cpuregs[13][5]));
DFFcell _31007_ (.C(clk), .D(_00816_), .Q(cpuregs[13][6]));
DFFcell _31008_ (.C(clk), .D(_00817_), .Q(cpuregs[13][7]));
DFFcell _31009_ (.C(clk), .D(_00818_), .Q(cpuregs[13][8]));
DFFcell _31010_ (.C(clk), .D(_00819_), .Q(cpuregs[13][9]));
DFFcell _31011_ (.C(clk), .D(_00820_), .Q(cpuregs[13][10]));
DFFcell _31012_ (.C(clk), .D(_00821_), .Q(cpuregs[13][11]));
DFFcell _31013_ (.C(clk), .D(_00822_), .Q(cpuregs[13][12]));
DFFcell _31014_ (.C(clk), .D(_00823_), .Q(cpuregs[13][13]));
DFFcell _31015_ (.C(clk), .D(_00824_), .Q(cpuregs[13][14]));
DFFcell _31016_ (.C(clk), .D(_00825_), .Q(cpuregs[13][15]));
DFFcell _31017_ (.C(clk), .D(_00826_), .Q(cpuregs[13][16]));
DFFcell _31018_ (.C(clk), .D(_00827_), .Q(cpuregs[13][17]));
DFFcell _31019_ (.C(clk), .D(_00828_), .Q(cpuregs[13][18]));
DFFcell _31020_ (.C(clk), .D(_00829_), .Q(cpuregs[13][19]));
DFFcell _31021_ (.C(clk), .D(_00830_), .Q(cpuregs[13][20]));
DFFcell _31022_ (.C(clk), .D(_00831_), .Q(cpuregs[13][21]));
DFFcell _31023_ (.C(clk), .D(_00832_), .Q(cpuregs[13][22]));
DFFcell _31024_ (.C(clk), .D(_00833_), .Q(cpuregs[13][23]));
DFFcell _31025_ (.C(clk), .D(_00834_), .Q(cpuregs[13][24]));
DFFcell _31026_ (.C(clk), .D(_00835_), .Q(cpuregs[13][25]));
DFFcell _31027_ (.C(clk), .D(_00836_), .Q(cpuregs[13][26]));
DFFcell _31028_ (.C(clk), .D(_00837_), .Q(cpuregs[13][27]));
DFFcell _31029_ (.C(clk), .D(_00838_), .Q(cpuregs[13][28]));
DFFcell _31030_ (.C(clk), .D(_00839_), .Q(cpuregs[13][29]));
DFFcell _31031_ (.C(clk), .D(_00840_), .Q(cpuregs[13][30]));
DFFcell _31032_ (.C(clk), .D(_00841_), .Q(cpuregs[13][31]));
DFFcell _31033_ (.C(clk), .D(_00842_), .Q(cpuregs[11][0]));
DFFcell _31034_ (.C(clk), .D(_00843_), .Q(cpuregs[11][1]));
DFFcell _31035_ (.C(clk), .D(_00844_), .Q(cpuregs[11][2]));
DFFcell _31036_ (.C(clk), .D(_00845_), .Q(cpuregs[11][3]));
DFFcell _31037_ (.C(clk), .D(_00846_), .Q(cpuregs[11][4]));
DFFcell _31038_ (.C(clk), .D(_00847_), .Q(cpuregs[11][5]));
DFFcell _31039_ (.C(clk), .D(_00848_), .Q(cpuregs[11][6]));
DFFcell _31040_ (.C(clk), .D(_00849_), .Q(cpuregs[11][7]));
DFFcell _31041_ (.C(clk), .D(_00850_), .Q(cpuregs[11][8]));
DFFcell _31042_ (.C(clk), .D(_00851_), .Q(cpuregs[11][9]));
DFFcell _31043_ (.C(clk), .D(_00852_), .Q(cpuregs[11][10]));
DFFcell _31044_ (.C(clk), .D(_00853_), .Q(cpuregs[11][11]));
DFFcell _31045_ (.C(clk), .D(_00854_), .Q(cpuregs[11][12]));
DFFcell _31046_ (.C(clk), .D(_00855_), .Q(cpuregs[11][13]));
DFFcell _31047_ (.C(clk), .D(_00856_), .Q(cpuregs[11][14]));
DFFcell _31048_ (.C(clk), .D(_00857_), .Q(cpuregs[11][15]));
DFFcell _31049_ (.C(clk), .D(_00858_), .Q(cpuregs[11][16]));
DFFcell _31050_ (.C(clk), .D(_00859_), .Q(cpuregs[11][17]));
DFFcell _31051_ (.C(clk), .D(_00860_), .Q(cpuregs[11][18]));
DFFcell _31052_ (.C(clk), .D(_00861_), .Q(cpuregs[11][19]));
DFFcell _31053_ (.C(clk), .D(_00862_), .Q(cpuregs[11][20]));
DFFcell _31054_ (.C(clk), .D(_00863_), .Q(cpuregs[11][21]));
DFFcell _31055_ (.C(clk), .D(_00864_), .Q(cpuregs[11][22]));
DFFcell _31056_ (.C(clk), .D(_00865_), .Q(cpuregs[11][23]));
DFFcell _31057_ (.C(clk), .D(_00866_), .Q(cpuregs[11][24]));
DFFcell _31058_ (.C(clk), .D(_00867_), .Q(cpuregs[11][25]));
DFFcell _31059_ (.C(clk), .D(_00868_), .Q(cpuregs[11][26]));
DFFcell _31060_ (.C(clk), .D(_00869_), .Q(cpuregs[11][27]));
DFFcell _31061_ (.C(clk), .D(_00870_), .Q(cpuregs[11][28]));
DFFcell _31062_ (.C(clk), .D(_00871_), .Q(cpuregs[11][29]));
DFFcell _31063_ (.C(clk), .D(_00872_), .Q(cpuregs[11][30]));
DFFcell _31064_ (.C(clk), .D(_00873_), .Q(cpuregs[11][31]));
DFFcell _31065_ (.C(clk), .D(_00874_), .Q(cpuregs[18][0]));
DFFcell _31066_ (.C(clk), .D(_00875_), .Q(cpuregs[18][1]));
DFFcell _31067_ (.C(clk), .D(_00876_), .Q(cpuregs[18][2]));
DFFcell _31068_ (.C(clk), .D(_00877_), .Q(cpuregs[18][3]));
DFFcell _31069_ (.C(clk), .D(_00878_), .Q(cpuregs[18][4]));
DFFcell _31070_ (.C(clk), .D(_00879_), .Q(cpuregs[18][5]));
DFFcell _31071_ (.C(clk), .D(_00880_), .Q(cpuregs[18][6]));
DFFcell _31072_ (.C(clk), .D(_00881_), .Q(cpuregs[18][7]));
DFFcell _31073_ (.C(clk), .D(_00882_), .Q(cpuregs[18][8]));
DFFcell _31074_ (.C(clk), .D(_00883_), .Q(cpuregs[18][9]));
DFFcell _31075_ (.C(clk), .D(_00884_), .Q(cpuregs[18][10]));
DFFcell _31076_ (.C(clk), .D(_00885_), .Q(cpuregs[18][11]));
DFFcell _31077_ (.C(clk), .D(_00886_), .Q(cpuregs[18][12]));
DFFcell _31078_ (.C(clk), .D(_00887_), .Q(cpuregs[18][13]));
DFFcell _31079_ (.C(clk), .D(_00888_), .Q(cpuregs[18][14]));
DFFcell _31080_ (.C(clk), .D(_00889_), .Q(cpuregs[18][15]));
DFFcell _31081_ (.C(clk), .D(_00890_), .Q(cpuregs[18][16]));
DFFcell _31082_ (.C(clk), .D(_00891_), .Q(cpuregs[18][17]));
DFFcell _31083_ (.C(clk), .D(_00892_), .Q(cpuregs[18][18]));
DFFcell _31084_ (.C(clk), .D(_00893_), .Q(cpuregs[18][19]));
DFFcell _31085_ (.C(clk), .D(_00894_), .Q(cpuregs[18][20]));
DFFcell _31086_ (.C(clk), .D(_00895_), .Q(cpuregs[18][21]));
DFFcell _31087_ (.C(clk), .D(_00896_), .Q(cpuregs[18][22]));
DFFcell _31088_ (.C(clk), .D(_00897_), .Q(cpuregs[18][23]));
DFFcell _31089_ (.C(clk), .D(_00898_), .Q(cpuregs[18][24]));
DFFcell _31090_ (.C(clk), .D(_00899_), .Q(cpuregs[18][25]));
DFFcell _31091_ (.C(clk), .D(_00900_), .Q(cpuregs[18][26]));
DFFcell _31092_ (.C(clk), .D(_00901_), .Q(cpuregs[18][27]));
DFFcell _31093_ (.C(clk), .D(_00902_), .Q(cpuregs[18][28]));
DFFcell _31094_ (.C(clk), .D(_00903_), .Q(cpuregs[18][29]));
DFFcell _31095_ (.C(clk), .D(_00904_), .Q(cpuregs[18][30]));
DFFcell _31096_ (.C(clk), .D(_00905_), .Q(cpuregs[18][31]));
DFFcell _31097_ (.C(clk), .D(_00906_), .Q(cpuregs[14][0]));
DFFcell _31098_ (.C(clk), .D(_00907_), .Q(cpuregs[14][1]));
DFFcell _31099_ (.C(clk), .D(_00908_), .Q(cpuregs[14][2]));
DFFcell _31100_ (.C(clk), .D(_00909_), .Q(cpuregs[14][3]));
DFFcell _31101_ (.C(clk), .D(_00910_), .Q(cpuregs[14][4]));
DFFcell _31102_ (.C(clk), .D(_00911_), .Q(cpuregs[14][5]));
DFFcell _31103_ (.C(clk), .D(_00912_), .Q(cpuregs[14][6]));
DFFcell _31104_ (.C(clk), .D(_00913_), .Q(cpuregs[14][7]));
DFFcell _31105_ (.C(clk), .D(_00914_), .Q(cpuregs[14][8]));
DFFcell _31106_ (.C(clk), .D(_00915_), .Q(cpuregs[14][9]));
DFFcell _31107_ (.C(clk), .D(_00916_), .Q(cpuregs[14][10]));
DFFcell _31108_ (.C(clk), .D(_00917_), .Q(cpuregs[14][11]));
DFFcell _31109_ (.C(clk), .D(_00918_), .Q(cpuregs[14][12]));
DFFcell _31110_ (.C(clk), .D(_00919_), .Q(cpuregs[14][13]));
DFFcell _31111_ (.C(clk), .D(_00920_), .Q(cpuregs[14][14]));
DFFcell _31112_ (.C(clk), .D(_00921_), .Q(cpuregs[14][15]));
DFFcell _31113_ (.C(clk), .D(_00922_), .Q(cpuregs[14][16]));
DFFcell _31114_ (.C(clk), .D(_00923_), .Q(cpuregs[14][17]));
DFFcell _31115_ (.C(clk), .D(_00924_), .Q(cpuregs[14][18]));
DFFcell _31116_ (.C(clk), .D(_00925_), .Q(cpuregs[14][19]));
DFFcell _31117_ (.C(clk), .D(_00926_), .Q(cpuregs[14][20]));
DFFcell _31118_ (.C(clk), .D(_00927_), .Q(cpuregs[14][21]));
DFFcell _31119_ (.C(clk), .D(_00928_), .Q(cpuregs[14][22]));
DFFcell _31120_ (.C(clk), .D(_00929_), .Q(cpuregs[14][23]));
DFFcell _31121_ (.C(clk), .D(_00930_), .Q(cpuregs[14][24]));
DFFcell _31122_ (.C(clk), .D(_00931_), .Q(cpuregs[14][25]));
DFFcell _31123_ (.C(clk), .D(_00932_), .Q(cpuregs[14][26]));
DFFcell _31124_ (.C(clk), .D(_00933_), .Q(cpuregs[14][27]));
DFFcell _31125_ (.C(clk), .D(_00934_), .Q(cpuregs[14][28]));
DFFcell _31126_ (.C(clk), .D(_00935_), .Q(cpuregs[14][29]));
DFFcell _31127_ (.C(clk), .D(_00936_), .Q(cpuregs[14][30]));
DFFcell _31128_ (.C(clk), .D(_00937_), .Q(cpuregs[14][31]));
DFFcell _31129_ (.C(clk), .D(_00938_), .Q(cpuregs[17][0]));
DFFcell _31130_ (.C(clk), .D(_00939_), .Q(cpuregs[17][1]));
DFFcell _31131_ (.C(clk), .D(_00940_), .Q(cpuregs[17][2]));
DFFcell _31132_ (.C(clk), .D(_00941_), .Q(cpuregs[17][3]));
DFFcell _31133_ (.C(clk), .D(_00942_), .Q(cpuregs[17][4]));
DFFcell _31134_ (.C(clk), .D(_00943_), .Q(cpuregs[17][5]));
DFFcell _31135_ (.C(clk), .D(_00944_), .Q(cpuregs[17][6]));
DFFcell _31136_ (.C(clk), .D(_00945_), .Q(cpuregs[17][7]));
DFFcell _31137_ (.C(clk), .D(_00946_), .Q(cpuregs[17][8]));
DFFcell _31138_ (.C(clk), .D(_00947_), .Q(cpuregs[17][9]));
DFFcell _31139_ (.C(clk), .D(_00948_), .Q(cpuregs[17][10]));
DFFcell _31140_ (.C(clk), .D(_00949_), .Q(cpuregs[17][11]));
DFFcell _31141_ (.C(clk), .D(_00950_), .Q(cpuregs[17][12]));
DFFcell _31142_ (.C(clk), .D(_00951_), .Q(cpuregs[17][13]));
DFFcell _31143_ (.C(clk), .D(_00952_), .Q(cpuregs[17][14]));
DFFcell _31144_ (.C(clk), .D(_00953_), .Q(cpuregs[17][15]));
DFFcell _31145_ (.C(clk), .D(_00954_), .Q(cpuregs[17][16]));
DFFcell _31146_ (.C(clk), .D(_00955_), .Q(cpuregs[17][17]));
DFFcell _31147_ (.C(clk), .D(_00956_), .Q(cpuregs[17][18]));
DFFcell _31148_ (.C(clk), .D(_00957_), .Q(cpuregs[17][19]));
DFFcell _31149_ (.C(clk), .D(_00958_), .Q(cpuregs[17][20]));
DFFcell _31150_ (.C(clk), .D(_00959_), .Q(cpuregs[17][21]));
DFFcell _31151_ (.C(clk), .D(_00960_), .Q(cpuregs[17][22]));
DFFcell _31152_ (.C(clk), .D(_00961_), .Q(cpuregs[17][23]));
DFFcell _31153_ (.C(clk), .D(_00962_), .Q(cpuregs[17][24]));
DFFcell _31154_ (.C(clk), .D(_00963_), .Q(cpuregs[17][25]));
DFFcell _31155_ (.C(clk), .D(_00964_), .Q(cpuregs[17][26]));
DFFcell _31156_ (.C(clk), .D(_00965_), .Q(cpuregs[17][27]));
DFFcell _31157_ (.C(clk), .D(_00966_), .Q(cpuregs[17][28]));
DFFcell _31158_ (.C(clk), .D(_00967_), .Q(cpuregs[17][29]));
DFFcell _31159_ (.C(clk), .D(_00968_), .Q(cpuregs[17][30]));
DFFcell _31160_ (.C(clk), .D(_00969_), .Q(cpuregs[17][31]));
DFFcell _31161_ (.C(clk), .D(_00970_), .Q(decoded_imm_j[12]));
DFFcell _31162_ (.C(clk), .D(_00971_), .Q(decoded_imm_j[13]));
DFFcell _31163_ (.C(clk), .D(_00972_), .Q(decoded_imm_j[14]));
DFFcell _31164_ (.C(clk), .D(_00973_), .Q(decoded_imm_j[15]));
DFFcell _31165_ (.C(clk), .D(_00974_), .Q(decoded_imm_j[16]));
DFFcell _31166_ (.C(clk), .D(_00975_), .Q(decoded_imm_j[17]));
DFFcell _31167_ (.C(clk), .D(_00976_), .Q(decoded_imm_j[18]));
DFFcell _31168_ (.C(clk), .D(_00977_), .Q(decoded_imm_j[19]));
DFFcell _31169_ (.C(clk), .D(_00978_), .Q(cpu_state[0]));
DFFcell _31170_ (.C(clk), .D(_00979_), .Q(cpu_state[1]));
DFFcell _31171_ (.C(clk), .D(_00980_), .Q(cpu_state[2]));
DFFcell _31172_ (.C(clk), .D(_00981_), .Q(cpu_state[3]));
DFFcell _31173_ (.C(clk), .D(_00982_), .Q(cpu_state[4]));
DFFcell _31174_ (.C(clk), .D(_00983_), .Q(cpu_state[5]));
DFFcell _31175_ (.C(clk), .D(_00984_), .Q(cpu_state[6]));
DFFcell _31176_ (.C(clk), .D(_00985_), .Q(cpu_state[7]));
DFFcell _31177_ (.C(clk), .D(_00986_), .Q(cpuregs[5][0]));
DFFcell _31178_ (.C(clk), .D(_00987_), .Q(cpuregs[5][1]));
DFFcell _31179_ (.C(clk), .D(_00988_), .Q(cpuregs[5][2]));
DFFcell _31180_ (.C(clk), .D(_00989_), .Q(cpuregs[5][3]));
DFFcell _31181_ (.C(clk), .D(_00990_), .Q(cpuregs[5][4]));
DFFcell _31182_ (.C(clk), .D(_00991_), .Q(cpuregs[5][5]));
DFFcell _31183_ (.C(clk), .D(_00992_), .Q(cpuregs[5][6]));
DFFcell _31184_ (.C(clk), .D(_00993_), .Q(cpuregs[5][7]));
DFFcell _31185_ (.C(clk), .D(_00994_), .Q(cpuregs[5][8]));
DFFcell _31186_ (.C(clk), .D(_00995_), .Q(cpuregs[5][9]));
DFFcell _31187_ (.C(clk), .D(_00996_), .Q(cpuregs[5][10]));
DFFcell _31188_ (.C(clk), .D(_00997_), .Q(cpuregs[5][11]));
DFFcell _31189_ (.C(clk), .D(_00998_), .Q(cpuregs[5][12]));
DFFcell _31190_ (.C(clk), .D(_00999_), .Q(cpuregs[5][13]));
DFFcell _31191_ (.C(clk), .D(_01000_), .Q(cpuregs[5][14]));
DFFcell _31192_ (.C(clk), .D(_01001_), .Q(cpuregs[5][15]));
DFFcell _31193_ (.C(clk), .D(_01002_), .Q(cpuregs[5][16]));
DFFcell _31194_ (.C(clk), .D(_01003_), .Q(cpuregs[5][17]));
DFFcell _31195_ (.C(clk), .D(_01004_), .Q(cpuregs[5][18]));
DFFcell _31196_ (.C(clk), .D(_01005_), .Q(cpuregs[5][19]));
DFFcell _31197_ (.C(clk), .D(_01006_), .Q(cpuregs[5][20]));
DFFcell _31198_ (.C(clk), .D(_01007_), .Q(cpuregs[5][21]));
DFFcell _31199_ (.C(clk), .D(_01008_), .Q(cpuregs[5][22]));
DFFcell _31200_ (.C(clk), .D(_01009_), .Q(cpuregs[5][23]));
DFFcell _31201_ (.C(clk), .D(_01010_), .Q(cpuregs[5][24]));
DFFcell _31202_ (.C(clk), .D(_01011_), .Q(cpuregs[5][25]));
DFFcell _31203_ (.C(clk), .D(_01012_), .Q(cpuregs[5][26]));
DFFcell _31204_ (.C(clk), .D(_01013_), .Q(cpuregs[5][27]));
DFFcell _31205_ (.C(clk), .D(_01014_), .Q(cpuregs[5][28]));
DFFcell _31206_ (.C(clk), .D(_01015_), .Q(cpuregs[5][29]));
DFFcell _31207_ (.C(clk), .D(_01016_), .Q(cpuregs[5][30]));
DFFcell _31208_ (.C(clk), .D(_01017_), .Q(cpuregs[5][31]));
DFFcell _31209_ (.C(clk), .D(_01018_), .Q(pcpi_rs1[0]));
DFFcell _31210_ (.C(clk), .D(_01019_), .Q(pcpi_rs1[1]));
DFFcell _31211_ (.C(clk), .D(_01020_), .Q(pcpi_rs1[2]));
DFFcell _31212_ (.C(clk), .D(_01021_), .Q(pcpi_rs1[3]));
DFFcell _31213_ (.C(clk), .D(_01022_), .Q(pcpi_rs1[4]));
DFFcell _31214_ (.C(clk), .D(_01023_), .Q(pcpi_rs1[5]));
DFFcell _31215_ (.C(clk), .D(_01024_), .Q(pcpi_rs1[6]));
DFFcell _31216_ (.C(clk), .D(_01025_), .Q(pcpi_rs1[7]));
DFFcell _31217_ (.C(clk), .D(_01026_), .Q(pcpi_rs1[8]));
DFFcell _31218_ (.C(clk), .D(_01027_), .Q(pcpi_rs1[9]));
DFFcell _31219_ (.C(clk), .D(_01028_), .Q(pcpi_rs1[10]));
DFFcell _31220_ (.C(clk), .D(_01029_), .Q(pcpi_rs1[11]));
DFFcell _31221_ (.C(clk), .D(_01030_), .Q(pcpi_rs1[12]));
DFFcell _31222_ (.C(clk), .D(_01031_), .Q(pcpi_rs1[13]));
DFFcell _31223_ (.C(clk), .D(_01032_), .Q(pcpi_rs1[14]));
DFFcell _31224_ (.C(clk), .D(_01033_), .Q(pcpi_rs1[15]));
DFFcell _31225_ (.C(clk), .D(_01034_), .Q(pcpi_rs1[16]));
DFFcell _31226_ (.C(clk), .D(_01035_), .Q(pcpi_rs1[17]));
DFFcell _31227_ (.C(clk), .D(_01036_), .Q(pcpi_rs1[18]));
DFFcell _31228_ (.C(clk), .D(_01037_), .Q(pcpi_rs1[19]));
DFFcell _31229_ (.C(clk), .D(_01038_), .Q(pcpi_rs1[20]));
DFFcell _31230_ (.C(clk), .D(_01039_), .Q(pcpi_rs1[21]));
DFFcell _31231_ (.C(clk), .D(_01040_), .Q(pcpi_rs1[22]));
DFFcell _31232_ (.C(clk), .D(_01041_), .Q(pcpi_rs1[23]));
DFFcell _31233_ (.C(clk), .D(_01042_), .Q(pcpi_rs1[24]));
DFFcell _31234_ (.C(clk), .D(_01043_), .Q(pcpi_rs1[25]));
DFFcell _31235_ (.C(clk), .D(_01044_), .Q(pcpi_rs1[26]));
DFFcell _31236_ (.C(clk), .D(_01045_), .Q(pcpi_rs1[27]));
DFFcell _31237_ (.C(clk), .D(_01046_), .Q(pcpi_rs1[28]));
DFFcell _31238_ (.C(clk), .D(_01047_), .Q(pcpi_rs1[29]));
DFFcell _31239_ (.C(clk), .D(_01048_), .Q(pcpi_rs1[30]));
DFFcell _31240_ (.C(clk), .D(_01049_), .Q(cpuregs[7][0]));
DFFcell _31241_ (.C(clk), .D(_01050_), .Q(cpuregs[7][1]));
DFFcell _31242_ (.C(clk), .D(_01051_), .Q(cpuregs[7][2]));
DFFcell _31243_ (.C(clk), .D(_01052_), .Q(cpuregs[7][3]));
DFFcell _31244_ (.C(clk), .D(_01053_), .Q(cpuregs[7][4]));
DFFcell _31245_ (.C(clk), .D(_01054_), .Q(cpuregs[7][5]));
DFFcell _31246_ (.C(clk), .D(_01055_), .Q(cpuregs[7][6]));
DFFcell _31247_ (.C(clk), .D(_01056_), .Q(cpuregs[7][7]));
DFFcell _31248_ (.C(clk), .D(_01057_), .Q(cpuregs[7][8]));
DFFcell _31249_ (.C(clk), .D(_01058_), .Q(cpuregs[7][9]));
DFFcell _31250_ (.C(clk), .D(_01059_), .Q(cpuregs[7][10]));
DFFcell _31251_ (.C(clk), .D(_01060_), .Q(cpuregs[7][11]));
DFFcell _31252_ (.C(clk), .D(_01061_), .Q(cpuregs[7][12]));
DFFcell _31253_ (.C(clk), .D(_01062_), .Q(cpuregs[7][13]));
DFFcell _31254_ (.C(clk), .D(_01063_), .Q(cpuregs[7][14]));
DFFcell _31255_ (.C(clk), .D(_01064_), .Q(cpuregs[7][15]));
DFFcell _31256_ (.C(clk), .D(_01065_), .Q(cpuregs[7][16]));
DFFcell _31257_ (.C(clk), .D(_01066_), .Q(cpuregs[7][17]));
DFFcell _31258_ (.C(clk), .D(_01067_), .Q(cpuregs[7][18]));
DFFcell _31259_ (.C(clk), .D(_01068_), .Q(cpuregs[7][19]));
DFFcell _31260_ (.C(clk), .D(_01069_), .Q(cpuregs[7][20]));
DFFcell _31261_ (.C(clk), .D(_01070_), .Q(cpuregs[7][21]));
DFFcell _31262_ (.C(clk), .D(_01071_), .Q(cpuregs[7][22]));
DFFcell _31263_ (.C(clk), .D(_01072_), .Q(cpuregs[7][23]));
DFFcell _31264_ (.C(clk), .D(_01073_), .Q(cpuregs[7][24]));
DFFcell _31265_ (.C(clk), .D(_01074_), .Q(cpuregs[7][25]));
DFFcell _31266_ (.C(clk), .D(_01075_), .Q(cpuregs[7][26]));
DFFcell _31267_ (.C(clk), .D(_01076_), .Q(cpuregs[7][27]));
DFFcell _31268_ (.C(clk), .D(_01077_), .Q(cpuregs[7][28]));
DFFcell _31269_ (.C(clk), .D(_01078_), .Q(cpuregs[7][29]));
DFFcell _31270_ (.C(clk), .D(_01079_), .Q(cpuregs[7][30]));
DFFcell _31271_ (.C(clk), .D(_01080_), .Q(cpuregs[7][31]));
DFFcell _31272_ (.C(clk), .D(_01081_), .Q(cpuregs[8][0]));
DFFcell _31273_ (.C(clk), .D(_01082_), .Q(cpuregs[8][1]));
DFFcell _31274_ (.C(clk), .D(_01083_), .Q(cpuregs[8][2]));
DFFcell _31275_ (.C(clk), .D(_01084_), .Q(cpuregs[8][3]));
DFFcell _31276_ (.C(clk), .D(_01085_), .Q(cpuregs[8][4]));
DFFcell _31277_ (.C(clk), .D(_01086_), .Q(cpuregs[8][5]));
DFFcell _31278_ (.C(clk), .D(_01087_), .Q(cpuregs[8][6]));
DFFcell _31279_ (.C(clk), .D(_01088_), .Q(cpuregs[8][7]));
DFFcell _31280_ (.C(clk), .D(_01089_), .Q(cpuregs[8][8]));
DFFcell _31281_ (.C(clk), .D(_01090_), .Q(cpuregs[8][9]));
DFFcell _31282_ (.C(clk), .D(_01091_), .Q(cpuregs[8][10]));
DFFcell _31283_ (.C(clk), .D(_01092_), .Q(cpuregs[8][11]));
DFFcell _31284_ (.C(clk), .D(_01093_), .Q(cpuregs[8][12]));
DFFcell _31285_ (.C(clk), .D(_01094_), .Q(cpuregs[8][13]));
DFFcell _31286_ (.C(clk), .D(_01095_), .Q(cpuregs[8][14]));
DFFcell _31287_ (.C(clk), .D(_01096_), .Q(cpuregs[8][15]));
DFFcell _31288_ (.C(clk), .D(_01097_), .Q(cpuregs[8][16]));
DFFcell _31289_ (.C(clk), .D(_01098_), .Q(cpuregs[8][17]));
DFFcell _31290_ (.C(clk), .D(_01099_), .Q(cpuregs[8][18]));
DFFcell _31291_ (.C(clk), .D(_01100_), .Q(cpuregs[8][19]));
DFFcell _31292_ (.C(clk), .D(_01101_), .Q(cpuregs[8][20]));
DFFcell _31293_ (.C(clk), .D(_01102_), .Q(cpuregs[8][21]));
DFFcell _31294_ (.C(clk), .D(_01103_), .Q(cpuregs[8][22]));
DFFcell _31295_ (.C(clk), .D(_01104_), .Q(cpuregs[8][23]));
DFFcell _31296_ (.C(clk), .D(_01105_), .Q(cpuregs[8][24]));
DFFcell _31297_ (.C(clk), .D(_01106_), .Q(cpuregs[8][25]));
DFFcell _31298_ (.C(clk), .D(_01107_), .Q(cpuregs[8][26]));
DFFcell _31299_ (.C(clk), .D(_01108_), .Q(cpuregs[8][27]));
DFFcell _31300_ (.C(clk), .D(_01109_), .Q(cpuregs[8][28]));
DFFcell _31301_ (.C(clk), .D(_01110_), .Q(cpuregs[8][29]));
DFFcell _31302_ (.C(clk), .D(_01111_), .Q(cpuregs[8][30]));
DFFcell _31303_ (.C(clk), .D(_01112_), .Q(cpuregs[8][31]));
DFFcell _31304_ (.C(clk), .D(_01113_), .Q(cpuregs[0][0]));
DFFcell _31305_ (.C(clk), .D(_01114_), .Q(cpuregs[0][1]));
DFFcell _31306_ (.C(clk), .D(_01115_), .Q(cpuregs[0][2]));
DFFcell _31307_ (.C(clk), .D(_01116_), .Q(cpuregs[0][3]));
DFFcell _31308_ (.C(clk), .D(_01117_), .Q(cpuregs[0][4]));
DFFcell _31309_ (.C(clk), .D(_01118_), .Q(cpuregs[0][5]));
DFFcell _31310_ (.C(clk), .D(_01119_), .Q(cpuregs[0][6]));
DFFcell _31311_ (.C(clk), .D(_01120_), .Q(cpuregs[0][7]));
DFFcell _31312_ (.C(clk), .D(_01121_), .Q(cpuregs[0][8]));
DFFcell _31313_ (.C(clk), .D(_01122_), .Q(cpuregs[0][9]));
DFFcell _31314_ (.C(clk), .D(_01123_), .Q(cpuregs[0][10]));
DFFcell _31315_ (.C(clk), .D(_01124_), .Q(cpuregs[0][11]));
DFFcell _31316_ (.C(clk), .D(_01125_), .Q(cpuregs[0][12]));
DFFcell _31317_ (.C(clk), .D(_01126_), .Q(cpuregs[0][13]));
DFFcell _31318_ (.C(clk), .D(_01127_), .Q(cpuregs[0][14]));
DFFcell _31319_ (.C(clk), .D(_01128_), .Q(cpuregs[0][15]));
DFFcell _31320_ (.C(clk), .D(_01129_), .Q(cpuregs[0][16]));
DFFcell _31321_ (.C(clk), .D(_01130_), .Q(cpuregs[0][17]));
DFFcell _31322_ (.C(clk), .D(_01131_), .Q(cpuregs[0][18]));
DFFcell _31323_ (.C(clk), .D(_01132_), .Q(cpuregs[0][19]));
DFFcell _31324_ (.C(clk), .D(_01133_), .Q(cpuregs[0][20]));
DFFcell _31325_ (.C(clk), .D(_01134_), .Q(cpuregs[0][21]));
DFFcell _31326_ (.C(clk), .D(_01135_), .Q(cpuregs[0][22]));
DFFcell _31327_ (.C(clk), .D(_01136_), .Q(cpuregs[0][23]));
DFFcell _31328_ (.C(clk), .D(_01137_), .Q(cpuregs[0][24]));
DFFcell _31329_ (.C(clk), .D(_01138_), .Q(cpuregs[0][25]));
DFFcell _31330_ (.C(clk), .D(_01139_), .Q(cpuregs[0][26]));
DFFcell _31331_ (.C(clk), .D(_01140_), .Q(cpuregs[0][27]));
DFFcell _31332_ (.C(clk), .D(_01141_), .Q(cpuregs[0][28]));
DFFcell _31333_ (.C(clk), .D(_01142_), .Q(cpuregs[0][29]));
DFFcell _31334_ (.C(clk), .D(_01143_), .Q(cpuregs[0][30]));
DFFcell _31335_ (.C(clk), .D(_01144_), .Q(cpuregs[0][31]));
DFFcell _31336_ (.C(clk), .D(_01145_), .Q(decoded_imm_j[8]));
DFFcell _31337_ (.C(clk), .D(_01146_), .Q(decoded_imm_j[9]));
DFFcell _31338_ (.C(clk), .D(_01147_), .Q(cpuregs[26][0]));
DFFcell _31339_ (.C(clk), .D(_01148_), .Q(cpuregs[26][1]));
DFFcell _31340_ (.C(clk), .D(_01149_), .Q(cpuregs[26][2]));
DFFcell _31341_ (.C(clk), .D(_01150_), .Q(cpuregs[26][3]));
DFFcell _31342_ (.C(clk), .D(_01151_), .Q(cpuregs[26][4]));
DFFcell _31343_ (.C(clk), .D(_01152_), .Q(cpuregs[26][5]));
DFFcell _31344_ (.C(clk), .D(_01153_), .Q(cpuregs[26][6]));
DFFcell _31345_ (.C(clk), .D(_01154_), .Q(cpuregs[26][7]));
DFFcell _31346_ (.C(clk), .D(_01155_), .Q(cpuregs[26][8]));
DFFcell _31347_ (.C(clk), .D(_01156_), .Q(cpuregs[26][9]));
DFFcell _31348_ (.C(clk), .D(_01157_), .Q(cpuregs[26][10]));
DFFcell _31349_ (.C(clk), .D(_01158_), .Q(cpuregs[26][11]));
DFFcell _31350_ (.C(clk), .D(_01159_), .Q(cpuregs[26][12]));
DFFcell _31351_ (.C(clk), .D(_01160_), .Q(cpuregs[26][13]));
DFFcell _31352_ (.C(clk), .D(_01161_), .Q(cpuregs[26][14]));
DFFcell _31353_ (.C(clk), .D(_01162_), .Q(cpuregs[26][15]));
DFFcell _31354_ (.C(clk), .D(_01163_), .Q(cpuregs[26][16]));
DFFcell _31355_ (.C(clk), .D(_01164_), .Q(cpuregs[26][17]));
DFFcell _31356_ (.C(clk), .D(_01165_), .Q(cpuregs[26][18]));
DFFcell _31357_ (.C(clk), .D(_01166_), .Q(cpuregs[26][19]));
DFFcell _31358_ (.C(clk), .D(_01167_), .Q(cpuregs[26][20]));
DFFcell _31359_ (.C(clk), .D(_01168_), .Q(cpuregs[26][21]));
DFFcell _31360_ (.C(clk), .D(_01169_), .Q(cpuregs[26][22]));
DFFcell _31361_ (.C(clk), .D(_01170_), .Q(cpuregs[26][23]));
DFFcell _31362_ (.C(clk), .D(_01171_), .Q(cpuregs[26][24]));
DFFcell _31363_ (.C(clk), .D(_01172_), .Q(cpuregs[26][25]));
DFFcell _31364_ (.C(clk), .D(_01173_), .Q(cpuregs[26][26]));
DFFcell _31365_ (.C(clk), .D(_01174_), .Q(cpuregs[26][27]));
DFFcell _31366_ (.C(clk), .D(_01175_), .Q(cpuregs[26][28]));
DFFcell _31367_ (.C(clk), .D(_01176_), .Q(cpuregs[26][29]));
DFFcell _31368_ (.C(clk), .D(_01177_), .Q(cpuregs[26][30]));
DFFcell _31369_ (.C(clk), .D(_01178_), .Q(cpuregs[26][31]));
DFFcell _31370_ (.C(clk), .D(_01179_), .Q(cpuregs[31][0]));
DFFcell _31371_ (.C(clk), .D(_01180_), .Q(cpuregs[31][1]));
DFFcell _31372_ (.C(clk), .D(_01181_), .Q(cpuregs[31][2]));
DFFcell _31373_ (.C(clk), .D(_01182_), .Q(cpuregs[31][3]));
DFFcell _31374_ (.C(clk), .D(_01183_), .Q(cpuregs[31][4]));
DFFcell _31375_ (.C(clk), .D(_01184_), .Q(cpuregs[31][5]));
DFFcell _31376_ (.C(clk), .D(_01185_), .Q(cpuregs[31][6]));
DFFcell _31377_ (.C(clk), .D(_01186_), .Q(cpuregs[31][7]));
DFFcell _31378_ (.C(clk), .D(_01187_), .Q(cpuregs[31][8]));
DFFcell _31379_ (.C(clk), .D(_01188_), .Q(cpuregs[31][9]));
DFFcell _31380_ (.C(clk), .D(_01189_), .Q(cpuregs[31][10]));
DFFcell _31381_ (.C(clk), .D(_01190_), .Q(cpuregs[31][11]));
DFFcell _31382_ (.C(clk), .D(_01191_), .Q(cpuregs[31][12]));
DFFcell _31383_ (.C(clk), .D(_01192_), .Q(cpuregs[31][13]));
DFFcell _31384_ (.C(clk), .D(_01193_), .Q(cpuregs[31][14]));
DFFcell _31385_ (.C(clk), .D(_01194_), .Q(cpuregs[31][15]));
DFFcell _31386_ (.C(clk), .D(_01195_), .Q(cpuregs[31][16]));
DFFcell _31387_ (.C(clk), .D(_01196_), .Q(cpuregs[31][17]));
DFFcell _31388_ (.C(clk), .D(_01197_), .Q(cpuregs[31][18]));
DFFcell _31389_ (.C(clk), .D(_01198_), .Q(cpuregs[31][19]));
DFFcell _31390_ (.C(clk), .D(_01199_), .Q(cpuregs[31][20]));
DFFcell _31391_ (.C(clk), .D(_01200_), .Q(cpuregs[31][21]));
DFFcell _31392_ (.C(clk), .D(_01201_), .Q(cpuregs[31][22]));
DFFcell _31393_ (.C(clk), .D(_01202_), .Q(cpuregs[31][23]));
DFFcell _31394_ (.C(clk), .D(_01203_), .Q(cpuregs[31][24]));
DFFcell _31395_ (.C(clk), .D(_01204_), .Q(cpuregs[31][25]));
DFFcell _31396_ (.C(clk), .D(_01205_), .Q(cpuregs[31][26]));
DFFcell _31397_ (.C(clk), .D(_01206_), .Q(cpuregs[31][27]));
DFFcell _31398_ (.C(clk), .D(_01207_), .Q(cpuregs[31][28]));
DFFcell _31399_ (.C(clk), .D(_01208_), .Q(cpuregs[31][29]));
DFFcell _31400_ (.C(clk), .D(_01209_), .Q(cpuregs[31][30]));
DFFcell _31401_ (.C(clk), .D(_01210_), .Q(cpuregs[31][31]));
DFFcell _31402_ (.C(clk), .D(_01211_), .Q(cpuregs[19][0]));
DFFcell _31403_ (.C(clk), .D(_01212_), .Q(cpuregs[19][1]));
DFFcell _31404_ (.C(clk), .D(_01213_), .Q(cpuregs[19][2]));
DFFcell _31405_ (.C(clk), .D(_01214_), .Q(cpuregs[19][3]));
DFFcell _31406_ (.C(clk), .D(_01215_), .Q(cpuregs[19][4]));
DFFcell _31407_ (.C(clk), .D(_01216_), .Q(cpuregs[19][5]));
DFFcell _31408_ (.C(clk), .D(_01217_), .Q(cpuregs[19][6]));
DFFcell _31409_ (.C(clk), .D(_01218_), .Q(cpuregs[19][7]));
DFFcell _31410_ (.C(clk), .D(_01219_), .Q(cpuregs[19][8]));
DFFcell _31411_ (.C(clk), .D(_01220_), .Q(cpuregs[19][9]));
DFFcell _31412_ (.C(clk), .D(_01221_), .Q(cpuregs[19][10]));
DFFcell _31413_ (.C(clk), .D(_01222_), .Q(cpuregs[19][11]));
DFFcell _31414_ (.C(clk), .D(_01223_), .Q(cpuregs[19][12]));
DFFcell _31415_ (.C(clk), .D(_01224_), .Q(cpuregs[19][13]));
DFFcell _31416_ (.C(clk), .D(_01225_), .Q(cpuregs[19][14]));
DFFcell _31417_ (.C(clk), .D(_01226_), .Q(cpuregs[19][15]));
DFFcell _31418_ (.C(clk), .D(_01227_), .Q(cpuregs[19][16]));
DFFcell _31419_ (.C(clk), .D(_01228_), .Q(cpuregs[19][17]));
DFFcell _31420_ (.C(clk), .D(_01229_), .Q(cpuregs[19][18]));
DFFcell _31421_ (.C(clk), .D(_01230_), .Q(cpuregs[19][19]));
DFFcell _31422_ (.C(clk), .D(_01231_), .Q(cpuregs[19][20]));
DFFcell _31423_ (.C(clk), .D(_01232_), .Q(cpuregs[19][21]));
DFFcell _31424_ (.C(clk), .D(_01233_), .Q(cpuregs[19][22]));
DFFcell _31425_ (.C(clk), .D(_01234_), .Q(cpuregs[19][23]));
DFFcell _31426_ (.C(clk), .D(_01235_), .Q(cpuregs[19][24]));
DFFcell _31427_ (.C(clk), .D(_01236_), .Q(cpuregs[19][25]));
DFFcell _31428_ (.C(clk), .D(_01237_), .Q(cpuregs[19][26]));
DFFcell _31429_ (.C(clk), .D(_01238_), .Q(cpuregs[19][27]));
DFFcell _31430_ (.C(clk), .D(_01239_), .Q(cpuregs[19][28]));
DFFcell _31431_ (.C(clk), .D(_01240_), .Q(cpuregs[19][29]));
DFFcell _31432_ (.C(clk), .D(_01241_), .Q(cpuregs[19][30]));
DFFcell _31433_ (.C(clk), .D(_01242_), .Q(cpuregs[19][31]));
DFFcell _31434_ (.C(clk), .D(_01243_), .Q(decoded_imm_j[6]));
DFFcell _31435_ (.C(clk), .D(_01244_), .Q(cpuregs[25][0]));
DFFcell _31436_ (.C(clk), .D(_01245_), .Q(cpuregs[25][1]));
DFFcell _31437_ (.C(clk), .D(_01246_), .Q(cpuregs[25][2]));
DFFcell _31438_ (.C(clk), .D(_01247_), .Q(cpuregs[25][3]));
DFFcell _31439_ (.C(clk), .D(_01248_), .Q(cpuregs[25][4]));
DFFcell _31440_ (.C(clk), .D(_01249_), .Q(cpuregs[25][5]));
DFFcell _31441_ (.C(clk), .D(_01250_), .Q(cpuregs[25][6]));
DFFcell _31442_ (.C(clk), .D(_01251_), .Q(cpuregs[25][7]));
DFFcell _31443_ (.C(clk), .D(_01252_), .Q(cpuregs[25][8]));
DFFcell _31444_ (.C(clk), .D(_01253_), .Q(cpuregs[25][9]));
DFFcell _31445_ (.C(clk), .D(_01254_), .Q(cpuregs[25][10]));
DFFcell _31446_ (.C(clk), .D(_01255_), .Q(cpuregs[25][11]));
DFFcell _31447_ (.C(clk), .D(_01256_), .Q(cpuregs[25][12]));
DFFcell _31448_ (.C(clk), .D(_01257_), .Q(cpuregs[25][13]));
DFFcell _31449_ (.C(clk), .D(_01258_), .Q(cpuregs[25][14]));
DFFcell _31450_ (.C(clk), .D(_01259_), .Q(cpuregs[25][15]));
DFFcell _31451_ (.C(clk), .D(_01260_), .Q(cpuregs[25][16]));
DFFcell _31452_ (.C(clk), .D(_01261_), .Q(cpuregs[25][17]));
DFFcell _31453_ (.C(clk), .D(_01262_), .Q(cpuregs[25][18]));
DFFcell _31454_ (.C(clk), .D(_01263_), .Q(cpuregs[25][19]));
DFFcell _31455_ (.C(clk), .D(_01264_), .Q(cpuregs[25][20]));
DFFcell _31456_ (.C(clk), .D(_01265_), .Q(cpuregs[25][21]));
DFFcell _31457_ (.C(clk), .D(_01266_), .Q(cpuregs[25][22]));
DFFcell _31458_ (.C(clk), .D(_01267_), .Q(cpuregs[25][23]));
DFFcell _31459_ (.C(clk), .D(_01268_), .Q(cpuregs[25][24]));
DFFcell _31460_ (.C(clk), .D(_01269_), .Q(cpuregs[25][25]));
DFFcell _31461_ (.C(clk), .D(_01270_), .Q(cpuregs[25][26]));
DFFcell _31462_ (.C(clk), .D(_01271_), .Q(cpuregs[25][27]));
DFFcell _31463_ (.C(clk), .D(_01272_), .Q(cpuregs[25][28]));
DFFcell _31464_ (.C(clk), .D(_01273_), .Q(cpuregs[25][29]));
DFFcell _31465_ (.C(clk), .D(_01274_), .Q(cpuregs[25][30]));
DFFcell _31466_ (.C(clk), .D(_01275_), .Q(cpuregs[25][31]));
DFFcell _31467_ (.C(clk), .D(_01276_), .Q(cpuregs[9][0]));
DFFcell _31468_ (.C(clk), .D(_01277_), .Q(cpuregs[9][1]));
DFFcell _31469_ (.C(clk), .D(_01278_), .Q(cpuregs[9][2]));
DFFcell _31470_ (.C(clk), .D(_01279_), .Q(cpuregs[9][3]));
DFFcell _31471_ (.C(clk), .D(_01280_), .Q(cpuregs[9][4]));
DFFcell _31472_ (.C(clk), .D(_01281_), .Q(cpuregs[9][5]));
DFFcell _31473_ (.C(clk), .D(_01282_), .Q(cpuregs[9][6]));
DFFcell _31474_ (.C(clk), .D(_01283_), .Q(cpuregs[9][7]));
DFFcell _31475_ (.C(clk), .D(_01284_), .Q(cpuregs[9][8]));
DFFcell _31476_ (.C(clk), .D(_01285_), .Q(cpuregs[9][9]));
DFFcell _31477_ (.C(clk), .D(_01286_), .Q(cpuregs[9][10]));
DFFcell _31478_ (.C(clk), .D(_01287_), .Q(cpuregs[9][11]));
DFFcell _31479_ (.C(clk), .D(_01288_), .Q(cpuregs[9][12]));
DFFcell _31480_ (.C(clk), .D(_01289_), .Q(cpuregs[9][13]));
DFFcell _31481_ (.C(clk), .D(_01290_), .Q(cpuregs[9][14]));
DFFcell _31482_ (.C(clk), .D(_01291_), .Q(cpuregs[9][15]));
DFFcell _31483_ (.C(clk), .D(_01292_), .Q(cpuregs[9][16]));
DFFcell _31484_ (.C(clk), .D(_01293_), .Q(cpuregs[9][17]));
DFFcell _31485_ (.C(clk), .D(_01294_), .Q(cpuregs[9][18]));
DFFcell _31486_ (.C(clk), .D(_01295_), .Q(cpuregs[9][19]));
DFFcell _31487_ (.C(clk), .D(_01296_), .Q(cpuregs[9][20]));
DFFcell _31488_ (.C(clk), .D(_01297_), .Q(cpuregs[9][21]));
DFFcell _31489_ (.C(clk), .D(_01298_), .Q(cpuregs[9][22]));
DFFcell _31490_ (.C(clk), .D(_01299_), .Q(cpuregs[9][23]));
DFFcell _31491_ (.C(clk), .D(_01300_), .Q(cpuregs[9][24]));
DFFcell _31492_ (.C(clk), .D(_01301_), .Q(cpuregs[9][25]));
DFFcell _31493_ (.C(clk), .D(_01302_), .Q(cpuregs[9][26]));
DFFcell _31494_ (.C(clk), .D(_01303_), .Q(cpuregs[9][27]));
DFFcell _31495_ (.C(clk), .D(_01304_), .Q(cpuregs[9][28]));
DFFcell _31496_ (.C(clk), .D(_01305_), .Q(cpuregs[9][29]));
DFFcell _31497_ (.C(clk), .D(_01306_), .Q(cpuregs[9][30]));
DFFcell _31498_ (.C(clk), .D(_01307_), .Q(cpuregs[9][31]));
DFFcell _31499_ (.C(clk), .D(_01308_), .Q(cpuregs[21][0]));
DFFcell _31500_ (.C(clk), .D(_01309_), .Q(cpuregs[21][1]));
DFFcell _31501_ (.C(clk), .D(_01310_), .Q(cpuregs[21][2]));
DFFcell _31502_ (.C(clk), .D(_01311_), .Q(cpuregs[21][3]));
DFFcell _31503_ (.C(clk), .D(_01312_), .Q(cpuregs[21][4]));
DFFcell _31504_ (.C(clk), .D(_01313_), .Q(cpuregs[21][5]));
DFFcell _31505_ (.C(clk), .D(_01314_), .Q(cpuregs[21][6]));
DFFcell _31506_ (.C(clk), .D(_01315_), .Q(cpuregs[21][7]));
DFFcell _31507_ (.C(clk), .D(_01316_), .Q(cpuregs[21][8]));
DFFcell _31508_ (.C(clk), .D(_01317_), .Q(cpuregs[21][9]));
DFFcell _31509_ (.C(clk), .D(_01318_), .Q(cpuregs[21][10]));
DFFcell _31510_ (.C(clk), .D(_01319_), .Q(cpuregs[21][11]));
DFFcell _31511_ (.C(clk), .D(_01320_), .Q(cpuregs[21][12]));
DFFcell _31512_ (.C(clk), .D(_01321_), .Q(cpuregs[21][13]));
DFFcell _31513_ (.C(clk), .D(_01322_), .Q(cpuregs[21][14]));
DFFcell _31514_ (.C(clk), .D(_01323_), .Q(cpuregs[21][15]));
DFFcell _31515_ (.C(clk), .D(_01324_), .Q(cpuregs[21][16]));
DFFcell _31516_ (.C(clk), .D(_01325_), .Q(cpuregs[21][17]));
DFFcell _31517_ (.C(clk), .D(_01326_), .Q(cpuregs[21][18]));
DFFcell _31518_ (.C(clk), .D(_01327_), .Q(cpuregs[21][19]));
DFFcell _31519_ (.C(clk), .D(_01328_), .Q(cpuregs[21][20]));
DFFcell _31520_ (.C(clk), .D(_01329_), .Q(cpuregs[21][21]));
DFFcell _31521_ (.C(clk), .D(_01330_), .Q(cpuregs[21][22]));
DFFcell _31522_ (.C(clk), .D(_01331_), .Q(cpuregs[21][23]));
DFFcell _31523_ (.C(clk), .D(_01332_), .Q(cpuregs[21][24]));
DFFcell _31524_ (.C(clk), .D(_01333_), .Q(cpuregs[21][25]));
DFFcell _31525_ (.C(clk), .D(_01334_), .Q(cpuregs[21][26]));
DFFcell _31526_ (.C(clk), .D(_01335_), .Q(cpuregs[21][27]));
DFFcell _31527_ (.C(clk), .D(_01336_), .Q(cpuregs[21][28]));
DFFcell _31528_ (.C(clk), .D(_01337_), .Q(cpuregs[21][29]));
DFFcell _31529_ (.C(clk), .D(_01338_), .Q(cpuregs[21][30]));
DFFcell _31530_ (.C(clk), .D(_01339_), .Q(cpuregs[21][31]));
DFFcell _31531_ (.C(clk), .D(_01340_), .Q(cpuregs[6][0]));
DFFcell _31532_ (.C(clk), .D(_01341_), .Q(cpuregs[6][1]));
DFFcell _31533_ (.C(clk), .D(_01342_), .Q(cpuregs[6][2]));
DFFcell _31534_ (.C(clk), .D(_01343_), .Q(cpuregs[6][3]));
DFFcell _31535_ (.C(clk), .D(_01344_), .Q(cpuregs[6][4]));
DFFcell _31536_ (.C(clk), .D(_01345_), .Q(cpuregs[6][5]));
DFFcell _31537_ (.C(clk), .D(_01346_), .Q(cpuregs[6][6]));
DFFcell _31538_ (.C(clk), .D(_01347_), .Q(cpuregs[6][7]));
DFFcell _31539_ (.C(clk), .D(_01348_), .Q(cpuregs[6][8]));
DFFcell _31540_ (.C(clk), .D(_01349_), .Q(cpuregs[6][9]));
DFFcell _31541_ (.C(clk), .D(_01350_), .Q(cpuregs[6][10]));
DFFcell _31542_ (.C(clk), .D(_01351_), .Q(cpuregs[6][11]));
DFFcell _31543_ (.C(clk), .D(_01352_), .Q(cpuregs[6][12]));
DFFcell _31544_ (.C(clk), .D(_01353_), .Q(cpuregs[6][13]));
DFFcell _31545_ (.C(clk), .D(_01354_), .Q(cpuregs[6][14]));
DFFcell _31546_ (.C(clk), .D(_01355_), .Q(cpuregs[6][15]));
DFFcell _31547_ (.C(clk), .D(_01356_), .Q(cpuregs[6][16]));
DFFcell _31548_ (.C(clk), .D(_01357_), .Q(cpuregs[6][17]));
DFFcell _31549_ (.C(clk), .D(_01358_), .Q(cpuregs[6][18]));
DFFcell _31550_ (.C(clk), .D(_01359_), .Q(cpuregs[6][19]));
DFFcell _31551_ (.C(clk), .D(_01360_), .Q(cpuregs[6][20]));
DFFcell _31552_ (.C(clk), .D(_01361_), .Q(cpuregs[6][21]));
DFFcell _31553_ (.C(clk), .D(_01362_), .Q(cpuregs[6][22]));
DFFcell _31554_ (.C(clk), .D(_01363_), .Q(cpuregs[6][23]));
DFFcell _31555_ (.C(clk), .D(_01364_), .Q(cpuregs[6][24]));
DFFcell _31556_ (.C(clk), .D(_01365_), .Q(cpuregs[6][25]));
DFFcell _31557_ (.C(clk), .D(_01366_), .Q(cpuregs[6][26]));
DFFcell _31558_ (.C(clk), .D(_01367_), .Q(cpuregs[6][27]));
DFFcell _31559_ (.C(clk), .D(_01368_), .Q(cpuregs[6][28]));
DFFcell _31560_ (.C(clk), .D(_01369_), .Q(cpuregs[6][29]));
DFFcell _31561_ (.C(clk), .D(_01370_), .Q(cpuregs[6][30]));
DFFcell _31562_ (.C(clk), .D(_01371_), .Q(cpuregs[6][31]));
DFFcell _31563_ (.C(clk), .D(_01372_), .Q(cpuregs[10][0]));
DFFcell _31564_ (.C(clk), .D(_01373_), .Q(cpuregs[10][1]));
DFFcell _31565_ (.C(clk), .D(_01374_), .Q(cpuregs[10][2]));
DFFcell _31566_ (.C(clk), .D(_01375_), .Q(cpuregs[10][3]));
DFFcell _31567_ (.C(clk), .D(_01376_), .Q(cpuregs[10][4]));
DFFcell _31568_ (.C(clk), .D(_01377_), .Q(cpuregs[10][5]));
DFFcell _31569_ (.C(clk), .D(_01378_), .Q(cpuregs[10][6]));
DFFcell _31570_ (.C(clk), .D(_01379_), .Q(cpuregs[10][7]));
DFFcell _31571_ (.C(clk), .D(_01380_), .Q(cpuregs[10][8]));
DFFcell _31572_ (.C(clk), .D(_01381_), .Q(cpuregs[10][9]));
DFFcell _31573_ (.C(clk), .D(_01382_), .Q(cpuregs[10][10]));
DFFcell _31574_ (.C(clk), .D(_01383_), .Q(cpuregs[10][11]));
DFFcell _31575_ (.C(clk), .D(_01384_), .Q(cpuregs[10][12]));
DFFcell _31576_ (.C(clk), .D(_01385_), .Q(cpuregs[10][13]));
DFFcell _31577_ (.C(clk), .D(_01386_), .Q(cpuregs[10][14]));
DFFcell _31578_ (.C(clk), .D(_01387_), .Q(cpuregs[10][15]));
DFFcell _31579_ (.C(clk), .D(_01388_), .Q(cpuregs[10][16]));
DFFcell _31580_ (.C(clk), .D(_01389_), .Q(cpuregs[10][17]));
DFFcell _31581_ (.C(clk), .D(_01390_), .Q(cpuregs[10][18]));
DFFcell _31582_ (.C(clk), .D(_01391_), .Q(cpuregs[10][19]));
DFFcell _31583_ (.C(clk), .D(_01392_), .Q(cpuregs[10][20]));
DFFcell _31584_ (.C(clk), .D(_01393_), .Q(cpuregs[10][21]));
DFFcell _31585_ (.C(clk), .D(_01394_), .Q(cpuregs[10][22]));
DFFcell _31586_ (.C(clk), .D(_01395_), .Q(cpuregs[10][23]));
DFFcell _31587_ (.C(clk), .D(_01396_), .Q(cpuregs[10][24]));
DFFcell _31588_ (.C(clk), .D(_01397_), .Q(cpuregs[10][25]));
DFFcell _31589_ (.C(clk), .D(_01398_), .Q(cpuregs[10][26]));
DFFcell _31590_ (.C(clk), .D(_01399_), .Q(cpuregs[10][27]));
DFFcell _31591_ (.C(clk), .D(_01400_), .Q(cpuregs[10][28]));
DFFcell _31592_ (.C(clk), .D(_01401_), .Q(cpuregs[10][29]));
DFFcell _31593_ (.C(clk), .D(_01402_), .Q(cpuregs[10][30]));
DFFcell _31594_ (.C(clk), .D(_01403_), .Q(cpuregs[10][31]));
DFFcell _31595_ (.C(clk), .D(_01404_), .Q(cpuregs[24][0]));
DFFcell _31596_ (.C(clk), .D(_01405_), .Q(cpuregs[24][1]));
DFFcell _31597_ (.C(clk), .D(_01406_), .Q(cpuregs[24][2]));
DFFcell _31598_ (.C(clk), .D(_01407_), .Q(cpuregs[24][3]));
DFFcell _31599_ (.C(clk), .D(_01408_), .Q(cpuregs[24][4]));
DFFcell _31600_ (.C(clk), .D(_01409_), .Q(cpuregs[24][5]));
DFFcell _31601_ (.C(clk), .D(_01410_), .Q(cpuregs[24][6]));
DFFcell _31602_ (.C(clk), .D(_01411_), .Q(cpuregs[24][7]));
DFFcell _31603_ (.C(clk), .D(_01412_), .Q(cpuregs[24][8]));
DFFcell _31604_ (.C(clk), .D(_01413_), .Q(cpuregs[24][9]));
DFFcell _31605_ (.C(clk), .D(_01414_), .Q(cpuregs[24][10]));
DFFcell _31606_ (.C(clk), .D(_01415_), .Q(cpuregs[24][11]));
DFFcell _31607_ (.C(clk), .D(_01416_), .Q(cpuregs[24][12]));
DFFcell _31608_ (.C(clk), .D(_01417_), .Q(cpuregs[24][13]));
DFFcell _31609_ (.C(clk), .D(_01418_), .Q(cpuregs[24][14]));
DFFcell _31610_ (.C(clk), .D(_01419_), .Q(cpuregs[24][15]));
DFFcell _31611_ (.C(clk), .D(_01420_), .Q(cpuregs[24][16]));
DFFcell _31612_ (.C(clk), .D(_01421_), .Q(cpuregs[24][17]));
DFFcell _31613_ (.C(clk), .D(_01422_), .Q(cpuregs[24][18]));
DFFcell _31614_ (.C(clk), .D(_01423_), .Q(cpuregs[24][19]));
DFFcell _31615_ (.C(clk), .D(_01424_), .Q(cpuregs[24][20]));
DFFcell _31616_ (.C(clk), .D(_01425_), .Q(cpuregs[24][21]));
DFFcell _31617_ (.C(clk), .D(_01426_), .Q(cpuregs[24][22]));
DFFcell _31618_ (.C(clk), .D(_01427_), .Q(cpuregs[24][23]));
DFFcell _31619_ (.C(clk), .D(_01428_), .Q(cpuregs[24][24]));
DFFcell _31620_ (.C(clk), .D(_01429_), .Q(cpuregs[24][25]));
DFFcell _31621_ (.C(clk), .D(_01430_), .Q(cpuregs[24][26]));
DFFcell _31622_ (.C(clk), .D(_01431_), .Q(cpuregs[24][27]));
DFFcell _31623_ (.C(clk), .D(_01432_), .Q(cpuregs[24][28]));
DFFcell _31624_ (.C(clk), .D(_01433_), .Q(cpuregs[24][29]));
DFFcell _31625_ (.C(clk), .D(_01434_), .Q(cpuregs[24][30]));
DFFcell _31626_ (.C(clk), .D(_01435_), .Q(cpuregs[24][31]));
DFFcell _31627_ (.C(clk), .D(_01436_), .Q(decoded_imm_j[31]));
DFFcell _31628_ (.C(clk), .D(_01437_), .Q(decoded_imm_j[5]));
DFFcell _31629_ (.C(clk), .D(_01438_), .Q(decoded_imm_j[7]));
DFFcell _31630_ (.C(clk), .D(_01439_), .Q(cpuregs[16][0]));
DFFcell _31631_ (.C(clk), .D(_01440_), .Q(cpuregs[16][1]));
DFFcell _31632_ (.C(clk), .D(_01441_), .Q(cpuregs[16][2]));
DFFcell _31633_ (.C(clk), .D(_01442_), .Q(cpuregs[16][3]));
DFFcell _31634_ (.C(clk), .D(_01443_), .Q(cpuregs[16][4]));
DFFcell _31635_ (.C(clk), .D(_01444_), .Q(cpuregs[16][5]));
DFFcell _31636_ (.C(clk), .D(_01445_), .Q(cpuregs[16][6]));
DFFcell _31637_ (.C(clk), .D(_01446_), .Q(cpuregs[16][7]));
DFFcell _31638_ (.C(clk), .D(_01447_), .Q(cpuregs[16][8]));
DFFcell _31639_ (.C(clk), .D(_01448_), .Q(cpuregs[16][9]));
DFFcell _31640_ (.C(clk), .D(_01449_), .Q(cpuregs[16][10]));
DFFcell _31641_ (.C(clk), .D(_01450_), .Q(cpuregs[16][11]));
DFFcell _31642_ (.C(clk), .D(_01451_), .Q(cpuregs[16][12]));
DFFcell _31643_ (.C(clk), .D(_01452_), .Q(cpuregs[16][13]));
DFFcell _31644_ (.C(clk), .D(_01453_), .Q(cpuregs[16][14]));
DFFcell _31645_ (.C(clk), .D(_01454_), .Q(cpuregs[16][15]));
DFFcell _31646_ (.C(clk), .D(_01455_), .Q(cpuregs[16][16]));
DFFcell _31647_ (.C(clk), .D(_01456_), .Q(cpuregs[16][17]));
DFFcell _31648_ (.C(clk), .D(_01457_), .Q(cpuregs[16][18]));
DFFcell _31649_ (.C(clk), .D(_01458_), .Q(cpuregs[16][19]));
DFFcell _31650_ (.C(clk), .D(_01459_), .Q(cpuregs[16][20]));
DFFcell _31651_ (.C(clk), .D(_01460_), .Q(cpuregs[16][21]));
DFFcell _31652_ (.C(clk), .D(_01461_), .Q(cpuregs[16][22]));
DFFcell _31653_ (.C(clk), .D(_01462_), .Q(cpuregs[16][23]));
DFFcell _31654_ (.C(clk), .D(_01463_), .Q(cpuregs[16][24]));
DFFcell _31655_ (.C(clk), .D(_01464_), .Q(cpuregs[16][25]));
DFFcell _31656_ (.C(clk), .D(_01465_), .Q(cpuregs[16][26]));
DFFcell _31657_ (.C(clk), .D(_01466_), .Q(cpuregs[16][27]));
DFFcell _31658_ (.C(clk), .D(_01467_), .Q(cpuregs[16][28]));
DFFcell _31659_ (.C(clk), .D(_01468_), .Q(cpuregs[16][29]));
DFFcell _31660_ (.C(clk), .D(_01469_), .Q(cpuregs[16][30]));
DFFcell _31661_ (.C(clk), .D(_01470_), .Q(cpuregs[16][31]));
DFFcell _31662_ (.C(clk), .D(_01471_), .Q(cpuregs[27][0]));
DFFcell _31663_ (.C(clk), .D(_01472_), .Q(cpuregs[27][1]));
DFFcell _31664_ (.C(clk), .D(_01473_), .Q(cpuregs[27][2]));
DFFcell _31665_ (.C(clk), .D(_01474_), .Q(cpuregs[27][3]));
DFFcell _31666_ (.C(clk), .D(_01475_), .Q(cpuregs[27][4]));
DFFcell _31667_ (.C(clk), .D(_01476_), .Q(cpuregs[27][5]));
DFFcell _31668_ (.C(clk), .D(_01477_), .Q(cpuregs[27][6]));
DFFcell _31669_ (.C(clk), .D(_01478_), .Q(cpuregs[27][7]));
DFFcell _31670_ (.C(clk), .D(_01479_), .Q(cpuregs[27][8]));
DFFcell _31671_ (.C(clk), .D(_01480_), .Q(cpuregs[27][9]));
DFFcell _31672_ (.C(clk), .D(_01481_), .Q(cpuregs[27][10]));
DFFcell _31673_ (.C(clk), .D(_01482_), .Q(cpuregs[27][11]));
DFFcell _31674_ (.C(clk), .D(_01483_), .Q(cpuregs[27][12]));
DFFcell _31675_ (.C(clk), .D(_01484_), .Q(cpuregs[27][13]));
DFFcell _31676_ (.C(clk), .D(_01485_), .Q(cpuregs[27][14]));
DFFcell _31677_ (.C(clk), .D(_01486_), .Q(cpuregs[27][15]));
DFFcell _31678_ (.C(clk), .D(_01487_), .Q(cpuregs[27][16]));
DFFcell _31679_ (.C(clk), .D(_01488_), .Q(cpuregs[27][17]));
DFFcell _31680_ (.C(clk), .D(_01489_), .Q(cpuregs[27][18]));
DFFcell _31681_ (.C(clk), .D(_01490_), .Q(cpuregs[27][19]));
DFFcell _31682_ (.C(clk), .D(_01491_), .Q(cpuregs[27][20]));
DFFcell _31683_ (.C(clk), .D(_01492_), .Q(cpuregs[27][21]));
DFFcell _31684_ (.C(clk), .D(_01493_), .Q(cpuregs[27][22]));
DFFcell _31685_ (.C(clk), .D(_01494_), .Q(cpuregs[27][23]));
DFFcell _31686_ (.C(clk), .D(_01495_), .Q(cpuregs[27][24]));
DFFcell _31687_ (.C(clk), .D(_01496_), .Q(cpuregs[27][25]));
DFFcell _31688_ (.C(clk), .D(_01497_), .Q(cpuregs[27][26]));
DFFcell _31689_ (.C(clk), .D(_01498_), .Q(cpuregs[27][27]));
DFFcell _31690_ (.C(clk), .D(_01499_), .Q(cpuregs[27][28]));
DFFcell _31691_ (.C(clk), .D(_01500_), .Q(cpuregs[27][29]));
DFFcell _31692_ (.C(clk), .D(_01501_), .Q(cpuregs[27][30]));
DFFcell _31693_ (.C(clk), .D(_01502_), .Q(cpuregs[27][31]));
DFFcell _31694_ (.C(clk), .D(_01503_), .Q(cpuregs[28][0]));
DFFcell _31695_ (.C(clk), .D(_01504_), .Q(cpuregs[28][1]));
DFFcell _31696_ (.C(clk), .D(_01505_), .Q(cpuregs[28][2]));
DFFcell _31697_ (.C(clk), .D(_01506_), .Q(cpuregs[28][3]));
DFFcell _31698_ (.C(clk), .D(_01507_), .Q(cpuregs[28][4]));
DFFcell _31699_ (.C(clk), .D(_01508_), .Q(cpuregs[28][5]));
DFFcell _31700_ (.C(clk), .D(_01509_), .Q(cpuregs[28][6]));
DFFcell _31701_ (.C(clk), .D(_01510_), .Q(cpuregs[28][7]));
DFFcell _31702_ (.C(clk), .D(_01511_), .Q(cpuregs[28][8]));
DFFcell _31703_ (.C(clk), .D(_01512_), .Q(cpuregs[28][9]));
DFFcell _31704_ (.C(clk), .D(_01513_), .Q(cpuregs[28][10]));
DFFcell _31705_ (.C(clk), .D(_01514_), .Q(cpuregs[28][11]));
DFFcell _31706_ (.C(clk), .D(_01515_), .Q(cpuregs[28][12]));
DFFcell _31707_ (.C(clk), .D(_01516_), .Q(cpuregs[28][13]));
DFFcell _31708_ (.C(clk), .D(_01517_), .Q(cpuregs[28][14]));
DFFcell _31709_ (.C(clk), .D(_01518_), .Q(cpuregs[28][15]));
DFFcell _31710_ (.C(clk), .D(_01519_), .Q(cpuregs[28][16]));
DFFcell _31711_ (.C(clk), .D(_01520_), .Q(cpuregs[28][17]));
DFFcell _31712_ (.C(clk), .D(_01521_), .Q(cpuregs[28][18]));
DFFcell _31713_ (.C(clk), .D(_01522_), .Q(cpuregs[28][19]));
DFFcell _31714_ (.C(clk), .D(_01523_), .Q(cpuregs[28][20]));
DFFcell _31715_ (.C(clk), .D(_01524_), .Q(cpuregs[28][21]));
DFFcell _31716_ (.C(clk), .D(_01525_), .Q(cpuregs[28][22]));
DFFcell _31717_ (.C(clk), .D(_01526_), .Q(cpuregs[28][23]));
DFFcell _31718_ (.C(clk), .D(_01527_), .Q(cpuregs[28][24]));
DFFcell _31719_ (.C(clk), .D(_01528_), .Q(cpuregs[28][25]));
DFFcell _31720_ (.C(clk), .D(_01529_), .Q(cpuregs[28][26]));
DFFcell _31721_ (.C(clk), .D(_01530_), .Q(cpuregs[28][27]));
DFFcell _31722_ (.C(clk), .D(_01531_), .Q(cpuregs[28][28]));
DFFcell _31723_ (.C(clk), .D(_01532_), .Q(cpuregs[28][29]));
DFFcell _31724_ (.C(clk), .D(_01533_), .Q(cpuregs[28][30]));
DFFcell _31725_ (.C(clk), .D(_01534_), .Q(cpuregs[28][31]));
DFFcell _31726_ (.C(clk), .D(_00014_), .Q(_00008_[0]));
DFFcell _31727_ (.C(clk), .D(_00015_), .Q(_00008_[1]));
DFFcell _31728_ (.C(clk), .D(_00016_), .Q(_00008_[2]));
DFFcell _31729_ (.C(clk), .D(_00017_), .Q(_00008_[3]));
DFFcell _31730_ (.C(clk), .D(_00018_), .Q(_00008_[4]));
assign { decoded_imm_j[30:20], decoded_imm_j[0] } = { decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], decoded_imm_j[31], 1'h0 };
assign eoi = 32'd0;
assign mem_addr[1:0] = 2'h0;
assign mem_la_addr[1:0] = 2'h0;
assign pcpi_insn = 32'hxxxxxxxx;
assign pcpi_valid = 1'h0;
assign reg_pc[0] = reg_next_pc[0];
assign trace_data = 36'hxxxxxxxxx;
assign trace_valid = 1'h0;
endmodule
