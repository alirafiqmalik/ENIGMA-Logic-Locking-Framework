module top(inputs,key,Q,Z);
input [7:0] inputs;
input [7:0] key;
wire [1:0] out_enc, out_org;
orgcir org(.inputs(inputs),.key(key),.out(out_org));
enccir enc(.inputs(inputs),.key(key),.out(out_enc));
output Z;
output [1:0]Q;
assign Q[0]=out_enc[0]==out_org[0];
assign Q[1]=out_enc[1]==out_org[1];
assign Z= Q[0]&Q[1];
endmodule



module enccir(inputs,key,out);
input [7:0] inputs;
input [7:0] key;
output [1:0] out;
wire _060_;
wire _015_;
wire _069_;
wire _009_;
wire [4:0] s.c.c;
wire _058_;
wire _055_;
wire _046_;
wire _057_;
wire _030_;
wire [4:0] s1.c.c;
wire _035_;
wire _023_;
wire _048_;
wire _059_;
wire _021_;
wire _043_;
wire _028_;
wire _062_;
wire _010_;
wire _025_;
wire _044_;
wire _018_;
wire _063_;
wire _033_;
wire _051_;
wire _029_;
wire _038_;
wire _020_;
wire _027_;
wire _016_;
wire _041_;
wire _070_;
wire _054_;
wire _065_;
wire _017_;
wire _011_;
wire _014_;
wire _000_;
wire _034_;
wire _071_;
wire _031_;
wire _042_;
wire _052_;
wire _004_;
wire _067_;
wire _002_;
wire _061_;
wire _032_;
wire _006_;
wire _012_;
wire _022_;
wire _007_;
wire _056_;
wire _003_;
wire _024_;
wire _045_;
wire _049_;
wire _013_;
wire _047_;
wire _050_;
wire _019_;
wire _036_;
wire _008_;
wire _066_;
wire _037_;
wire _068_;
wire _040_;
wire _039_;
wire _005_;
wire _001_;
wire _064_;
wire _053_;
wire _026_;
NOT_g NOT_g_072_(.A(inputs[3]), .Y(_000_));
NOT_g NOT_g_114_(.A(inputs[3]), .Y(_036_));
XNOR_g XNOR_g_073_(.A(key[0]), .B(inputs[0]), .Y(_001_));
XNOR_g XNOR_g_074_(.A(key[7]), .B(inputs[7]), .Y(_002_));
XNOR_g XNOR_g_076_(.A(key[1]), .B(inputs[1]), .Y(_004_));
XNOR_g XNOR_g_077_(.A(key[3]), .B(inputs[3]), .Y(_005_));
XNOR_g XNOR_g_087_(.A(key[5]), .B(inputs[5]), .Y(_015_));
XNOR_g XNOR_g_088_(.A(key[2]), .B(inputs[2]), .Y(_016_));
XNOR_g XNOR_g_090_(.A(key[6]), .B(inputs[6]), .Y(_018_));
XNOR_g XNOR_g_091_(.A(key[4]), .B(inputs[4]), .Y(_019_));
XNOR_g XNOR_g_096_(.A(_023_), .B(s.c.c[0]), .Y(out[0]));
XNOR_g XNOR_g_115_(.A(key[0]), .B(inputs[0]), .Y(_037_));
XNOR_g XNOR_g_116_(.A(key[7]), .B(inputs[7]), .Y(_038_));
XNOR_g XNOR_g_118_(.A(key[1]), .B(inputs[1]), .Y(_040_));
XNOR_g XNOR_g_119_(.A(key[3]), .B(inputs[3]), .Y(_041_));
XNOR_g XNOR_g_129_(.A(key[5]), .B(inputs[5]), .Y(_051_));
XNOR_g XNOR_g_130_(.A(key[2]), .B(inputs[2]), .Y(_052_));
XNOR_g XNOR_g_132_(.A(key[6]), .B(inputs[6]), .Y(_054_));
XNOR_g XNOR_g_133_(.A(key[4]), .B(inputs[4]), .Y(_055_));
XNOR_g XNOR_g_138_(.A(_059_), .B(s1.c.c[0]), .Y(out[1]));
AND_g AND_g_075_(.A(_002_), .B(_001_), .Y(_003_));
AND_g AND_g_078_(.A(_005_), .B(_004_), .Y(_006_));
AND_g AND_g_079_(.A(_006_), .B(_003_), .Y(_007_));
AND_g AND_g_082_(.A(_009_), .B(_008_), .Y(_010_));
AND_g AND_g_084_(.A(_000_), .B(inputs[0]), .Y(_012_));
AND_g AND_g_085_(.A(_012_), .B(_011_), .Y(_013_));
AND_g AND_g_089_(.A(_016_), .B(_015_), .Y(_017_));
AND_g AND_g_092_(.A(_019_), .B(_018_), .Y(_020_));
AND_g AND_g_093_(.A(_020_), .B(_017_), .Y(_021_));
AND_g AND_g_094_(.A(_021_), .B(_014_), .Y(_022_));
AND_g AND_g_097_(.A(inputs[4]), .B(inputs[0]), .Y(_024_));
AND_g AND_g_117_(.A(_038_), .B(_037_), .Y(_039_));
AND_g AND_g_120_(.A(_041_), .B(_040_), .Y(_042_));
AND_g AND_g_121_(.A(_042_), .B(_039_), .Y(_043_));
AND_g AND_g_124_(.A(_045_), .B(_044_), .Y(_046_));
AND_g AND_g_126_(.A(_036_), .B(inputs[0]), .Y(_048_));
AND_g AND_g_127_(.A(_048_), .B(_047_), .Y(_049_));
AND_g AND_g_131_(.A(_052_), .B(_051_), .Y(_053_));
AND_g AND_g_134_(.A(_055_), .B(_054_), .Y(_056_));
AND_g AND_g_135_(.A(_056_), .B(_053_), .Y(_057_));
AND_g AND_g_136_(.A(_057_), .B(_050_), .Y(_058_));
AND_g AND_g_139_(.A(inputs[4]), .B(inputs[0]), .Y(_060_));
NOR_g NOR_g_080_(.A(inputs[6]), .B(inputs[5]), .Y(_008_));
NOR_g NOR_g_081_(.A(inputs[7]), .B(inputs[4]), .Y(_009_));
NOR_g NOR_g_083_(.A(inputs[2]), .B(inputs[1]), .Y(_011_));
NOR_g NOR_g_122_(.A(inputs[6]), .B(inputs[5]), .Y(_044_));
NOR_g NOR_g_123_(.A(inputs[7]), .B(inputs[4]), .Y(_045_));
NOR_g NOR_g_125_(.A(inputs[2]), .B(inputs[1]), .Y(_047_));
NAND_g NAND_g_086_(.A(_013_), .B(_010_), .Y(_014_));
NAND_g NAND_g_095_(.A(_022_), .B(_007_), .Y(_023_));
NAND_g NAND_g_098_(.A(inputs[5]), .B(inputs[1]), .Y(_025_));
NAND_g NAND_g_100_(.A(_026_), .B(_024_), .Y(_027_));
NAND_g NAND_g_102_(.A(_027_), .B(_025_), .Y(_028_));
NAND_g NAND_g_103_(.A(inputs[6]), .B(inputs[2]), .Y(_029_));
NAND_g NAND_g_105_(.A(_030_), .B(_028_), .Y(_031_));
NAND_g NAND_g_107_(.A(_031_), .B(_029_), .Y(_032_));
NAND_g NAND_g_108_(.A(inputs[7]), .B(inputs[3]), .Y(_033_));
NAND_g NAND_g_110_(.A(_034_), .B(_032_), .Y(_035_));
NAND_g NAND_g_113_(.A(_035_), .B(_033_), .Y(s.c.c[4]));
NAND_g NAND_g_128_(.A(_049_), .B(_046_), .Y(_050_));
NAND_g NAND_g_137_(.A(_058_), .B(_043_), .Y(_059_));
NAND_g NAND_g_140_(.A(inputs[5]), .B(inputs[1]), .Y(_061_));
NAND_g NAND_g_142_(.A(_062_), .B(_060_), .Y(_063_));
NAND_g NAND_g_144_(.A(_063_), .B(_061_), .Y(_064_));
NAND_g NAND_g_145_(.A(inputs[6]), .B(inputs[2]), .Y(_065_));
NAND_g NAND_g_147_(.A(_066_), .B(_064_), .Y(_067_));
NAND_g NAND_g_149_(.A(_067_), .B(_065_), .Y(_068_));
NAND_g NAND_g_150_(.A(inputs[7]), .B(inputs[3]), .Y(_069_));
NAND_g NAND_g_152_(.A(_070_), .B(_068_), .Y(_071_));
NAND_g NAND_g_155_(.A(_071_), .B(_069_), .Y(s1.c.c[4]));
XOR_g XOR_g_099_(.A(inputs[5]), .B(inputs[1]), .Y(_026_));
XOR_g XOR_g_101_(.A(_026_), .B(_024_), .Y(s.c.c[1]));
XOR_g XOR_g_104_(.A(inputs[6]), .B(inputs[2]), .Y(_030_));
XOR_g XOR_g_106_(.A(_030_), .B(_028_), .Y(s.c.c[2]));
XOR_g XOR_g_109_(.A(inputs[7]), .B(inputs[3]), .Y(_034_));
XOR_g XOR_g_111_(.A(_034_), .B(_032_), .Y(s.c.c[3]));
XOR_g XOR_g_112_(.A(inputs[4]), .B(inputs[0]), .Y(s.c.c[0]));
XOR_g XOR_g_141_(.A(inputs[5]), .B(inputs[1]), .Y(_062_));
XOR_g XOR_g_143_(.A(_062_), .B(_060_), .Y(s1.c.c[1]));
XOR_g XOR_g_146_(.A(inputs[6]), .B(inputs[2]), .Y(_066_));
XOR_g XOR_g_148_(.A(_066_), .B(_064_), .Y(s1.c.c[2]));
XOR_g XOR_g_151_(.A(inputs[7]), .B(inputs[3]), .Y(_070_));
XOR_g XOR_g_153_(.A(_070_), .B(_068_), .Y(s1.c.c[3]));
XOR_g XOR_g_154_(.A(inputs[4]), .B(inputs[0]), .Y(s1.c.c[0]));
endmodule





module orgcir(inputs, key, out);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
input [7:0] inputs;
wire [7:0] inputs;
input [7:0] key;
wire [7:0] key;
output [1:0] out;
wire [1:0] out;
wire [4:0] s.c.c;
wire [4:0] s1.c.c;
NOT_g _072_ ( .A(inputs[3]), .Y(_000_) );
XNOR_g _073_ ( .A(inputs[0]), .B(key[0]), .Y(_001_) );
XNOR_g _074_ ( .A(inputs[7]), .B(key[7]), .Y(_002_) );
AND_g _075_ ( .A(_001_), .B(_002_), .Y(_003_) );
XNOR_g _076_ ( .A(inputs[1]), .B(key[1]), .Y(_004_) );
XNOR_g _077_ ( .A(inputs[3]), .B(key[3]), .Y(_005_) );
AND_g _078_ ( .A(_004_), .B(_005_), .Y(_006_) );
AND_g _079_ ( .A(_003_), .B(_006_), .Y(_007_) );
NOR_g _080_ ( .A(inputs[5]), .B(inputs[6]), .Y(_008_) );
NOR_g _081_ ( .A(inputs[4]), .B(inputs[7]), .Y(_009_) );
AND_g _082_ ( .A(_008_), .B(_009_), .Y(_010_) );
NOR_g _083_ ( .A(inputs[1]), .B(inputs[2]), .Y(_011_) );
AND_g _084_ ( .A(inputs[0]), .B(_000_), .Y(_012_) );
AND_g _085_ ( .A(_011_), .B(_012_), .Y(_013_) );
NAND_g _086_ ( .A(_010_), .B(_013_), .Y(_014_) );
XNOR_g _087_ ( .A(inputs[5]), .B(key[5]), .Y(_015_) );
XNOR_g _088_ ( .A(inputs[2]), .B(key[2]), .Y(_016_) );
AND_g _089_ ( .A(_015_), .B(_016_), .Y(_017_) );
XNOR_g _090_ ( .A(inputs[6]), .B(key[6]), .Y(_018_) );
XNOR_g _091_ ( .A(inputs[4]), .B(key[4]), .Y(_019_) );
AND_g _092_ ( .A(_018_), .B(_019_), .Y(_020_) );
AND_g _093_ ( .A(_017_), .B(_020_), .Y(_021_) );
AND_g _094_ ( .A(_014_), .B(_021_), .Y(_022_) );
NAND_g _095_ ( .A(_007_), .B(_022_), .Y(_023_) );
XNOR_g _096_ ( .A(s.c.c[0]), .B(_023_), .Y(out[0]) );
AND_g _097_ ( .A(inputs[0]), .B(inputs[4]), .Y(_024_) );
NAND_g _098_ ( .A(inputs[1]), .B(inputs[5]), .Y(_025_) );
XOR_g _099_ ( .A(inputs[1]), .B(inputs[5]), .Y(_026_) );
NAND_g _100_ ( .A(_024_), .B(_026_), .Y(_027_) );
XOR_g _101_ ( .A(_024_), .B(_026_), .Y(s.c.c[1]) );
NAND_g _102_ ( .A(_025_), .B(_027_), .Y(_028_) );
NAND_g _103_ ( .A(inputs[2]), .B(inputs[6]), .Y(_029_) );
XOR_g _104_ ( .A(inputs[2]), .B(inputs[6]), .Y(_030_) );
NAND_g _105_ ( .A(_028_), .B(_030_), .Y(_031_) );
XOR_g _106_ ( .A(_028_), .B(_030_), .Y(s.c.c[2]) );
NAND_g _107_ ( .A(_029_), .B(_031_), .Y(_032_) );
NAND_g _108_ ( .A(inputs[3]), .B(inputs[7]), .Y(_033_) );
XOR_g _109_ ( .A(inputs[3]), .B(inputs[7]), .Y(_034_) );
NAND_g _110_ ( .A(_032_), .B(_034_), .Y(_035_) );
XOR_g _111_ ( .A(_032_), .B(_034_), .Y(s.c.c[3]) );
XOR_g _112_ ( .A(inputs[0]), .B(inputs[4]), .Y(s.c.c[0]) );
NAND_g _113_ ( .A(_033_), .B(_035_), .Y(s.c.c[4]) );
NOT_g _114_ ( .A(inputs[3]), .Y(_036_) );
XNOR_g _115_ ( .A(inputs[0]), .B(key[0]), .Y(_037_) );
XNOR_g _116_ ( .A(inputs[7]), .B(key[7]), .Y(_038_) );
AND_g _117_ ( .A(_037_), .B(_038_), .Y(_039_) );
XNOR_g _118_ ( .A(inputs[1]), .B(key[1]), .Y(_040_) );
XNOR_g _119_ ( .A(inputs[3]), .B(key[3]), .Y(_041_) );
AND_g _120_ ( .A(_040_), .B(_041_), .Y(_042_) );
AND_g _121_ ( .A(_039_), .B(_042_), .Y(_043_) );
NOR_g _122_ ( .A(inputs[5]), .B(inputs[6]), .Y(_044_) );
NOR_g _123_ ( .A(inputs[4]), .B(inputs[7]), .Y(_045_) );
AND_g _124_ ( .A(_044_), .B(_045_), .Y(_046_) );
NOR_g _125_ ( .A(inputs[1]), .B(inputs[2]), .Y(_047_) );
AND_g _126_ ( .A(inputs[0]), .B(_036_), .Y(_048_) );
AND_g _127_ ( .A(_047_), .B(_048_), .Y(_049_) );
NAND_g _128_ ( .A(_046_), .B(_049_), .Y(_050_) );
XNOR_g _129_ ( .A(inputs[5]), .B(key[5]), .Y(_051_) );
XNOR_g _130_ ( .A(inputs[2]), .B(key[2]), .Y(_052_) );
AND_g _131_ ( .A(_051_), .B(_052_), .Y(_053_) );
XNOR_g _132_ ( .A(inputs[6]), .B(key[6]), .Y(_054_) );
XNOR_g _133_ ( .A(inputs[4]), .B(key[4]), .Y(_055_) );
AND_g _134_ ( .A(_054_), .B(_055_), .Y(_056_) );
AND_g _135_ ( .A(_053_), .B(_056_), .Y(_057_) );
AND_g _136_ ( .A(_050_), .B(_057_), .Y(_058_) );
NAND_g _137_ ( .A(_043_), .B(_058_), .Y(_059_) );
XNOR_g _138_ ( .A(s1.c.c[0]), .B(_059_), .Y(out[1]) );
AND_g _139_ ( .A(inputs[0]), .B(inputs[4]), .Y(_060_) );
NAND_g _140_ ( .A(inputs[1]), .B(inputs[5]), .Y(_061_) );
XOR_g _141_ ( .A(inputs[1]), .B(inputs[5]), .Y(_062_) );
NAND_g _142_ ( .A(_060_), .B(_062_), .Y(_063_) );
XOR_g _143_ ( .A(_060_), .B(_062_), .Y(s1.c.c[1]) );
NAND_g _144_ ( .A(_061_), .B(_063_), .Y(_064_) );
NAND_g _145_ ( .A(inputs[2]), .B(inputs[6]), .Y(_065_) );
XOR_g _146_ ( .A(inputs[2]), .B(inputs[6]), .Y(_066_) );
NAND_g _147_ ( .A(_064_), .B(_066_), .Y(_067_) );
XOR_g _148_ ( .A(_064_), .B(_066_), .Y(s1.c.c[2]) );
NAND_g _149_ ( .A(_065_), .B(_067_), .Y(_068_) );
NAND_g _150_ ( .A(inputs[3]), .B(inputs[7]), .Y(_069_) );
XOR_g _151_ ( .A(inputs[3]), .B(inputs[7]), .Y(_070_) );
NAND_g _152_ ( .A(_068_), .B(_070_), .Y(_071_) );
XOR_g _153_ ( .A(_068_), .B(_070_), .Y(s1.c.c[3]) );
XOR_g _154_ ( .A(inputs[0]), .B(inputs[4]), .Y(s1.c.c[0]) );
NAND_g _155_ ( .A(_069_), .B(_071_), .Y(s1.c.c[4]) );
endmodule
module BUF_g(A, Y);
input A;
output Y;
assign Y=A;
endmodule

 
module NOT_g(A, Y);
input A;
output Y;
assign Y=~A;
endmodule

module AND_g(A, B, Y);
input A, B;
output Y;
assign Y=(A & B);
endmodule

module OR_g(A, B, Y);
input A, B;
output Y;
assign Y= (A | B);
endmodule

module NAND_g(A, B, Y);
input A, B;
output Y;
assign Y= ~(A & B);

endmodule

module NOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A | B);
endmodule


module XOR_g(A, B, Y);
input A, B;
output Y;
assign Y = (A ^ B);
endmodule

module XNOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A ^ B);
endmodule

module DFFcell(C, D, Q);
input C, D;
output reg Q;
always @(posedge C)
	Q <= D;
endmodule


module DFFRcell(C, D, Q, R);
input C, D, R;
output reg Q;
always @(posedge C, negedge R)
	if (!R)
		Q <= 1'b0;
	else
		Q <= D;
endmodule
