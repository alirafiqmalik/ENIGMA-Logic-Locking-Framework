module top(inputs,key,lockingkeyinput,Q,Z);
input [7:0] inputs;
input [7:0] key;
input [255:0] lockingkeyinput;
wire [1:0] out_enc, out_org;
orgcir org(.inputs(inputs),.key(key),.out(out_org));
enccir enc(.inputs(inputs),.key(key),.lockingkeyinput(lockingkeyinput),.out(out_enc));
output Z;
output [1:0]Q;
assign Q[0]=out_enc[0]==out_org[0];
assign Q[1]=out_enc[1]==out_org[1];
assign Z= Q[0]&Q[1];
endmodule



module enccir(inputs,key,lockingkeyinput,out);
input [7:0] inputs;
input [7:0] key;
input [255:0] lockingkeyinput;
output [1:0] out;
wire _058_;
wire [4:0] s1cc;
wire _040_;
wire _002_;
wire _010_;
wire _052_;
wire _003_;
wire _060_;
wire _053_;
wire _042_;
wire _046_;
wire _056_;
wire _034_;
wire _032_;
wire _022_;
wire _024_;
wire _065_;
wire _012_;
wire _069_;
wire _015_;
wire _029_;
wire _039_;
wire _036_;
wire _066_;
wire _007_;
wire _008_;
wire _017_;
wire _070_;
wire _011_;
wire _064_;
wire _051_;
wire _021_;
wire _030_;
wire _059_;
wire _025_;
wire _001_;
wire [4:0] scc;
wire _067_;
wire _057_;
wire _019_;
wire _049_;
wire _054_;
wire _005_;
wire _023_;
wire _006_;
wire _037_;
wire _045_;
wire _068_;
wire _004_;
wire _055_;
wire _018_;
wire _043_;
wire _062_;
wire _044_;
wire _027_;
wire _038_;
wire _009_;
wire _000_;
wire _047_;
wire _061_;
wire _071_;
wire _031_;
wire _014_;
wire _013_;
wire _048_;
wire _026_;
wire _050_;
wire _016_;
wire _063_;
wire _035_;
wire _041_;
wire _028_;
wire _033_;
wire _020_;
wire keywire74;
wire keywire75;
wire keywire76;
wire keywire77;
wire keywire78;
wire keywire79;
wire keywire80;
wire keywire81;
wire keywire82;
wire keywire83;
wire keywire84;
wire keywire85;
wire keywire86;
wire keywire87;
wire keywire88;
wire keywire89;
wire keywire90;
wire keywire91;
wire keywire92;
wire keywire93;
wire keywire94;
wire keywire95;
wire keywire96;
wire keywire97;
wire keywire98;
wire keywire99;
wire keywire100;
wire keywire101;
wire keywire102;
wire keywire103;
wire keywire104;
wire keywire105;
wire keywire106;
wire keywire107;
wire keywire108;
wire keywire109;
wire keywire110;
wire keywire111;
wire keywire112;
wire keywire113;
wire keywire114;
wire keywire115;
wire keywire116;
wire keywire117;
wire keywire118;
wire keywire119;
wire keywire120;
wire keywire121;
wire keywire122;
wire keywire123;
wire keywire124;
wire keywire125;
wire keywire126;
wire keywire127;
wire keywire128;
wire keywire129;
wire keywire130;
wire keywire131;
wire keywire132;
wire keywire133;
wire keywire134;
wire keywire135;
wire keywire136;
wire keywire137;
wire keywire138;
wire keywire139;
wire keywire140;
wire keywire141;
wire keywire142;
wire keywire143;
wire keywire144;
wire keywire145;
wire keywire146;
wire keywire147;
wire keywire148;
wire keywire149;
wire keywire150;
wire keywire151;
wire keywire152;
wire keywire153;
wire keywire154;
wire keywire155;
wire keywire156;
wire keywire157;
wire keywire158;
wire keywire159;
wire keywire160;
wire keywire161;
wire keywire162;
wire keywire163;
wire keywire164;
wire keywire165;
wire keywire166;
wire keywire167;
wire keywire168;
wire keywire169;
wire keywire170;
wire keywire171;
wire keywire172;
wire keywire173;
wire keywire174;
wire keywire175;
wire keywire176;
wire keywire177;
wire keywire178;
wire keywire179;
wire keywire180;
wire keywire181;
wire keywire182;
wire keywire183;
wire keywire184;
wire keywire185;
wire keywire186;
wire keywire187;
wire keywire188;
wire keywire189;
wire keywire190;
wire keywire191;
wire keywire192;
wire keywire193;
wire keywire194;
wire keywire195;
wire keywire196;
wire keywire197;
wire keywire198;
wire keywire199;
wire keywire200;
wire keywire201;
wire keywire202;
wire keywire203;
wire keywire204;
wire keywire205;
wire keywire206;
wire keywire207;
wire keywire208;
wire keywire209;
wire keywire210;
wire keywire211;
wire keywire212;
wire keywire213;
wire keywire214;
wire keywire215;
wire keywire216;
wire keywire217;
wire keywire218;
wire keywire219;
wire keywire220;
wire keywire221;
wire keywire222;
wire keywire223;
wire keywire224;
wire keywire225;
wire keywire226;
wire keywire227;
wire keywire228;
wire keywire229;
wire keywire230;
wire keywire231;
wire keywire232;
wire keywire233;
wire keywire234;
wire keywire235;
wire keywire236;
wire keywire237;
wire keywire238;
wire keywire239;
wire keywire240;
wire keywire241;
wire keywire242;
wire keywire243;
wire keywire244;
wire keywire245;
wire keywire246;
wire keywire247;
wire keywire248;
wire keywire249;
wire keywire250;
wire keywire251;
wire keywire252;
wire keywire253;
wire keywire254;
wire keywire255;
wire keywire256;
wire keywire257;
wire keywire258;
wire keywire259;
wire keywire260;
wire keywire261;
wire keywire262;
wire keywire263;
wire keywire264;
wire keywire265;
wire keywire266;
wire keywire267;
wire keywire268;
wire keywire269;
wire keywire270;
wire keywire271;
wire keywire272;
wire keywire273;
wire keywire274;
wire keywire275;
wire keywire276;
wire keywire277;
wire keywire278;
wire keywire279;
wire keywire280;
wire keywire281;
wire keywire282;
wire keywire283;
wire keywire284;
wire keywire285;
wire keywire286;
wire keywire287;
wire keywire288;
wire keywire289;
wire keywire290;
wire keywire291;
wire keywire292;
wire keywire293;
wire keywire294;
wire keywire295;
wire keywire296;
wire keywire297;
wire keywire298;
wire keywire299;
wire keywire300;
wire keywire301;
wire keywire302;
wire keywire303;
wire keywire304;
wire keywire305;
wire keywire306;
wire keywire307;
wire keywire308;
wire keywire309;
wire keywire310;
wire keywire311;
wire keywire312;
wire keywire313;
wire keywire314;
wire keywire315;
wire keywire316;
wire keywire317;
wire keywire318;
wire keywire319;
wire keywire320;
wire keywire321;
wire keywire322;
wire keywire323;
wire keywire324;
wire keywire325;
wire keywire326;
wire keywire327;
wire keywire328;
wire keywire329;
NOT_g NOT_g_072_(.A(inputs[3]), .Y(keywire237));
NOT_g NOT_g_114_(.A(inputs[3]), .Y(keywire297));
XNOR_g XNOR_g_073_(.A(key[0]), .B(inputs[0]), .Y(keywire321));
XNOR_g XNOR_g_074_(.A(key[7]), .B(inputs[7]), .Y(keywire320));
XNOR_g XNOR_g_076_(.A(key[1]), .B(inputs[1]), .Y(keywire319));
XNOR_g XNOR_g_077_(.A(key[3]), .B(inputs[3]), .Y(keywire318));
XNOR_g XNOR_g_087_(.A(key[5]), .B(inputs[5]), .Y(keywire249));
XNOR_g XNOR_g_088_(.A(key[2]), .B(inputs[2]), .Y(keywire231));
XNOR_g XNOR_g_090_(.A(key[6]), .B(inputs[6]), .Y(keywire253));
XNOR_g XNOR_g_091_(.A(key[4]), .B(inputs[4]), .Y(keywire245));
XNOR_g XNOR_g_096_(.A(_023_), .B(scc[0]), .Y(keywire295));
XNOR_g XNOR_g_115_(.A(key[0]), .B(inputs[0]), .Y(keywire329));
XNOR_g XNOR_g_116_(.A(key[7]), .B(inputs[7]), .Y(keywire328));
XNOR_g XNOR_g_118_(.A(key[1]), .B(inputs[1]), .Y(keywire327));
XNOR_g XNOR_g_119_(.A(key[3]), .B(inputs[3]), .Y(keywire326));
XNOR_g XNOR_g_129_(.A(key[5]), .B(inputs[5]), .Y(keywire250));
XNOR_g XNOR_g_130_(.A(key[2]), .B(inputs[2]), .Y(keywire232));
XNOR_g XNOR_g_132_(.A(key[6]), .B(inputs[6]), .Y(keywire254));
XNOR_g XNOR_g_133_(.A(key[4]), .B(inputs[4]), .Y(keywire246));
XNOR_g XNOR_g_138_(.A(_059_), .B(s1cc[0]), .Y(keywire296));
XNOR_g keygate_XNOR_0(.A(keywire74), .B(lockingkeyinput[0]), .Y(_049_));
XNOR_g keygate_XNOR_3(.A(keywire77), .B(lockingkeyinput[3]), .Y(_059_));
XNOR_g keygate_XNOR_4(.A(keywire78), .B(lockingkeyinput[4]), .Y(out[1]));
XNOR_g keygate_XNOR_5(.A(keywire79), .B(lockingkeyinput[5]), .Y(_001_));
XNOR_g keygate_XNOR_7(.A(keywire81), .B(lockingkeyinput[7]), .Y(_012_));
XNOR_g keygate_XNOR_8(.A(keywire82), .B(lockingkeyinput[8]), .Y(_024_));
XNOR_g keygate_XNOR_9(.A(keywire83), .B(lockingkeyinput[9]), .Y(_048_));
XNOR_g keygate_XNOR_11(.A(keywire85), .B(lockingkeyinput[11]), .Y(scc[0]));
XNOR_g keygate_XNOR_14(.A(keywire88), .B(lockingkeyinput[14]), .Y(_040_));
XNOR_g keygate_XNOR_15(.A(keywire89), .B(lockingkeyinput[15]), .Y(_011_));
XNOR_g keygate_XNOR_17(.A(keywire91), .B(lockingkeyinput[17]), .Y(_025_));
XNOR_g keygate_XNOR_19(.A(keywire93), .B(lockingkeyinput[19]), .Y(_026_));
XNOR_g keygate_XNOR_21(.A(keywire95), .B(lockingkeyinput[21]), .Y(_016_));
XNOR_g keygate_XNOR_22(.A(keywire96), .B(lockingkeyinput[22]), .Y(_052_));
XNOR_g keygate_XNOR_26(.A(keywire100), .B(lockingkeyinput[26]), .Y(_066_));
XNOR_g keygate_XNOR_27(.A(keywire101), .B(lockingkeyinput[27]), .Y(_000_));
XNOR_g keygate_XNOR_28(.A(keywire102), .B(lockingkeyinput[28]), .Y(_036_));
XNOR_g keygate_XNOR_29(.A(keywire103), .B(lockingkeyinput[29]), .Y(_005_));
XNOR_g keygate_XNOR_31(.A(keywire105), .B(lockingkeyinput[31]), .Y(_033_));
XNOR_g keygate_XNOR_34(.A(keywire108), .B(lockingkeyinput[34]), .Y(_070_));
XNOR_g keygate_XNOR_38(.A(keywire112), .B(lockingkeyinput[38]), .Y(_045_));
XNOR_g keygate_XNOR_39(.A(keywire113), .B(lockingkeyinput[39]), .Y(_015_));
XNOR_g keygate_XNOR_42(.A(keywire116), .B(lockingkeyinput[42]), .Y(_044_));
XNOR_g keygate_XNOR_43(.A(keywire117), .B(lockingkeyinput[43]), .Y(_018_));
XNOR_g keygate_XNOR_45(.A(keywire119), .B(lockingkeyinput[45]), .Y(_002_));
XNOR_g keygate_XNOR_50(.A(keywire124), .B(lockingkeyinput[50]), .Y(_027_));
XNOR_g keygate_XNOR_52(.A(keywire126), .B(lockingkeyinput[52]), .Y(_063_));
XNOR_g keygate_XNOR_57(.A(keywire131), .B(lockingkeyinput[57]), .Y(_028_));
XNOR_g keygate_XNOR_58(.A(keywire132), .B(lockingkeyinput[58]), .Y(_064_));
XNOR_g keygate_XNOR_59(.A(keywire133), .B(lockingkeyinput[59]), .Y(_017_));
XNOR_g keygate_XNOR_61(.A(keywire135), .B(lockingkeyinput[61]), .Y(_032_));
XNOR_g keygate_XNOR_62(.A(keywire136), .B(lockingkeyinput[62]), .Y(_068_));
XNOR_g keygate_XNOR_64(.A(keywire138), .B(lockingkeyinput[64]), .Y(scc[2]));
XNOR_g keygate_XNOR_65(.A(keywire139), .B(lockingkeyinput[65]), .Y(_067_));
XNOR_g keygate_XNOR_66(.A(keywire140), .B(lockingkeyinput[66]), .Y(s1cc[2]));
XNOR_g keygate_XNOR_67(.A(keywire141), .B(lockingkeyinput[67]), .Y(scc[4]));
XNOR_g keygate_XNOR_68(.A(keywire142), .B(lockingkeyinput[68]), .Y(s1cc[4]));
XNOR_g keygate_XNOR_72(.A(keywire146), .B(lockingkeyinput[72]), .Y(s1cc[3]));
XNOR_g keygate_XNOR_77(.A(keywire151), .B(lockingkeyinput[77]), .Y(_007_));
XNOR_g keygate_XNOR_81(.A(keywire155), .B(lockingkeyinput[81]), .Y(_057_));
XNOR_g keygate_XNOR_82(.A(keywire156), .B(lockingkeyinput[82]), .Y(_023_));
XNOR_g keygate_XNOR_83(.A(keywire157), .B(lockingkeyinput[83]), .Y(_022_));
XNOR_g keygate_XNOR_84(.A(keywire158), .B(lockingkeyinput[84]), .Y(keywire83));
XNOR_g keygate_XNOR_87(.A(keywire161), .B(lockingkeyinput[87]), .Y(keywire78));
XNOR_g keygate_XNOR_92(.A(keywire166), .B(lockingkeyinput[92]), .Y(keywire157));
XNOR_g keygate_XNOR_95(.A(keywire169), .B(lockingkeyinput[95]), .Y(keywire152));
XNOR_g keygate_XNOR_96(.A(keywire170), .B(lockingkeyinput[96]), .Y(keywire154));
XNOR_g keygate_XNOR_97(.A(keywire171), .B(lockingkeyinput[97]), .Y(keywire153));
XNOR_g keygate_XNOR_98(.A(keywire172), .B(lockingkeyinput[98]), .Y(keywire129));
XNOR_g keygate_XNOR_99(.A(keywire173), .B(lockingkeyinput[99]), .Y(keywire121));
XNOR_g keygate_XNOR_101(.A(keywire175), .B(lockingkeyinput[101]), .Y(keywire75));
XNOR_g keygate_XNOR_103(.A(keywire177), .B(lockingkeyinput[103]), .Y(keywire122));
XNOR_g keygate_XNOR_107(.A(keywire181), .B(lockingkeyinput[107]), .Y(keywire149));
XNOR_g keygate_XNOR_108(.A(keywire182), .B(lockingkeyinput[108]), .Y(keywire103));
XNOR_g keygate_XNOR_112(.A(keywire186), .B(lockingkeyinput[112]), .Y(keywire148));
XNOR_g keygate_XNOR_114(.A(keywire188), .B(lockingkeyinput[114]), .Y(keywire74));
XNOR_g keygate_XNOR_116(.A(keywire190), .B(lockingkeyinput[116]), .Y(keywire104));
XNOR_g keygate_XNOR_118(.A(keywire192), .B(lockingkeyinput[118]), .Y(keywire120));
XNOR_g keygate_XNOR_120(.A(keywire194), .B(lockingkeyinput[120]), .Y(keywire109));
XNOR_g keygate_XNOR_122(.A(keywire196), .B(lockingkeyinput[122]), .Y(keywire95));
XNOR_g keygate_XNOR_123(.A(keywire197), .B(lockingkeyinput[123]), .Y(keywire113));
XNOR_g keygate_XNOR_125(.A(keywire199), .B(lockingkeyinput[125]), .Y(keywire89));
XNOR_g keygate_XNOR_126(.A(keywire200), .B(lockingkeyinput[126]), .Y(keywire111));
XNOR_g keygate_XNOR_128(.A(keywire202), .B(lockingkeyinput[128]), .Y(keywire110));
XNOR_g keygate_XNOR_129(.A(keywire203), .B(lockingkeyinput[129]), .Y(keywire118));
XNOR_g keygate_XNOR_131(.A(keywire205), .B(lockingkeyinput[131]), .Y(keywire114));
XNOR_g keygate_XNOR_132(.A(keywire206), .B(lockingkeyinput[132]), .Y(keywire90));
XNOR_g keygate_XNOR_135(.A(keywire209), .B(lockingkeyinput[135]), .Y(keywire101));
XNOR_g keygate_XNOR_138(.A(keywire212), .B(lockingkeyinput[138]), .Y(keywire168));
XNOR_g keygate_XNOR_141(.A(keywire215), .B(lockingkeyinput[141]), .Y(keywire185));
XNOR_g keygate_XNOR_142(.A(keywire216), .B(lockingkeyinput[142]), .Y(keywire193));
XNOR_g keygate_XNOR_143(.A(keywire217), .B(lockingkeyinput[143]), .Y(keywire198));
XNOR_g keygate_XNOR_144(.A(keywire218), .B(lockingkeyinput[144]), .Y(keywire82));
XNOR_g keygate_XNOR_147(.A(keywire221), .B(lockingkeyinput[147]), .Y(keywire163));
XNOR_g keygate_XNOR_148(.A(keywire222), .B(lockingkeyinput[148]), .Y(keywire165));
XNOR_g keygate_XNOR_149(.A(keywire223), .B(lockingkeyinput[149]), .Y(keywire183));
XNOR_g keygate_XNOR_150(.A(keywire224), .B(lockingkeyinput[150]), .Y(keywire191));
XNOR_g keygate_XNOR_151(.A(keywire225), .B(lockingkeyinput[151]), .Y(keywire199));
XNOR_g keygate_XNOR_152(.A(keywire226), .B(lockingkeyinput[152]), .Y(keywire206));
XNOR_g keygate_XNOR_153(.A(keywire227), .B(lockingkeyinput[153]), .Y(keywire91));
XNOR_g keygate_XNOR_154(.A(keywire228), .B(lockingkeyinput[154]), .Y(keywire92));
XNOR_g keygate_XNOR_155(.A(keywire229), .B(lockingkeyinput[155]), .Y(keywire93));
XNOR_g keygate_XNOR_156(.A(keywire230), .B(lockingkeyinput[156]), .Y(keywire94));
XNOR_g keygate_XNOR_157(.A(keywire231), .B(lockingkeyinput[157]), .Y(keywire196));
XNOR_g keygate_XNOR_159(.A(keywire233), .B(lockingkeyinput[159]), .Y(keywire97));
XNOR_g keygate_XNOR_160(.A(keywire234), .B(lockingkeyinput[160]), .Y(keywire98));
XNOR_g keygate_XNOR_162(.A(keywire236), .B(lockingkeyinput[162]), .Y(keywire100));
XNOR_g keygate_XNOR_163(.A(keywire237), .B(lockingkeyinput[163]), .Y(keywire209));
XNOR_g keygate_XNOR_164(.A(keywire238), .B(lockingkeyinput[164]), .Y(keywire159));
XNOR_g keygate_XNOR_165(.A(keywire239), .B(lockingkeyinput[165]), .Y(keywire182));
XNOR_g keygate_XNOR_168(.A(keywire242), .B(lockingkeyinput[168]), .Y(keywire106));
XNOR_g keygate_XNOR_169(.A(keywire243), .B(lockingkeyinput[169]), .Y(keywire107));
XNOR_g keygate_XNOR_170(.A(keywire244), .B(lockingkeyinput[170]), .Y(keywire108));
XNOR_g keygate_XNOR_172(.A(keywire246), .B(lockingkeyinput[172]), .Y(keywire202));
XNOR_g keygate_XNOR_173(.A(keywire247), .B(lockingkeyinput[173]), .Y(keywire200));
XNOR_g keygate_XNOR_174(.A(keywire248), .B(lockingkeyinput[174]), .Y(keywire207));
XNOR_g keygate_XNOR_179(.A(keywire253), .B(lockingkeyinput[179]), .Y(keywire195));
XNOR_g keygate_XNOR_180(.A(keywire254), .B(lockingkeyinput[180]), .Y(keywire203));
XNOR_g keygate_XNOR_181(.A(keywire255), .B(lockingkeyinput[181]), .Y(keywire184));
XNOR_g keygate_XNOR_182(.A(keywire256), .B(lockingkeyinput[182]), .Y(keywire192));
XNOR_g keygate_XNOR_189(.A(keywire263), .B(lockingkeyinput[189]), .Y(keywire127));
XNOR_g keygate_XNOR_195(.A(keywire269), .B(lockingkeyinput[195]), .Y(keywire179));
XNOR_g keygate_XNOR_196(.A(keywire270), .B(lockingkeyinput[196]), .Y(keywire187));
XNOR_g keygate_XNOR_197(.A(keywire271), .B(lockingkeyinput[197]), .Y(keywire135));
XNOR_g keygate_XNOR_198(.A(keywire272), .B(lockingkeyinput[198]), .Y(keywire136));
XNOR_g keygate_XNOR_200(.A(keywire274), .B(lockingkeyinput[200]), .Y(keywire138));
XNOR_g keygate_XNOR_201(.A(keywire275), .B(lockingkeyinput[201]), .Y(keywire139));
XNOR_g keygate_XNOR_202(.A(keywire276), .B(lockingkeyinput[202]), .Y(keywire140));
XNOR_g keygate_XNOR_203(.A(keywire277), .B(lockingkeyinput[203]), .Y(keywire141));
XNOR_g keygate_XNOR_206(.A(keywire280), .B(lockingkeyinput[206]), .Y(keywire144));
XNOR_g keygate_XNOR_209(.A(keywire283), .B(lockingkeyinput[209]), .Y(keywire178));
XNOR_g keygate_XNOR_211(.A(keywire285), .B(lockingkeyinput[211]), .Y(keywire181));
XNOR_g keygate_XNOR_212(.A(keywire286), .B(lockingkeyinput[212]), .Y(keywire189));
XNOR_g keygate_XNOR_215(.A(keywire289), .B(lockingkeyinput[215]), .Y(keywire171));
XNOR_g keygate_XNOR_217(.A(keywire291), .B(lockingkeyinput[217]), .Y(keywire174));
XNOR_g keygate_XNOR_218(.A(keywire292), .B(lockingkeyinput[218]), .Y(keywire162));
XNOR_g keygate_XNOR_219(.A(keywire293), .B(lockingkeyinput[219]), .Y(keywire166));
XNOR_g keygate_XNOR_225(.A(keywire299), .B(lockingkeyinput[225]), .Y(keywire221));
XNOR_g keygate_XNOR_228(.A(keywire302), .B(lockingkeyinput[228]), .Y(keywire293));
XNOR_g keygate_XNOR_233(.A(keywire307), .B(lockingkeyinput[233]), .Y(keywire289));
XNOR_g keygate_XNOR_236(.A(keywire310), .B(lockingkeyinput[236]), .Y(keywire291));
XNOR_g keygate_XNOR_238(.A(keywire312), .B(lockingkeyinput[238]), .Y(keywire266));
XNOR_g keygate_XNOR_242(.A(keywire316), .B(lockingkeyinput[242]), .Y(keywire259));
XNOR_g keygate_XNOR_243(.A(keywire317), .B(lockingkeyinput[243]), .Y(keywire285));
XNOR_g keygate_XNOR_248(.A(keywire322), .B(lockingkeyinput[248]), .Y(keywire284));
XNOR_g keygate_XNOR_254(.A(keywire328), .B(lockingkeyinput[254]), .Y(keywire256));
XNOR_g keygate_XNOR_255(.A(keywire329), .B(lockingkeyinput[255]), .Y(keywire216));
AND_g AND_g_075_(.A(_002_), .B(_001_), .Y(keywire309));
AND_g AND_g_078_(.A(_005_), .B(_004_), .Y(keywire308));
AND_g AND_g_079_(.A(_006_), .B(_003_), .Y(keywire303));
AND_g AND_g_082_(.A(_009_), .B(_008_), .Y(keywire317));
AND_g AND_g_084_(.A(_000_), .B(inputs[0]), .Y(keywire217));
AND_g AND_g_085_(.A(_012_), .B(_011_), .Y(keywire316));
AND_g AND_g_089_(.A(_016_), .B(_015_), .Y(keywire315));
AND_g AND_g_092_(.A(_019_), .B(_018_), .Y(keywire314));
AND_g AND_g_093_(.A(_020_), .B(_017_), .Y(keywire306));
AND_g AND_g_094_(.A(_021_), .B(_014_), .Y(keywire302));
AND_g AND_g_097_(.A(inputs[4]), .B(inputs[0]), .Y(keywire218));
AND_g AND_g_117_(.A(_038_), .B(_037_), .Y(keywire313));
AND_g AND_g_120_(.A(_041_), .B(_040_), .Y(keywire312));
AND_g AND_g_121_(.A(_042_), .B(_039_), .Y(keywire305));
AND_g AND_g_124_(.A(_045_), .B(_044_), .Y(keywire325));
AND_g AND_g_126_(.A(_036_), .B(inputs[0]), .Y(keywire294));
AND_g AND_g_127_(.A(_048_), .B(_047_), .Y(keywire324));
AND_g AND_g_131_(.A(_052_), .B(_051_), .Y(keywire323));
AND_g AND_g_134_(.A(_055_), .B(_054_), .Y(keywire322));
AND_g AND_g_135_(.A(_056_), .B(_053_), .Y(keywire310));
AND_g AND_g_136_(.A(_057_), .B(_050_), .Y(keywire304));
AND_g AND_g_139_(.A(inputs[4]), .B(inputs[0]), .Y(keywire220));
NOR_g NOR_g_080_(.A(inputs[6]), .B(inputs[5]), .Y(keywire251));
NOR_g NOR_g_081_(.A(inputs[7]), .B(inputs[4]), .Y(keywire247));
NOR_g NOR_g_083_(.A(inputs[2]), .B(inputs[1]), .Y(keywire225));
NOR_g NOR_g_122_(.A(inputs[6]), .B(inputs[5]), .Y(keywire252));
NOR_g NOR_g_123_(.A(inputs[7]), .B(inputs[4]), .Y(keywire248));
NOR_g NOR_g_125_(.A(inputs[2]), .B(inputs[1]), .Y(keywire226));
NAND_g NAND_g_086_(.A(_013_), .B(_010_), .Y(keywire307));
NAND_g NAND_g_095_(.A(_022_), .B(_007_), .Y(keywire298));
NAND_g NAND_g_098_(.A(inputs[5]), .B(inputs[1]), .Y(keywire227));
NAND_g NAND_g_100_(.A(_026_), .B(_024_), .Y(keywire260));
NAND_g NAND_g_102_(.A(_027_), .B(_025_), .Y(keywire267));
NAND_g NAND_g_103_(.A(inputs[6]), .B(inputs[2]), .Y(keywire233));
NAND_g NAND_g_105_(.A(_030_), .B(_028_), .Y(keywire273));
NAND_g NAND_g_107_(.A(_031_), .B(_029_), .Y(keywire271));
NAND_g NAND_g_108_(.A(inputs[7]), .B(inputs[3]), .Y(keywire241));
NAND_g NAND_g_110_(.A(_034_), .B(_032_), .Y(keywire279));
NAND_g NAND_g_113_(.A(_035_), .B(_033_), .Y(keywire277));
NAND_g NAND_g_128_(.A(_049_), .B(_046_), .Y(keywire311));
NAND_g NAND_g_137_(.A(_058_), .B(_043_), .Y(keywire300));
NAND_g NAND_g_140_(.A(inputs[5]), .B(inputs[1]), .Y(keywire228));
NAND_g NAND_g_142_(.A(_062_), .B(_060_), .Y(keywire262));
NAND_g NAND_g_144_(.A(_063_), .B(_061_), .Y(keywire268));
NAND_g NAND_g_145_(.A(inputs[6]), .B(inputs[2]), .Y(keywire234));
NAND_g NAND_g_147_(.A(_066_), .B(_064_), .Y(keywire275));
NAND_g NAND_g_149_(.A(_067_), .B(_065_), .Y(keywire272));
NAND_g NAND_g_150_(.A(inputs[7]), .B(inputs[3]), .Y(keywire242));
NAND_g NAND_g_152_(.A(_070_), .B(_068_), .Y(keywire281));
NAND_g NAND_g_155_(.A(_071_), .B(_069_), .Y(keywire278));
XOR_g XOR_g_099_(.A(inputs[5]), .B(inputs[1]), .Y(keywire229));
XOR_g XOR_g_101_(.A(_026_), .B(_024_), .Y(keywire261));
XOR_g XOR_g_104_(.A(inputs[6]), .B(inputs[2]), .Y(keywire235));
XOR_g XOR_g_106_(.A(_030_), .B(_028_), .Y(keywire274));
XOR_g XOR_g_109_(.A(inputs[7]), .B(inputs[3]), .Y(keywire243));
XOR_g XOR_g_111_(.A(_034_), .B(_032_), .Y(keywire280));
XOR_g XOR_g_112_(.A(inputs[4]), .B(inputs[0]), .Y(keywire299));
XOR_g XOR_g_141_(.A(inputs[5]), .B(inputs[1]), .Y(keywire230));
XOR_g XOR_g_143_(.A(_062_), .B(_060_), .Y(keywire263));
XOR_g XOR_g_146_(.A(inputs[6]), .B(inputs[2]), .Y(keywire236));
XOR_g XOR_g_148_(.A(_066_), .B(_064_), .Y(keywire276));
XOR_g XOR_g_151_(.A(inputs[7]), .B(inputs[3]), .Y(keywire244));
XOR_g XOR_g_153_(.A(_070_), .B(_068_), .Y(keywire282));
XOR_g XOR_g_154_(.A(inputs[4]), .B(inputs[0]), .Y(keywire301));
XOR_g keygate_XOR_1(.A(keywire75), .B(lockingkeyinput[1]), .Y(_050_));
XOR_g keygate_XOR_2(.A(keywire76), .B(lockingkeyinput[2]), .Y(_058_));
XOR_g keygate_XOR_6(.A(keywire80), .B(lockingkeyinput[6]), .Y(_037_));
XOR_g keygate_XOR_10(.A(keywire84), .B(lockingkeyinput[10]), .Y(_060_));
XOR_g keygate_XOR_12(.A(keywire86), .B(lockingkeyinput[12]), .Y(s1cc[0]));
XOR_g keygate_XOR_13(.A(keywire87), .B(lockingkeyinput[13]), .Y(_004_));
XOR_g keygate_XOR_16(.A(keywire90), .B(lockingkeyinput[16]), .Y(_047_));
XOR_g keygate_XOR_18(.A(keywire92), .B(lockingkeyinput[18]), .Y(_061_));
XOR_g keygate_XOR_20(.A(keywire94), .B(lockingkeyinput[20]), .Y(_062_));
XOR_g keygate_XOR_23(.A(keywire97), .B(lockingkeyinput[23]), .Y(_029_));
XOR_g keygate_XOR_24(.A(keywire98), .B(lockingkeyinput[24]), .Y(_065_));
XOR_g keygate_XOR_25(.A(keywire99), .B(lockingkeyinput[25]), .Y(_030_));
XOR_g keygate_XOR_30(.A(keywire104), .B(lockingkeyinput[30]), .Y(_041_));
XOR_g keygate_XOR_32(.A(keywire106), .B(lockingkeyinput[32]), .Y(_069_));
XOR_g keygate_XOR_33(.A(keywire107), .B(lockingkeyinput[33]), .Y(_034_));
XOR_g keygate_XOR_35(.A(keywire109), .B(lockingkeyinput[35]), .Y(_019_));
XOR_g keygate_XOR_36(.A(keywire110), .B(lockingkeyinput[36]), .Y(_055_));
XOR_g keygate_XOR_37(.A(keywire111), .B(lockingkeyinput[37]), .Y(_009_));
XOR_g keygate_XOR_40(.A(keywire114), .B(lockingkeyinput[40]), .Y(_051_));
XOR_g keygate_XOR_41(.A(keywire115), .B(lockingkeyinput[41]), .Y(_008_));
XOR_g keygate_XOR_44(.A(keywire118), .B(lockingkeyinput[44]), .Y(_054_));
XOR_g keygate_XOR_46(.A(keywire120), .B(lockingkeyinput[46]), .Y(_038_));
XOR_g keygate_XOR_47(.A(keywire121), .B(lockingkeyinput[47]), .Y(_003_));
XOR_g keygate_XOR_48(.A(keywire122), .B(lockingkeyinput[48]), .Y(_039_));
XOR_g keygate_XOR_49(.A(keywire123), .B(lockingkeyinput[49]), .Y(_013_));
XOR_g keygate_XOR_51(.A(keywire125), .B(lockingkeyinput[51]), .Y(scc[1]));
XOR_g keygate_XOR_53(.A(keywire127), .B(lockingkeyinput[53]), .Y(s1cc[1]));
XOR_g keygate_XOR_54(.A(keywire128), .B(lockingkeyinput[54]), .Y(out[0]));
XOR_g keygate_XOR_55(.A(keywire129), .B(lockingkeyinput[55]), .Y(_006_));
XOR_g keygate_XOR_56(.A(keywire130), .B(lockingkeyinput[56]), .Y(_042_));
XOR_g keygate_XOR_60(.A(keywire134), .B(lockingkeyinput[60]), .Y(_053_));
XOR_g keygate_XOR_63(.A(keywire137), .B(lockingkeyinput[63]), .Y(_031_));
XOR_g keygate_XOR_69(.A(keywire143), .B(lockingkeyinput[69]), .Y(_035_));
XOR_g keygate_XOR_70(.A(keywire144), .B(lockingkeyinput[70]), .Y(scc[3]));
XOR_g keygate_XOR_71(.A(keywire145), .B(lockingkeyinput[71]), .Y(_071_));
XOR_g keygate_XOR_73(.A(keywire147), .B(lockingkeyinput[73]), .Y(_020_));
XOR_g keygate_XOR_74(.A(keywire148), .B(lockingkeyinput[74]), .Y(_056_));
XOR_g keygate_XOR_75(.A(keywire149), .B(lockingkeyinput[75]), .Y(_010_));
XOR_g keygate_XOR_76(.A(keywire150), .B(lockingkeyinput[76]), .Y(_046_));
XOR_g keygate_XOR_78(.A(keywire152), .B(lockingkeyinput[78]), .Y(_043_));
XOR_g keygate_XOR_79(.A(keywire153), .B(lockingkeyinput[79]), .Y(_014_));
XOR_g keygate_XOR_80(.A(keywire154), .B(lockingkeyinput[80]), .Y(_021_));
XOR_g keygate_XOR_85(.A(keywire159), .B(lockingkeyinput[85]), .Y(keywire102));
XOR_g keygate_XOR_86(.A(keywire160), .B(lockingkeyinput[86]), .Y(keywire128));
XOR_g keygate_XOR_88(.A(keywire162), .B(lockingkeyinput[88]), .Y(keywire156));
XOR_g keygate_XOR_89(.A(keywire163), .B(lockingkeyinput[89]), .Y(keywire85));
XOR_g keygate_XOR_90(.A(keywire164), .B(lockingkeyinput[90]), .Y(keywire77));
XOR_g keygate_XOR_91(.A(keywire165), .B(lockingkeyinput[91]), .Y(keywire86));
XOR_g keygate_XOR_93(.A(keywire167), .B(lockingkeyinput[93]), .Y(keywire151));
XOR_g keygate_XOR_94(.A(keywire168), .B(lockingkeyinput[94]), .Y(keywire76));
XOR_g keygate_XOR_100(.A(keywire174), .B(lockingkeyinput[100]), .Y(keywire155));
XOR_g keygate_XOR_102(.A(keywire176), .B(lockingkeyinput[102]), .Y(keywire130));
XOR_g keygate_XOR_104(.A(keywire178), .B(lockingkeyinput[104]), .Y(keywire147));
XOR_g keygate_XOR_105(.A(keywire179), .B(lockingkeyinput[105]), .Y(keywire133));
XOR_g keygate_XOR_106(.A(keywire180), .B(lockingkeyinput[106]), .Y(keywire123));
XOR_g keygate_XOR_109(.A(keywire183), .B(lockingkeyinput[109]), .Y(keywire87));
XOR_g keygate_XOR_110(.A(keywire184), .B(lockingkeyinput[110]), .Y(keywire119));
XOR_g keygate_XOR_111(.A(keywire185), .B(lockingkeyinput[111]), .Y(keywire79));
XOR_g keygate_XOR_113(.A(keywire187), .B(lockingkeyinput[113]), .Y(keywire134));
XOR_g keygate_XOR_115(.A(keywire189), .B(lockingkeyinput[115]), .Y(keywire150));
XOR_g keygate_XOR_117(.A(keywire191), .B(lockingkeyinput[117]), .Y(keywire88));
XOR_g keygate_XOR_119(.A(keywire193), .B(lockingkeyinput[119]), .Y(keywire80));
XOR_g keygate_XOR_121(.A(keywire195), .B(lockingkeyinput[121]), .Y(keywire117));
XOR_g keygate_XOR_124(.A(keywire198), .B(lockingkeyinput[124]), .Y(keywire81));
XOR_g keygate_XOR_127(.A(keywire201), .B(lockingkeyinput[127]), .Y(keywire115));
XOR_g keygate_XOR_130(.A(keywire204), .B(lockingkeyinput[130]), .Y(keywire96));
XOR_g keygate_XOR_133(.A(keywire207), .B(lockingkeyinput[133]), .Y(keywire112));
XOR_g keygate_XOR_134(.A(keywire208), .B(lockingkeyinput[134]), .Y(keywire116));
XOR_g keygate_XOR_136(.A(keywire210), .B(lockingkeyinput[136]), .Y(keywire188));
XOR_g keygate_XOR_137(.A(keywire211), .B(lockingkeyinput[137]), .Y(keywire175));
XOR_g keygate_XOR_139(.A(keywire213), .B(lockingkeyinput[139]), .Y(keywire164));
XOR_g keygate_XOR_140(.A(keywire214), .B(lockingkeyinput[140]), .Y(keywire161));
XOR_g keygate_XOR_145(.A(keywire219), .B(lockingkeyinput[145]), .Y(keywire158));
XOR_g keygate_XOR_146(.A(keywire220), .B(lockingkeyinput[146]), .Y(keywire84));
XOR_g keygate_XOR_158(.A(keywire232), .B(lockingkeyinput[158]), .Y(keywire204));
XOR_g keygate_XOR_161(.A(keywire235), .B(lockingkeyinput[161]), .Y(keywire99));
XOR_g keygate_XOR_166(.A(keywire240), .B(lockingkeyinput[166]), .Y(keywire190));
XOR_g keygate_XOR_167(.A(keywire241), .B(lockingkeyinput[167]), .Y(keywire105));
XOR_g keygate_XOR_171(.A(keywire245), .B(lockingkeyinput[171]), .Y(keywire194));
XOR_g keygate_XOR_175(.A(keywire249), .B(lockingkeyinput[175]), .Y(keywire197));
XOR_g keygate_XOR_176(.A(keywire250), .B(lockingkeyinput[176]), .Y(keywire205));
XOR_g keygate_XOR_177(.A(keywire251), .B(lockingkeyinput[177]), .Y(keywire201));
XOR_g keygate_XOR_178(.A(keywire252), .B(lockingkeyinput[178]), .Y(keywire208));
XOR_g keygate_XOR_183(.A(keywire257), .B(lockingkeyinput[183]), .Y(keywire173));
XOR_g keygate_XOR_184(.A(keywire258), .B(lockingkeyinput[184]), .Y(keywire177));
XOR_g keygate_XOR_185(.A(keywire259), .B(lockingkeyinput[185]), .Y(keywire180));
XOR_g keygate_XOR_186(.A(keywire260), .B(lockingkeyinput[186]), .Y(keywire124));
XOR_g keygate_XOR_187(.A(keywire261), .B(lockingkeyinput[187]), .Y(keywire125));
XOR_g keygate_XOR_188(.A(keywire262), .B(lockingkeyinput[188]), .Y(keywire126));
XOR_g keygate_XOR_190(.A(keywire264), .B(lockingkeyinput[190]), .Y(keywire160));
XOR_g keygate_XOR_191(.A(keywire265), .B(lockingkeyinput[191]), .Y(keywire172));
XOR_g keygate_XOR_192(.A(keywire266), .B(lockingkeyinput[192]), .Y(keywire176));
XOR_g keygate_XOR_193(.A(keywire267), .B(lockingkeyinput[193]), .Y(keywire131));
XOR_g keygate_XOR_194(.A(keywire268), .B(lockingkeyinput[194]), .Y(keywire132));
XOR_g keygate_XOR_199(.A(keywire273), .B(lockingkeyinput[199]), .Y(keywire137));
XOR_g keygate_XOR_204(.A(keywire278), .B(lockingkeyinput[204]), .Y(keywire142));
XOR_g keygate_XOR_205(.A(keywire279), .B(lockingkeyinput[205]), .Y(keywire143));
XOR_g keygate_XOR_207(.A(keywire281), .B(lockingkeyinput[207]), .Y(keywire145));
XOR_g keygate_XOR_208(.A(keywire282), .B(lockingkeyinput[208]), .Y(keywire146));
XOR_g keygate_XOR_210(.A(keywire284), .B(lockingkeyinput[210]), .Y(keywire186));
XOR_g keygate_XOR_213(.A(keywire287), .B(lockingkeyinput[213]), .Y(keywire167));
XOR_g keygate_XOR_214(.A(keywire288), .B(lockingkeyinput[214]), .Y(keywire169));
XOR_g keygate_XOR_216(.A(keywire290), .B(lockingkeyinput[216]), .Y(keywire170));
XOR_g keygate_XOR_220(.A(keywire294), .B(lockingkeyinput[220]), .Y(keywire219));
XOR_g keygate_XOR_221(.A(keywire295), .B(lockingkeyinput[221]), .Y(keywire264));
XOR_g keygate_XOR_222(.A(keywire296), .B(lockingkeyinput[222]), .Y(keywire214));
XOR_g keygate_XOR_223(.A(keywire297), .B(lockingkeyinput[223]), .Y(keywire238));
XOR_g keygate_XOR_224(.A(keywire298), .B(lockingkeyinput[224]), .Y(keywire292));
XOR_g keygate_XOR_226(.A(keywire300), .B(lockingkeyinput[226]), .Y(keywire213));
XOR_g keygate_XOR_227(.A(keywire301), .B(lockingkeyinput[227]), .Y(keywire222));
XOR_g keygate_XOR_229(.A(keywire303), .B(lockingkeyinput[229]), .Y(keywire287));
XOR_g keygate_XOR_230(.A(keywire304), .B(lockingkeyinput[230]), .Y(keywire212));
XOR_g keygate_XOR_231(.A(keywire305), .B(lockingkeyinput[231]), .Y(keywire288));
XOR_g keygate_XOR_232(.A(keywire306), .B(lockingkeyinput[232]), .Y(keywire290));
XOR_g keygate_XOR_234(.A(keywire308), .B(lockingkeyinput[234]), .Y(keywire265));
XOR_g keygate_XOR_235(.A(keywire309), .B(lockingkeyinput[235]), .Y(keywire257));
XOR_g keygate_XOR_237(.A(keywire311), .B(lockingkeyinput[237]), .Y(keywire211));
XOR_g keygate_XOR_239(.A(keywire313), .B(lockingkeyinput[239]), .Y(keywire258));
XOR_g keygate_XOR_240(.A(keywire314), .B(lockingkeyinput[240]), .Y(keywire283));
XOR_g keygate_XOR_241(.A(keywire315), .B(lockingkeyinput[241]), .Y(keywire269));
XOR_g keygate_XOR_244(.A(keywire318), .B(lockingkeyinput[244]), .Y(keywire239));
XOR_g keygate_XOR_245(.A(keywire319), .B(lockingkeyinput[245]), .Y(keywire223));
XOR_g keygate_XOR_246(.A(keywire320), .B(lockingkeyinput[246]), .Y(keywire255));
XOR_g keygate_XOR_247(.A(keywire321), .B(lockingkeyinput[247]), .Y(keywire215));
XOR_g keygate_XOR_249(.A(keywire323), .B(lockingkeyinput[249]), .Y(keywire270));
XOR_g keygate_XOR_250(.A(keywire324), .B(lockingkeyinput[250]), .Y(keywire210));
XOR_g keygate_XOR_251(.A(keywire325), .B(lockingkeyinput[251]), .Y(keywire286));
XOR_g keygate_XOR_252(.A(keywire326), .B(lockingkeyinput[252]), .Y(keywire240));
XOR_g keygate_XOR_253(.A(keywire327), .B(lockingkeyinput[253]), .Y(keywire224));
endmodule





module orgcir(inputs, key, out);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
input [7:0] inputs;
wire [7:0] inputs;
input [7:0] key;
wire [7:0] key;
output [1:0] out;
wire [1:0] out;
wire [4:0] scc;
wire [4:0] s1cc;
NOT_g _072_ ( .A(inputs[3]), .Y(_000_) );
XNOR_g _073_ ( .A(inputs[0]), .B(key[0]), .Y(_001_) );
XNOR_g _074_ ( .A(inputs[7]), .B(key[7]), .Y(_002_) );
AND_g _075_ ( .A(_001_), .B(_002_), .Y(_003_) );
XNOR_g _076_ ( .A(inputs[1]), .B(key[1]), .Y(_004_) );
XNOR_g _077_ ( .A(inputs[3]), .B(key[3]), .Y(_005_) );
AND_g _078_ ( .A(_004_), .B(_005_), .Y(_006_) );
AND_g _079_ ( .A(_003_), .B(_006_), .Y(_007_) );
NOR_g _080_ ( .A(inputs[5]), .B(inputs[6]), .Y(_008_) );
NOR_g _081_ ( .A(inputs[4]), .B(inputs[7]), .Y(_009_) );
AND_g _082_ ( .A(_008_), .B(_009_), .Y(_010_) );
NOR_g _083_ ( .A(inputs[1]), .B(inputs[2]), .Y(_011_) );
AND_g _084_ ( .A(inputs[0]), .B(_000_), .Y(_012_) );
AND_g _085_ ( .A(_011_), .B(_012_), .Y(_013_) );
NAND_g _086_ ( .A(_010_), .B(_013_), .Y(_014_) );
XNOR_g _087_ ( .A(inputs[5]), .B(key[5]), .Y(_015_) );
XNOR_g _088_ ( .A(inputs[2]), .B(key[2]), .Y(_016_) );
AND_g _089_ ( .A(_015_), .B(_016_), .Y(_017_) );
XNOR_g _090_ ( .A(inputs[6]), .B(key[6]), .Y(_018_) );
XNOR_g _091_ ( .A(inputs[4]), .B(key[4]), .Y(_019_) );
AND_g _092_ ( .A(_018_), .B(_019_), .Y(_020_) );
AND_g _093_ ( .A(_017_), .B(_020_), .Y(_021_) );
AND_g _094_ ( .A(_014_), .B(_021_), .Y(_022_) );
NAND_g _095_ ( .A(_007_), .B(_022_), .Y(_023_) );
XNOR_g _096_ ( .A(scc[0]), .B(_023_), .Y(out[0]) );
AND_g _097_ ( .A(inputs[0]), .B(inputs[4]), .Y(_024_) );
NAND_g _098_ ( .A(inputs[1]), .B(inputs[5]), .Y(_025_) );
XOR_g _099_ ( .A(inputs[1]), .B(inputs[5]), .Y(_026_) );
NAND_g _100_ ( .A(_024_), .B(_026_), .Y(_027_) );
XOR_g _101_ ( .A(_024_), .B(_026_), .Y(scc[1]) );
NAND_g _102_ ( .A(_025_), .B(_027_), .Y(_028_) );
NAND_g _103_ ( .A(inputs[2]), .B(inputs[6]), .Y(_029_) );
XOR_g _104_ ( .A(inputs[2]), .B(inputs[6]), .Y(_030_) );
NAND_g _105_ ( .A(_028_), .B(_030_), .Y(_031_) );
XOR_g _106_ ( .A(_028_), .B(_030_), .Y(scc[2]) );
NAND_g _107_ ( .A(_029_), .B(_031_), .Y(_032_) );
NAND_g _108_ ( .A(inputs[3]), .B(inputs[7]), .Y(_033_) );
XOR_g _109_ ( .A(inputs[3]), .B(inputs[7]), .Y(_034_) );
NAND_g _110_ ( .A(_032_), .B(_034_), .Y(_035_) );
XOR_g _111_ ( .A(_032_), .B(_034_), .Y(scc[3]) );
XOR_g _112_ ( .A(inputs[0]), .B(inputs[4]), .Y(scc[0]) );
NAND_g _113_ ( .A(_033_), .B(_035_), .Y(scc[4]) );
NOT_g _114_ ( .A(inputs[3]), .Y(_036_) );
XNOR_g _115_ ( .A(inputs[0]), .B(key[0]), .Y(_037_) );
XNOR_g _116_ ( .A(inputs[7]), .B(key[7]), .Y(_038_) );
AND_g _117_ ( .A(_037_), .B(_038_), .Y(_039_) );
XNOR_g _118_ ( .A(inputs[1]), .B(key[1]), .Y(_040_) );
XNOR_g _119_ ( .A(inputs[3]), .B(key[3]), .Y(_041_) );
AND_g _120_ ( .A(_040_), .B(_041_), .Y(_042_) );
AND_g _121_ ( .A(_039_), .B(_042_), .Y(_043_) );
NOR_g _122_ ( .A(inputs[5]), .B(inputs[6]), .Y(_044_) );
NOR_g _123_ ( .A(inputs[4]), .B(inputs[7]), .Y(_045_) );
AND_g _124_ ( .A(_044_), .B(_045_), .Y(_046_) );
NOR_g _125_ ( .A(inputs[1]), .B(inputs[2]), .Y(_047_) );
AND_g _126_ ( .A(inputs[0]), .B(_036_), .Y(_048_) );
AND_g _127_ ( .A(_047_), .B(_048_), .Y(_049_) );
NAND_g _128_ ( .A(_046_), .B(_049_), .Y(_050_) );
XNOR_g _129_ ( .A(inputs[5]), .B(key[5]), .Y(_051_) );
XNOR_g _130_ ( .A(inputs[2]), .B(key[2]), .Y(_052_) );
AND_g _131_ ( .A(_051_), .B(_052_), .Y(_053_) );
XNOR_g _132_ ( .A(inputs[6]), .B(key[6]), .Y(_054_) );
XNOR_g _133_ ( .A(inputs[4]), .B(key[4]), .Y(_055_) );
AND_g _134_ ( .A(_054_), .B(_055_), .Y(_056_) );
AND_g _135_ ( .A(_053_), .B(_056_), .Y(_057_) );
AND_g _136_ ( .A(_050_), .B(_057_), .Y(_058_) );
NAND_g _137_ ( .A(_043_), .B(_058_), .Y(_059_) );
XNOR_g _138_ ( .A(s1cc[0]), .B(_059_), .Y(out[1]) );
AND_g _139_ ( .A(inputs[0]), .B(inputs[4]), .Y(_060_) );
NAND_g _140_ ( .A(inputs[1]), .B(inputs[5]), .Y(_061_) );
XOR_g _141_ ( .A(inputs[1]), .B(inputs[5]), .Y(_062_) );
NAND_g _142_ ( .A(_060_), .B(_062_), .Y(_063_) );
XOR_g _143_ ( .A(_060_), .B(_062_), .Y(s1cc[1]) );
NAND_g _144_ ( .A(_061_), .B(_063_), .Y(_064_) );
NAND_g _145_ ( .A(inputs[2]), .B(inputs[6]), .Y(_065_) );
XOR_g _146_ ( .A(inputs[2]), .B(inputs[6]), .Y(_066_) );
NAND_g _147_ ( .A(_064_), .B(_066_), .Y(_067_) );
XOR_g _148_ ( .A(_064_), .B(_066_), .Y(s1cc[2]) );
NAND_g _149_ ( .A(_065_), .B(_067_), .Y(_068_) );
NAND_g _150_ ( .A(inputs[3]), .B(inputs[7]), .Y(_069_) );
XOR_g _151_ ( .A(inputs[3]), .B(inputs[7]), .Y(_070_) );
NAND_g _152_ ( .A(_068_), .B(_070_), .Y(_071_) );
XOR_g _153_ ( .A(_068_), .B(_070_), .Y(s1cc[3]) );
XOR_g _154_ ( .A(inputs[0]), .B(inputs[4]), .Y(s1cc[0]) );
NAND_g _155_ ( .A(_069_), .B(_071_), .Y(s1cc[4]) );
endmodule
module BUF_g(A, Y);
input A;
output Y;
assign Y=A;
endmodule

 
module NOT_g(A, Y);
input A;
output Y;
assign Y=~A;
endmodule

module AND_g(A, B, Y);
input A, B;
output Y;
assign Y=(A & B);
endmodule

module OR_g(A, B, Y);
input A, B;
output Y;
assign Y= (A | B);
endmodule

module NAND_g(A, B, Y);
input A, B;
output Y;
assign Y= ~(A & B);

endmodule

module NOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A | B);
endmodule


module XOR_g(A, B, Y);
input A, B;
output Y;
assign Y = (A ^ B);
endmodule

module XNOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A ^ B);
endmodule

module DFFcell(C, D, Q);
input C, D;
output reg Q;
always @(posedge C)
	Q <= D;
endmodule


module DFFRcell(C, D, Q, R);
input C, D, R;
output reg Q;
always @(posedge C, negedge R)
	if (!R)
		Q <= 1'b0;
	else
		Q <= D;
endmodule
