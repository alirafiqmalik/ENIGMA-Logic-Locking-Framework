module c17(N1, N2, N3, N6, N7, N22, N23);
wire _0_;
wire _1_;
wire _2_;
wire _3_;
input N1;
wire N1;
input N2;
wire N2;
output N22;
wire N22;
output N23;
wire N23;
input N3;
wire N3;
input N6;
wire N6;
input N7;
wire N7;
NAND_g _4_ ( .A(N3), .B(N6), .Y(_2_) );
NAND_g _5_ ( .A(N2), .B(_2_), .Y(_3_) );
NAND_g _6_ ( .A(N7), .B(_2_), .Y(_0_) );
NAND_g _7_ ( .A(_3_), .B(_0_), .Y(N23) );
NAND_g _8_ ( .A(N1), .B(N3), .Y(_1_) );
NAND_g _9_ ( .A(_3_), .B(_1_), .Y(N22) );
endmodule
