module picorv32(clk, resetn, trap, mem_valid, mem_instr, mem_ready, mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, irq, eoi, trace_valid, trace_data);
wire [31:0] _00000_;
wire _00001_;
wire [31:0] _00002_;
wire _00003_;
wire _00004_;
wire _00005_;
wire _00006_;
wire _00007_;
wire _00008_;
wire [31:0] _00009_;
wire [4:0] _00010_;
wire [4:0] _00011_;
wire [4:0] _00012_;
wire _00013_;
wire _00014_;
wire _00015_;
wire _00016_;
wire _00017_;
wire _00018_;
wire _00019_;
wire _00020_;
wire _00021_;
wire _00022_;
wire _00023_;
wire _00024_;
wire _00025_;
wire _00026_;
wire _00027_;
wire _00028_;
wire _00029_;
wire _00030_;
wire _00031_;
wire _00032_;
wire _00033_;
wire _00034_;
wire _00035_;
wire _00036_;
wire _00037_;
wire _00038_;
wire _00039_;
wire _00040_;
wire _00041_;
wire _00042_;
wire _00043_;
wire _00044_;
wire _00045_;
wire _00046_;
wire _00047_;
wire _00048_;
wire _00049_;
wire _00050_;
wire _00051_;
wire _00052_;
wire _00053_;
wire _00054_;
wire _00055_;
wire _00056_;
wire _00057_;
wire _00058_;
wire _00059_;
wire _00060_;
wire _00061_;
wire _00062_;
wire _00063_;
wire _00064_;
wire _00065_;
wire _00066_;
wire _00067_;
wire _00068_;
wire _00069_;
wire _00070_;
wire _00071_;
wire _00072_;
wire _00073_;
wire _00074_;
wire _00075_;
wire _00076_;
wire _00077_;
wire _00078_;
wire _00079_;
wire _00080_;
wire _00081_;
wire _00082_;
wire _00083_;
wire _00084_;
wire _00085_;
wire _00086_;
wire _00087_;
wire _00088_;
wire _00089_;
wire _00090_;
wire _00091_;
wire _00092_;
wire _00093_;
wire _00094_;
wire _00095_;
wire _00096_;
wire _00097_;
wire _00098_;
wire _00099_;
wire _00100_;
wire _00101_;
wire _00102_;
wire _00103_;
wire _00104_;
wire _00105_;
wire _00106_;
wire _00107_;
wire _00108_;
wire _00109_;
wire _00110_;
wire _00111_;
wire _00112_;
wire _00113_;
wire _00114_;
wire _00115_;
wire _00116_;
wire _00117_;
wire _00118_;
wire _00119_;
wire _00120_;
wire _00121_;
wire _00122_;
wire _00123_;
wire _00124_;
wire _00125_;
wire _00126_;
wire _00127_;
wire _00128_;
wire _00129_;
wire _00130_;
wire _00131_;
wire _00132_;
wire _00133_;
wire _00134_;
wire _00135_;
wire _00136_;
wire _00137_;
wire _00138_;
wire _00139_;
wire _00140_;
wire _00141_;
wire _00142_;
wire _00143_;
wire _00144_;
wire _00145_;
wire _00146_;
wire _00147_;
wire _00148_;
wire _00149_;
wire _00150_;
wire _00151_;
wire _00152_;
wire _00153_;
wire _00154_;
wire _00155_;
wire _00156_;
wire _00157_;
wire _00158_;
wire _00159_;
wire _00160_;
wire _00161_;
wire _00162_;
wire _00163_;
wire _00164_;
wire _00165_;
wire _00166_;
wire _00167_;
wire _00168_;
wire _00169_;
wire _00170_;
wire _00171_;
wire _00172_;
wire _00173_;
wire _00174_;
wire _00175_;
wire _00176_;
wire _00177_;
wire _00178_;
wire _00179_;
wire _00180_;
wire _00181_;
wire _00182_;
wire _00183_;
wire _00184_;
wire _00185_;
wire _00186_;
wire _00187_;
wire _00188_;
wire _00189_;
wire _00190_;
wire _00191_;
wire _00192_;
wire _00193_;
wire _00194_;
wire _00195_;
wire _00196_;
wire _00197_;
wire _00198_;
wire _00199_;
wire _00200_;
wire _00201_;
wire _00202_;
wire _00203_;
wire _00204_;
wire _00205_;
wire _00206_;
wire _00207_;
wire _00208_;
wire _00209_;
wire _00210_;
wire _00211_;
wire _00212_;
wire _00213_;
wire _00214_;
wire _00215_;
wire _00216_;
wire _00217_;
wire _00218_;
wire _00219_;
wire _00220_;
wire _00221_;
wire _00222_;
wire _00223_;
wire _00224_;
wire _00225_;
wire _00226_;
wire _00227_;
wire _00228_;
wire _00229_;
wire _00230_;
wire _00231_;
wire _00232_;
wire _00233_;
wire _00234_;
wire _00235_;
wire _00236_;
wire _00237_;
wire _00238_;
wire _00239_;
wire _00240_;
wire _00241_;
wire _00242_;
wire _00243_;
wire _00244_;
wire _00245_;
wire _00246_;
wire _00247_;
wire _00248_;
wire _00249_;
wire _00250_;
wire _00251_;
wire _00252_;
wire _00253_;
wire _00254_;
wire _00255_;
wire _00256_;
wire _00257_;
wire _00258_;
wire _00259_;
wire _00260_;
wire _00261_;
wire _00262_;
wire _00263_;
wire _00264_;
wire _00265_;
wire _00266_;
wire _00267_;
wire _00268_;
wire _00269_;
wire _00270_;
wire _00271_;
wire _00272_;
wire _00273_;
wire _00274_;
wire _00275_;
wire _00276_;
wire _00277_;
wire _00278_;
wire _00279_;
wire _00280_;
wire _00281_;
wire _00282_;
wire _00283_;
wire _00284_;
wire _00285_;
wire _00286_;
wire _00287_;
wire _00288_;
wire _00289_;
wire _00290_;
wire _00291_;
wire _00292_;
wire _00293_;
wire _00294_;
wire _00295_;
wire _00296_;
wire _00297_;
wire _00298_;
wire _00299_;
wire _00300_;
wire _00301_;
wire _00302_;
wire _00303_;
wire _00304_;
wire _00305_;
wire _00306_;
wire _00307_;
wire _00308_;
wire _00309_;
wire _00310_;
wire _00311_;
wire _00312_;
wire _00313_;
wire _00314_;
wire _00315_;
wire _00316_;
wire _00317_;
wire _00318_;
wire _00319_;
wire _00320_;
wire _00321_;
wire _00322_;
wire _00323_;
wire _00324_;
wire _00325_;
wire _00326_;
wire _00327_;
wire _00328_;
wire _00329_;
wire _00330_;
wire _00331_;
wire _00332_;
wire _00333_;
wire _00334_;
wire _00335_;
wire _00336_;
wire _00337_;
wire _00338_;
wire _00339_;
wire _00340_;
wire _00341_;
wire _00342_;
wire _00343_;
wire _00344_;
wire _00345_;
wire _00346_;
wire _00347_;
wire _00348_;
wire _00349_;
wire _00350_;
wire _00351_;
wire _00352_;
wire _00353_;
wire _00354_;
wire _00355_;
wire _00356_;
wire _00357_;
wire _00358_;
wire _00359_;
wire _00360_;
wire _00361_;
wire _00362_;
wire _00363_;
wire _00364_;
wire _00365_;
wire _00366_;
wire _00367_;
wire _00368_;
wire _00369_;
wire _00370_;
wire _00371_;
wire _00372_;
wire _00373_;
wire _00374_;
wire _00375_;
wire _00376_;
wire _00377_;
wire _00378_;
wire _00379_;
wire _00380_;
wire _00381_;
wire _00382_;
wire _00383_;
wire _00384_;
wire _00385_;
wire _00386_;
wire _00387_;
wire _00388_;
wire _00389_;
wire _00390_;
wire _00391_;
wire _00392_;
wire _00393_;
wire _00394_;
wire _00395_;
wire _00396_;
wire _00397_;
wire _00398_;
wire _00399_;
wire _00400_;
wire _00401_;
wire _00402_;
wire _00403_;
wire _00404_;
wire _00405_;
wire _00406_;
wire _00407_;
wire _00408_;
wire _00409_;
wire _00410_;
wire _00411_;
wire _00412_;
wire _00413_;
wire _00414_;
wire _00415_;
wire _00416_;
wire _00417_;
wire _00418_;
wire _00419_;
wire _00420_;
wire _00421_;
wire _00422_;
wire _00423_;
wire _00424_;
wire _00425_;
wire _00426_;
wire _00427_;
wire _00428_;
wire _00429_;
wire _00430_;
wire _00431_;
wire _00432_;
wire _00433_;
wire _00434_;
wire _00435_;
wire _00436_;
wire _00437_;
wire _00438_;
wire _00439_;
wire _00440_;
wire _00441_;
wire _00442_;
wire _00443_;
wire _00444_;
wire _00445_;
wire _00446_;
wire _00447_;
wire _00448_;
wire _00449_;
wire _00450_;
wire _00451_;
wire _00452_;
wire _00453_;
wire _00454_;
wire _00455_;
wire _00456_;
wire _00457_;
wire _00458_;
wire _00459_;
wire _00460_;
wire _00461_;
wire _00462_;
wire _00463_;
wire _00464_;
wire _00465_;
wire _00466_;
wire _00467_;
wire _00468_;
wire _00469_;
wire _00470_;
wire _00471_;
wire _00472_;
wire _00473_;
wire _00474_;
wire _00475_;
wire _00476_;
wire _00477_;
wire _00478_;
wire _00479_;
wire _00480_;
wire _00481_;
wire _00482_;
wire _00483_;
wire _00484_;
wire _00485_;
wire _00486_;
wire _00487_;
wire _00488_;
wire _00489_;
wire _00490_;
wire _00491_;
wire _00492_;
wire _00493_;
wire _00494_;
wire _00495_;
wire _00496_;
wire _00497_;
wire _00498_;
wire _00499_;
wire _00500_;
wire _00501_;
wire _00502_;
wire _00503_;
wire _00504_;
wire _00505_;
wire _00506_;
wire _00507_;
wire _00508_;
wire _00509_;
wire _00510_;
wire _00511_;
wire _00512_;
wire _00513_;
wire _00514_;
wire _00515_;
wire _00516_;
wire _00517_;
wire _00518_;
wire _00519_;
wire _00520_;
wire _00521_;
wire _00522_;
wire _00523_;
wire _00524_;
wire _00525_;
wire _00526_;
wire _00527_;
wire _00528_;
wire _00529_;
wire _00530_;
wire _00531_;
wire _00532_;
wire _00533_;
wire _00534_;
wire _00535_;
wire _00536_;
wire _00537_;
wire _00538_;
wire _00539_;
wire _00540_;
wire _00541_;
wire _00542_;
wire _00543_;
wire _00544_;
wire _00545_;
wire _00546_;
wire _00547_;
wire _00548_;
wire _00549_;
wire _00550_;
wire _00551_;
wire _00552_;
wire _00553_;
wire _00554_;
wire _00555_;
wire _00556_;
wire _00557_;
wire _00558_;
wire _00559_;
wire _00560_;
wire _00561_;
wire _00562_;
wire _00563_;
wire _00564_;
wire _00565_;
wire _00566_;
wire _00567_;
wire _00568_;
wire _00569_;
wire _00570_;
wire _00571_;
wire _00572_;
wire _00573_;
wire _00574_;
wire _00575_;
wire _00576_;
wire _00577_;
wire _00578_;
wire _00579_;
wire _00580_;
wire _00581_;
wire _00582_;
wire _00583_;
wire _00584_;
wire _00585_;
wire _00586_;
wire _00587_;
wire _00588_;
wire _00589_;
wire _00590_;
wire _00591_;
wire _00592_;
wire _00593_;
wire _00594_;
wire _00595_;
wire _00596_;
wire _00597_;
wire _00598_;
wire _00599_;
wire _00600_;
wire _00601_;
wire _00602_;
wire _00603_;
wire _00604_;
wire _00605_;
wire _00606_;
wire _00607_;
wire _00608_;
wire _00609_;
wire _00610_;
wire _00611_;
wire _00612_;
wire _00613_;
wire _00614_;
wire _00615_;
wire _00616_;
wire _00617_;
wire _00618_;
wire _00619_;
wire _00620_;
wire _00621_;
wire _00622_;
wire _00623_;
wire _00624_;
wire _00625_;
wire _00626_;
wire _00627_;
wire _00628_;
wire _00629_;
wire _00630_;
wire _00631_;
wire _00632_;
wire _00633_;
wire _00634_;
wire _00635_;
wire _00636_;
wire _00637_;
wire _00638_;
wire _00639_;
wire _00640_;
wire _00641_;
wire _00642_;
wire _00643_;
wire _00644_;
wire _00645_;
wire _00646_;
wire _00647_;
wire _00648_;
wire _00649_;
wire _00650_;
wire _00651_;
wire _00652_;
wire _00653_;
wire _00654_;
wire _00655_;
wire _00656_;
wire _00657_;
wire _00658_;
wire _00659_;
wire _00660_;
wire _00661_;
wire _00662_;
wire _00663_;
wire _00664_;
wire _00665_;
wire _00666_;
wire _00667_;
wire _00668_;
wire _00669_;
wire _00670_;
wire _00671_;
wire _00672_;
wire _00673_;
wire _00674_;
wire _00675_;
wire _00676_;
wire _00677_;
wire _00678_;
wire _00679_;
wire _00680_;
wire _00681_;
wire _00682_;
wire _00683_;
wire _00684_;
wire _00685_;
wire _00686_;
wire _00687_;
wire _00688_;
wire _00689_;
wire _00690_;
wire _00691_;
wire _00692_;
wire _00693_;
wire _00694_;
wire _00695_;
wire _00696_;
wire _00697_;
wire _00698_;
wire _00699_;
wire _00700_;
wire _00701_;
wire _00702_;
wire _00703_;
wire _00704_;
wire _00705_;
wire _00706_;
wire _00707_;
wire _00708_;
wire _00709_;
wire _00710_;
wire _00711_;
wire _00712_;
wire _00713_;
wire _00714_;
wire _00715_;
wire _00716_;
wire _00717_;
wire _00718_;
wire _00719_;
wire _00720_;
wire _00721_;
wire _00722_;
wire _00723_;
wire _00724_;
wire _00725_;
wire _00726_;
wire _00727_;
wire _00728_;
wire _00729_;
wire _00730_;
wire _00731_;
wire _00732_;
wire _00733_;
wire _00734_;
wire _00735_;
wire _00736_;
wire _00737_;
wire _00738_;
wire _00739_;
wire _00740_;
wire _00741_;
wire _00742_;
wire _00743_;
wire _00744_;
wire _00745_;
wire _00746_;
wire _00747_;
wire _00748_;
wire _00749_;
wire _00750_;
wire _00751_;
wire _00752_;
wire _00753_;
wire _00754_;
wire _00755_;
wire _00756_;
wire _00757_;
wire _00758_;
wire _00759_;
wire _00760_;
wire _00761_;
wire _00762_;
wire _00763_;
wire _00764_;
wire _00765_;
wire _00766_;
wire _00767_;
wire _00768_;
wire _00769_;
wire _00770_;
wire _00771_;
wire _00772_;
wire _00773_;
wire _00774_;
wire _00775_;
wire _00776_;
wire _00777_;
wire _00778_;
wire _00779_;
wire _00780_;
wire _00781_;
wire _00782_;
wire _00783_;
wire _00784_;
wire _00785_;
wire _00786_;
wire _00787_;
wire _00788_;
wire _00789_;
wire _00790_;
wire _00791_;
wire _00792_;
wire _00793_;
wire _00794_;
wire _00795_;
wire _00796_;
wire _00797_;
wire _00798_;
wire _00799_;
wire _00800_;
wire _00801_;
wire _00802_;
wire _00803_;
wire _00804_;
wire _00805_;
wire _00806_;
wire _00807_;
wire _00808_;
wire _00809_;
wire _00810_;
wire _00811_;
wire _00812_;
wire _00813_;
wire _00814_;
wire _00815_;
wire _00816_;
wire _00817_;
wire _00818_;
wire _00819_;
wire _00820_;
wire _00821_;
wire _00822_;
wire _00823_;
wire _00824_;
wire _00825_;
wire _00826_;
wire _00827_;
wire _00828_;
wire _00829_;
wire _00830_;
wire _00831_;
wire _00832_;
wire _00833_;
wire _00834_;
wire _00835_;
wire _00836_;
wire _00837_;
wire _00838_;
wire _00839_;
wire _00840_;
wire _00841_;
wire _00842_;
wire _00843_;
wire _00844_;
wire _00845_;
wire _00846_;
wire _00847_;
wire _00848_;
wire _00849_;
wire _00850_;
wire _00851_;
wire _00852_;
wire _00853_;
wire _00854_;
wire _00855_;
wire _00856_;
wire _00857_;
wire _00858_;
wire _00859_;
wire _00860_;
wire _00861_;
wire _00862_;
wire _00863_;
wire _00864_;
wire _00865_;
wire _00866_;
wire _00867_;
wire _00868_;
wire _00869_;
wire _00870_;
wire _00871_;
wire _00872_;
wire _00873_;
wire _00874_;
wire _00875_;
wire _00876_;
wire _00877_;
wire _00878_;
wire _00879_;
wire _00880_;
wire _00881_;
wire _00882_;
wire _00883_;
wire _00884_;
wire _00885_;
wire _00886_;
wire _00887_;
wire _00888_;
wire _00889_;
wire _00890_;
wire _00891_;
wire _00892_;
wire _00893_;
wire _00894_;
wire _00895_;
wire _00896_;
wire _00897_;
wire _00898_;
wire _00899_;
wire _00900_;
wire _00901_;
wire _00902_;
wire _00903_;
wire _00904_;
wire _00905_;
wire _00906_;
wire _00907_;
wire _00908_;
wire _00909_;
wire _00910_;
wire _00911_;
wire _00912_;
wire _00913_;
wire _00914_;
wire _00915_;
wire _00916_;
wire _00917_;
wire _00918_;
wire _00919_;
wire _00920_;
wire _00921_;
wire _00922_;
wire _00923_;
wire _00924_;
wire _00925_;
wire _00926_;
wire _00927_;
wire _00928_;
wire _00929_;
wire _00930_;
wire _00931_;
wire _00932_;
wire _00933_;
wire _00934_;
wire _00935_;
wire _00936_;
wire _00937_;
wire _00938_;
wire _00939_;
wire _00940_;
wire _00941_;
wire _00942_;
wire _00943_;
wire _00944_;
wire _00945_;
wire _00946_;
wire _00947_;
wire _00948_;
wire _00949_;
wire _00950_;
wire _00951_;
wire _00952_;
wire _00953_;
wire _00954_;
wire _00955_;
wire _00956_;
wire _00957_;
wire _00958_;
wire _00959_;
wire _00960_;
wire _00961_;
wire _00962_;
wire _00963_;
wire _00964_;
wire _00965_;
wire _00966_;
wire _00967_;
wire _00968_;
wire _00969_;
wire _00970_;
wire _00971_;
wire _00972_;
wire _00973_;
wire _00974_;
wire _00975_;
wire _00976_;
wire _00977_;
wire _00978_;
wire _00979_;
wire _00980_;
wire _00981_;
wire _00982_;
wire _00983_;
wire _00984_;
wire _00985_;
wire _00986_;
wire _00987_;
wire _00988_;
wire _00989_;
wire _00990_;
wire _00991_;
wire _00992_;
wire _00993_;
wire _00994_;
wire _00995_;
wire _00996_;
wire _00997_;
wire _00998_;
wire _00999_;
wire _01000_;
wire _01001_;
wire _01002_;
wire _01003_;
wire _01004_;
wire _01005_;
wire _01006_;
wire _01007_;
wire _01008_;
wire _01009_;
wire _01010_;
wire _01011_;
wire _01012_;
wire _01013_;
wire _01014_;
wire _01015_;
wire _01016_;
wire _01017_;
wire _01018_;
wire _01019_;
wire _01020_;
wire _01021_;
wire _01022_;
wire _01023_;
wire _01024_;
wire _01025_;
wire _01026_;
wire _01027_;
wire _01028_;
wire _01029_;
wire _01030_;
wire _01031_;
wire _01032_;
wire _01033_;
wire _01034_;
wire _01035_;
wire _01036_;
wire _01037_;
wire _01038_;
wire _01039_;
wire _01040_;
wire _01041_;
wire _01042_;
wire _01043_;
wire _01044_;
wire _01045_;
wire _01046_;
wire _01047_;
wire _01048_;
wire _01049_;
wire _01050_;
wire _01051_;
wire _01052_;
wire _01053_;
wire _01054_;
wire _01055_;
wire _01056_;
wire _01057_;
wire _01058_;
wire _01059_;
wire _01060_;
wire _01061_;
wire _01062_;
wire _01063_;
wire _01064_;
wire _01065_;
wire _01066_;
wire _01067_;
wire _01068_;
wire _01069_;
wire _01070_;
wire _01071_;
wire _01072_;
wire _01073_;
wire _01074_;
wire _01075_;
wire _01076_;
wire _01077_;
wire _01078_;
wire _01079_;
wire _01080_;
wire _01081_;
wire _01082_;
wire _01083_;
wire _01084_;
wire _01085_;
wire _01086_;
wire _01087_;
wire _01088_;
wire _01089_;
wire _01090_;
wire _01091_;
wire _01092_;
wire _01093_;
wire _01094_;
wire _01095_;
wire _01096_;
wire _01097_;
wire _01098_;
wire _01099_;
wire _01100_;
wire _01101_;
wire _01102_;
wire _01103_;
wire _01104_;
wire _01105_;
wire _01106_;
wire _01107_;
wire _01108_;
wire _01109_;
wire _01110_;
wire _01111_;
wire _01112_;
wire _01113_;
wire _01114_;
wire _01115_;
wire _01116_;
wire _01117_;
wire _01118_;
wire _01119_;
wire _01120_;
wire _01121_;
wire _01122_;
wire _01123_;
wire _01124_;
wire _01125_;
wire _01126_;
wire _01127_;
wire _01128_;
wire _01129_;
wire _01130_;
wire _01131_;
wire _01132_;
wire _01133_;
wire _01134_;
wire _01135_;
wire _01136_;
wire _01137_;
wire _01138_;
wire _01139_;
wire _01140_;
wire _01141_;
wire _01142_;
wire _01143_;
wire _01144_;
wire _01145_;
wire _01146_;
wire _01147_;
wire _01148_;
wire _01149_;
wire _01150_;
wire _01151_;
wire _01152_;
wire _01153_;
wire _01154_;
wire _01155_;
wire _01156_;
wire _01157_;
wire _01158_;
wire _01159_;
wire _01160_;
wire _01161_;
wire _01162_;
wire _01163_;
wire _01164_;
wire _01165_;
wire _01166_;
wire _01167_;
wire _01168_;
wire _01169_;
wire _01170_;
wire _01171_;
wire _01172_;
wire _01173_;
wire _01174_;
wire _01175_;
wire _01176_;
wire _01177_;
wire _01178_;
wire _01179_;
wire _01180_;
wire _01181_;
wire _01182_;
wire _01183_;
wire _01184_;
wire _01185_;
wire _01186_;
wire _01187_;
wire _01188_;
wire _01189_;
wire _01190_;
wire _01191_;
wire _01192_;
wire _01193_;
wire _01194_;
wire _01195_;
wire _01196_;
wire _01197_;
wire _01198_;
wire _01199_;
wire _01200_;
wire _01201_;
wire _01202_;
wire _01203_;
wire _01204_;
wire _01205_;
wire _01206_;
wire _01207_;
wire _01208_;
wire _01209_;
wire _01210_;
wire _01211_;
wire _01212_;
wire _01213_;
wire _01214_;
wire _01215_;
wire _01216_;
wire _01217_;
wire _01218_;
wire _01219_;
wire _01220_;
wire _01221_;
wire _01222_;
wire _01223_;
wire _01224_;
wire _01225_;
wire _01226_;
wire _01227_;
wire _01228_;
wire _01229_;
wire _01230_;
wire _01231_;
wire _01232_;
wire _01233_;
wire _01234_;
wire _01235_;
wire _01236_;
wire _01237_;
wire _01238_;
wire _01239_;
wire _01240_;
wire _01241_;
wire _01242_;
wire _01243_;
wire _01244_;
wire _01245_;
wire _01246_;
wire _01247_;
wire _01248_;
wire _01249_;
wire _01250_;
wire _01251_;
wire _01252_;
wire _01253_;
wire _01254_;
wire _01255_;
wire _01256_;
wire _01257_;
wire _01258_;
wire _01259_;
wire _01260_;
wire _01261_;
wire _01262_;
wire _01263_;
wire _01264_;
wire _01265_;
wire _01266_;
wire _01267_;
wire _01268_;
wire _01269_;
wire _01270_;
wire _01271_;
wire _01272_;
wire _01273_;
wire _01274_;
wire _01275_;
wire _01276_;
wire _01277_;
wire _01278_;
wire _01279_;
wire _01280_;
wire _01281_;
wire _01282_;
wire _01283_;
wire _01284_;
wire _01285_;
wire _01286_;
wire _01287_;
wire _01288_;
wire _01289_;
wire _01290_;
wire _01291_;
wire _01292_;
wire _01293_;
wire _01294_;
wire _01295_;
wire _01296_;
wire _01297_;
wire _01298_;
wire _01299_;
wire _01300_;
wire _01301_;
wire _01302_;
wire _01303_;
wire _01304_;
wire _01305_;
wire _01306_;
wire _01307_;
wire _01308_;
wire _01309_;
wire _01310_;
wire _01311_;
wire _01312_;
wire _01313_;
wire _01314_;
wire _01315_;
wire _01316_;
wire _01317_;
wire _01318_;
wire _01319_;
wire _01320_;
wire _01321_;
wire _01322_;
wire _01323_;
wire _01324_;
wire _01325_;
wire _01326_;
wire _01327_;
wire _01328_;
wire _01329_;
wire _01330_;
wire _01331_;
wire _01332_;
wire _01333_;
wire _01334_;
wire _01335_;
wire _01336_;
wire _01337_;
wire _01338_;
wire _01339_;
wire _01340_;
wire _01341_;
wire _01342_;
wire _01343_;
wire _01344_;
wire _01345_;
wire _01346_;
wire _01347_;
wire _01348_;
wire _01349_;
wire _01350_;
wire _01351_;
wire _01352_;
wire _01353_;
wire _01354_;
wire _01355_;
wire _01356_;
wire _01357_;
wire _01358_;
wire _01359_;
wire _01360_;
wire _01361_;
wire _01362_;
wire _01363_;
wire _01364_;
wire _01365_;
wire _01366_;
wire _01367_;
wire _01368_;
wire _01369_;
wire _01370_;
wire _01371_;
wire _01372_;
wire _01373_;
wire _01374_;
wire _01375_;
wire _01376_;
wire _01377_;
wire _01378_;
wire _01379_;
wire _01380_;
wire _01381_;
wire _01382_;
wire _01383_;
wire _01384_;
wire _01385_;
wire _01386_;
wire _01387_;
wire _01388_;
wire _01389_;
wire _01390_;
wire _01391_;
wire _01392_;
wire _01393_;
wire _01394_;
wire _01395_;
wire _01396_;
wire _01397_;
wire _01398_;
wire _01399_;
wire _01400_;
wire _01401_;
wire _01402_;
wire _01403_;
wire _01404_;
wire _01405_;
wire _01406_;
wire _01407_;
wire _01408_;
wire _01409_;
wire _01410_;
wire _01411_;
wire _01412_;
wire _01413_;
wire _01414_;
wire _01415_;
wire _01416_;
wire _01417_;
wire _01418_;
wire _01419_;
wire _01420_;
wire _01421_;
wire _01422_;
wire _01423_;
wire _01424_;
wire _01425_;
wire _01426_;
wire _01427_;
wire _01428_;
wire _01429_;
wire _01430_;
wire _01431_;
wire _01432_;
wire _01433_;
wire _01434_;
wire _01435_;
wire _01436_;
wire _01437_;
wire _01438_;
wire _01439_;
wire _01440_;
wire _01441_;
wire _01442_;
wire _01443_;
wire _01444_;
wire _01445_;
wire _01446_;
wire _01447_;
wire _01448_;
wire _01449_;
wire _01450_;
wire _01451_;
wire _01452_;
wire _01453_;
wire _01454_;
wire _01455_;
wire _01456_;
wire _01457_;
wire _01458_;
wire _01459_;
wire _01460_;
wire _01461_;
wire _01462_;
wire _01463_;
wire _01464_;
wire _01465_;
wire _01466_;
wire _01467_;
wire _01468_;
wire _01469_;
wire _01470_;
wire _01471_;
wire _01472_;
wire _01473_;
wire _01474_;
wire _01475_;
wire _01476_;
wire _01477_;
wire _01478_;
wire _01479_;
wire _01480_;
wire _01481_;
wire _01482_;
wire _01483_;
wire _01484_;
wire _01485_;
wire _01486_;
wire _01487_;
wire _01488_;
wire _01489_;
wire _01490_;
wire _01491_;
wire _01492_;
wire _01493_;
wire _01494_;
wire _01495_;
wire _01496_;
wire _01497_;
wire _01498_;
wire _01499_;
wire _01500_;
wire _01501_;
wire _01502_;
wire _01503_;
wire _01504_;
wire _01505_;
wire _01506_;
wire _01507_;
wire _01508_;
wire _01509_;
wire _01510_;
wire _01511_;
wire _01512_;
wire _01513_;
wire _01514_;
wire _01515_;
wire _01516_;
wire _01517_;
wire _01518_;
wire _01519_;
wire _01520_;
wire _01521_;
wire _01522_;
wire _01523_;
wire _01524_;
wire _01525_;
wire _01526_;
wire _01527_;
wire _01528_;
wire _01529_;
wire _01530_;
wire _01531_;
wire _01532_;
wire _01533_;
wire _01534_;
wire _01535_;
wire _01536_;
wire _01537_;
wire _01538_;
wire _01539_;
wire _01540_;
wire _01541_;
wire _01542_;
wire _01543_;
wire _01544_;
wire _01545_;
wire _01546_;
wire _01547_;
wire _01548_;
wire _01549_;
wire _01550_;
wire _01551_;
wire _01552_;
wire _01553_;
wire _01554_;
wire _01555_;
wire _01556_;
wire _01557_;
wire _01558_;
wire _01559_;
wire _01560_;
wire _01561_;
wire _01562_;
wire _01563_;
wire _01564_;
wire _01565_;
wire _01566_;
wire _01567_;
wire _01568_;
wire _01569_;
wire _01570_;
wire _01571_;
wire _01572_;
wire _01573_;
wire _01574_;
wire _01575_;
wire _01576_;
wire _01577_;
wire _01578_;
wire _01579_;
wire _01580_;
wire _01581_;
wire _01582_;
wire _01583_;
wire _01584_;
wire _01585_;
wire _01586_;
wire _01587_;
wire _01588_;
wire _01589_;
wire _01590_;
wire _01591_;
wire _01592_;
wire _01593_;
wire _01594_;
wire _01595_;
wire _01596_;
wire _01597_;
wire _01598_;
wire _01599_;
wire _01600_;
wire _01601_;
wire _01602_;
wire _01603_;
wire _01604_;
wire _01605_;
wire _01606_;
wire _01607_;
wire _01608_;
wire _01609_;
wire _01610_;
wire _01611_;
wire _01612_;
wire _01613_;
wire _01614_;
wire _01615_;
wire _01616_;
wire _01617_;
wire _01618_;
wire _01619_;
wire _01620_;
wire _01621_;
wire _01622_;
wire _01623_;
wire _01624_;
wire _01625_;
wire _01626_;
wire _01627_;
wire _01628_;
wire _01629_;
wire _01630_;
wire _01631_;
wire _01632_;
wire _01633_;
wire _01634_;
wire _01635_;
wire _01636_;
wire _01637_;
wire _01638_;
wire _01639_;
wire _01640_;
wire _01641_;
wire _01642_;
wire _01643_;
wire _01644_;
wire _01645_;
wire _01646_;
wire _01647_;
wire _01648_;
wire _01649_;
wire _01650_;
wire _01651_;
wire _01652_;
wire _01653_;
wire _01654_;
wire _01655_;
wire _01656_;
wire _01657_;
wire _01658_;
wire _01659_;
wire _01660_;
wire _01661_;
wire _01662_;
wire _01663_;
wire _01664_;
wire _01665_;
wire _01666_;
wire _01667_;
wire _01668_;
wire _01669_;
wire _01670_;
wire _01671_;
wire _01672_;
wire _01673_;
wire _01674_;
wire _01675_;
wire _01676_;
wire _01677_;
wire _01678_;
wire _01679_;
wire _01680_;
wire _01681_;
wire _01682_;
wire _01683_;
wire _01684_;
wire _01685_;
wire _01686_;
wire _01687_;
wire _01688_;
wire _01689_;
wire _01690_;
wire _01691_;
wire _01692_;
wire _01693_;
wire _01694_;
wire _01695_;
wire _01696_;
wire _01697_;
wire _01698_;
wire _01699_;
wire _01700_;
wire _01701_;
wire _01702_;
wire _01703_;
wire _01704_;
wire _01705_;
wire _01706_;
wire _01707_;
wire _01708_;
wire _01709_;
wire _01710_;
wire _01711_;
wire _01712_;
wire _01713_;
wire _01714_;
wire _01715_;
wire _01716_;
wire _01717_;
wire _01718_;
wire _01719_;
wire _01720_;
wire _01721_;
wire _01722_;
wire _01723_;
wire _01724_;
wire _01725_;
wire _01726_;
wire _01727_;
wire _01728_;
wire _01729_;
wire _01730_;
wire _01731_;
wire _01732_;
wire _01733_;
wire _01734_;
wire _01735_;
wire _01736_;
wire _01737_;
wire _01738_;
wire _01739_;
wire _01740_;
wire _01741_;
wire _01742_;
wire _01743_;
wire _01744_;
wire _01745_;
wire _01746_;
wire _01747_;
wire _01748_;
wire _01749_;
wire _01750_;
wire _01751_;
wire _01752_;
wire _01753_;
wire _01754_;
wire _01755_;
wire _01756_;
wire _01757_;
wire _01758_;
wire _01759_;
wire _01760_;
wire _01761_;
wire _01762_;
wire _01763_;
wire _01764_;
wire _01765_;
wire _01766_;
wire _01767_;
wire _01768_;
wire _01769_;
wire _01770_;
wire _01771_;
wire _01772_;
wire _01773_;
wire _01774_;
wire _01775_;
wire _01776_;
wire _01777_;
wire _01778_;
wire _01779_;
wire _01780_;
wire _01781_;
wire _01782_;
wire _01783_;
wire _01784_;
wire _01785_;
wire _01786_;
wire _01787_;
wire _01788_;
wire _01789_;
wire _01790_;
wire _01791_;
wire _01792_;
wire _01793_;
wire _01794_;
wire _01795_;
wire _01796_;
wire _01797_;
wire _01798_;
wire _01799_;
wire _01800_;
wire _01801_;
wire _01802_;
wire _01803_;
wire _01804_;
wire _01805_;
wire _01806_;
wire _01807_;
wire _01808_;
wire _01809_;
wire _01810_;
wire _01811_;
wire _01812_;
wire _01813_;
wire _01814_;
wire _01815_;
wire _01816_;
wire _01817_;
wire _01818_;
wire _01819_;
wire _01820_;
wire _01821_;
wire _01822_;
wire _01823_;
wire _01824_;
wire _01825_;
wire _01826_;
wire _01827_;
wire _01828_;
wire _01829_;
wire _01830_;
wire _01831_;
wire _01832_;
wire _01833_;
wire _01834_;
wire _01835_;
wire _01836_;
wire _01837_;
wire _01838_;
wire _01839_;
wire _01840_;
wire _01841_;
wire _01842_;
wire _01843_;
wire _01844_;
wire _01845_;
wire _01846_;
wire _01847_;
wire _01848_;
wire _01849_;
wire _01850_;
wire _01851_;
wire _01852_;
wire _01853_;
wire _01854_;
wire _01855_;
wire _01856_;
wire _01857_;
wire _01858_;
wire _01859_;
wire _01860_;
wire _01861_;
wire _01862_;
wire _01863_;
wire _01864_;
wire _01865_;
wire _01866_;
wire _01867_;
wire _01868_;
wire _01869_;
wire _01870_;
wire _01871_;
wire _01872_;
wire _01873_;
wire _01874_;
wire _01875_;
wire _01876_;
wire _01877_;
wire _01878_;
wire _01879_;
wire _01880_;
wire _01881_;
wire _01882_;
wire _01883_;
wire _01884_;
wire _01885_;
wire _01886_;
wire _01887_;
wire _01888_;
wire _01889_;
wire _01890_;
wire _01891_;
wire _01892_;
wire _01893_;
wire _01894_;
wire _01895_;
wire _01896_;
wire _01897_;
wire _01898_;
wire _01899_;
wire _01900_;
wire _01901_;
wire _01902_;
wire _01903_;
wire _01904_;
wire _01905_;
wire _01906_;
wire _01907_;
wire _01908_;
wire _01909_;
wire _01910_;
wire _01911_;
wire _01912_;
wire _01913_;
wire _01914_;
wire _01915_;
wire _01916_;
wire _01917_;
wire _01918_;
wire _01919_;
wire _01920_;
wire _01921_;
wire _01922_;
wire _01923_;
wire _01924_;
wire _01925_;
wire _01926_;
wire _01927_;
wire _01928_;
wire _01929_;
wire _01930_;
wire _01931_;
wire _01932_;
wire _01933_;
wire _01934_;
wire _01935_;
wire _01936_;
wire _01937_;
wire _01938_;
wire _01939_;
wire _01940_;
wire _01941_;
wire _01942_;
wire _01943_;
wire _01944_;
wire _01945_;
wire _01946_;
wire _01947_;
wire _01948_;
wire _01949_;
wire _01950_;
wire _01951_;
wire _01952_;
wire _01953_;
wire _01954_;
wire _01955_;
wire _01956_;
wire _01957_;
wire _01958_;
wire _01959_;
wire _01960_;
wire _01961_;
wire _01962_;
wire _01963_;
wire _01964_;
wire _01965_;
wire _01966_;
wire _01967_;
wire _01968_;
wire _01969_;
wire _01970_;
wire _01971_;
wire _01972_;
wire _01973_;
wire _01974_;
wire _01975_;
wire _01976_;
wire _01977_;
wire _01978_;
wire _01979_;
wire _01980_;
wire _01981_;
wire _01982_;
wire _01983_;
wire _01984_;
wire _01985_;
wire _01986_;
wire _01987_;
wire _01988_;
wire _01989_;
wire _01990_;
wire _01991_;
wire _01992_;
wire _01993_;
wire _01994_;
wire _01995_;
wire _01996_;
wire _01997_;
wire _01998_;
wire _01999_;
wire _02000_;
wire _02001_;
wire _02002_;
wire _02003_;
wire _02004_;
wire _02005_;
wire _02006_;
wire _02007_;
wire _02008_;
wire _02009_;
wire _02010_;
wire _02011_;
wire _02012_;
wire _02013_;
wire _02014_;
wire _02015_;
wire _02016_;
wire _02017_;
wire _02018_;
wire _02019_;
wire _02020_;
wire _02021_;
wire _02022_;
wire _02023_;
wire _02024_;
wire _02025_;
wire _02026_;
wire _02027_;
wire _02028_;
wire _02029_;
wire _02030_;
wire _02031_;
wire _02032_;
wire _02033_;
wire _02034_;
wire _02035_;
wire _02036_;
wire _02037_;
wire _02038_;
wire _02039_;
wire _02040_;
wire _02041_;
wire _02042_;
wire _02043_;
wire _02044_;
wire _02045_;
wire _02046_;
wire _02047_;
wire _02048_;
wire _02049_;
wire _02050_;
wire _02051_;
wire _02052_;
wire _02053_;
wire _02054_;
wire _02055_;
wire _02056_;
wire _02057_;
wire _02058_;
wire _02059_;
wire _02060_;
wire _02061_;
wire _02062_;
wire _02063_;
wire _02064_;
wire _02065_;
wire _02066_;
wire _02067_;
wire _02068_;
wire _02069_;
wire _02070_;
wire _02071_;
wire _02072_;
wire _02073_;
wire _02074_;
wire _02075_;
wire _02076_;
wire _02077_;
wire _02078_;
wire _02079_;
wire _02080_;
wire _02081_;
wire _02082_;
wire _02083_;
wire _02084_;
wire _02085_;
wire _02086_;
wire _02087_;
wire _02088_;
wire _02089_;
wire _02090_;
wire _02091_;
wire _02092_;
wire _02093_;
wire _02094_;
wire _02095_;
wire _02096_;
wire _02097_;
wire _02098_;
wire _02099_;
wire _02100_;
wire _02101_;
wire _02102_;
wire _02103_;
wire _02104_;
wire _02105_;
wire _02106_;
wire _02107_;
wire _02108_;
wire _02109_;
wire _02110_;
wire _02111_;
wire _02112_;
wire _02113_;
wire _02114_;
wire _02115_;
wire _02116_;
wire _02117_;
wire _02118_;
wire _02119_;
wire _02120_;
wire _02121_;
wire _02122_;
wire _02123_;
wire _02124_;
wire _02125_;
wire _02126_;
wire _02127_;
wire _02128_;
wire _02129_;
wire _02130_;
wire _02131_;
wire _02132_;
wire _02133_;
wire _02134_;
wire _02135_;
wire _02136_;
wire _02137_;
wire _02138_;
wire _02139_;
wire _02140_;
wire _02141_;
wire _02142_;
wire _02143_;
wire _02144_;
wire _02145_;
wire _02146_;
wire _02147_;
wire _02148_;
wire _02149_;
wire _02150_;
wire _02151_;
wire _02152_;
wire _02153_;
wire _02154_;
wire _02155_;
wire _02156_;
wire _02157_;
wire _02158_;
wire _02159_;
wire _02160_;
wire _02161_;
wire _02162_;
wire _02163_;
wire _02164_;
wire _02165_;
wire _02166_;
wire _02167_;
wire _02168_;
wire _02169_;
wire _02170_;
wire _02171_;
wire _02172_;
wire _02173_;
wire _02174_;
wire _02175_;
wire _02176_;
wire _02177_;
wire _02178_;
wire _02179_;
wire _02180_;
wire _02181_;
wire _02182_;
wire _02183_;
wire _02184_;
wire _02185_;
wire _02186_;
wire _02187_;
wire _02188_;
wire _02189_;
wire _02190_;
wire _02191_;
wire _02192_;
wire _02193_;
wire _02194_;
wire _02195_;
wire _02196_;
wire _02197_;
wire _02198_;
wire _02199_;
wire _02200_;
wire _02201_;
wire _02202_;
wire _02203_;
wire _02204_;
wire _02205_;
wire _02206_;
wire _02207_;
wire _02208_;
wire _02209_;
wire _02210_;
wire _02211_;
wire _02212_;
wire _02213_;
wire _02214_;
wire _02215_;
wire _02216_;
wire _02217_;
wire _02218_;
wire _02219_;
wire _02220_;
wire _02221_;
wire _02222_;
wire _02223_;
wire _02224_;
wire _02225_;
wire _02226_;
wire _02227_;
wire _02228_;
wire _02229_;
wire _02230_;
wire _02231_;
wire _02232_;
wire _02233_;
wire _02234_;
wire _02235_;
wire _02236_;
wire _02237_;
wire _02238_;
wire _02239_;
wire _02240_;
wire _02241_;
wire _02242_;
wire _02243_;
wire _02244_;
wire _02245_;
wire _02246_;
wire _02247_;
wire _02248_;
wire _02249_;
wire _02250_;
wire _02251_;
wire _02252_;
wire _02253_;
wire _02254_;
wire _02255_;
wire _02256_;
wire _02257_;
wire _02258_;
wire _02259_;
wire _02260_;
wire _02261_;
wire _02262_;
wire _02263_;
wire _02264_;
wire _02265_;
wire _02266_;
wire _02267_;
wire _02268_;
wire _02269_;
wire _02270_;
wire _02271_;
wire _02272_;
wire _02273_;
wire _02274_;
wire _02275_;
wire _02276_;
wire _02277_;
wire _02278_;
wire _02279_;
wire _02280_;
wire _02281_;
wire _02282_;
wire _02283_;
wire _02284_;
wire _02285_;
wire _02286_;
wire _02287_;
wire _02288_;
wire _02289_;
wire _02290_;
wire _02291_;
wire _02292_;
wire _02293_;
wire _02294_;
wire _02295_;
wire _02296_;
wire _02297_;
wire _02298_;
wire _02299_;
wire _02300_;
wire _02301_;
wire _02302_;
wire _02303_;
wire _02304_;
wire _02305_;
wire _02306_;
wire _02307_;
wire _02308_;
wire _02309_;
wire _02310_;
wire _02311_;
wire _02312_;
wire _02313_;
wire _02314_;
wire _02315_;
wire _02316_;
wire _02317_;
wire _02318_;
wire _02319_;
wire _02320_;
wire _02321_;
wire _02322_;
wire _02323_;
wire _02324_;
wire _02325_;
wire _02326_;
wire _02327_;
wire _02328_;
wire _02329_;
wire _02330_;
wire _02331_;
wire _02332_;
wire _02333_;
wire _02334_;
wire _02335_;
wire _02336_;
wire _02337_;
wire _02338_;
wire _02339_;
wire _02340_;
wire _02341_;
wire _02342_;
wire _02343_;
wire _02344_;
wire _02345_;
wire _02346_;
wire _02347_;
wire _02348_;
wire _02349_;
wire _02350_;
wire _02351_;
wire _02352_;
wire _02353_;
wire _02354_;
wire _02355_;
wire _02356_;
wire _02357_;
wire _02358_;
wire _02359_;
wire _02360_;
wire _02361_;
wire _02362_;
wire _02363_;
wire _02364_;
wire _02365_;
wire _02366_;
wire _02367_;
wire _02368_;
wire _02369_;
wire _02370_;
wire _02371_;
wire _02372_;
wire _02373_;
wire _02374_;
wire _02375_;
wire _02376_;
wire _02377_;
wire _02378_;
wire _02379_;
wire _02380_;
wire _02381_;
wire _02382_;
wire _02383_;
wire _02384_;
wire _02385_;
wire _02386_;
wire _02387_;
wire _02388_;
wire _02389_;
wire _02390_;
wire _02391_;
wire _02392_;
wire _02393_;
wire _02394_;
wire _02395_;
wire _02396_;
wire _02397_;
wire _02398_;
wire _02399_;
wire _02400_;
wire _02401_;
wire _02402_;
wire _02403_;
wire _02404_;
wire _02405_;
wire _02406_;
wire _02407_;
wire _02408_;
wire _02409_;
wire _02410_;
wire _02411_;
wire _02412_;
wire _02413_;
wire _02414_;
wire _02415_;
wire _02416_;
wire _02417_;
wire _02418_;
wire _02419_;
wire _02420_;
wire _02421_;
wire _02422_;
wire _02423_;
wire _02424_;
wire _02425_;
wire _02426_;
wire _02427_;
wire _02428_;
wire _02429_;
wire _02430_;
wire _02431_;
wire _02432_;
wire _02433_;
wire _02434_;
wire _02435_;
wire _02436_;
wire _02437_;
wire _02438_;
wire _02439_;
wire _02440_;
wire _02441_;
wire _02442_;
wire _02443_;
wire _02444_;
wire _02445_;
wire _02446_;
wire _02447_;
wire _02448_;
wire _02449_;
wire _02450_;
wire _02451_;
wire _02452_;
wire _02453_;
wire _02454_;
wire _02455_;
wire _02456_;
wire _02457_;
wire _02458_;
wire _02459_;
wire _02460_;
wire _02461_;
wire _02462_;
wire _02463_;
wire _02464_;
wire _02465_;
wire _02466_;
wire _02467_;
wire _02468_;
wire _02469_;
wire _02470_;
wire _02471_;
wire _02472_;
wire _02473_;
wire _02474_;
wire _02475_;
wire _02476_;
wire _02477_;
wire _02478_;
wire _02479_;
wire _02480_;
wire _02481_;
wire _02482_;
wire _02483_;
wire _02484_;
wire _02485_;
wire _02486_;
wire _02487_;
wire _02488_;
wire _02489_;
wire _02490_;
wire _02491_;
wire _02492_;
wire _02493_;
wire _02494_;
wire _02495_;
wire _02496_;
wire _02497_;
wire _02498_;
wire _02499_;
wire _02500_;
wire _02501_;
wire _02502_;
wire _02503_;
wire _02504_;
wire _02505_;
wire _02506_;
wire _02507_;
wire _02508_;
wire _02509_;
wire _02510_;
wire _02511_;
wire _02512_;
wire _02513_;
wire _02514_;
wire _02515_;
wire _02516_;
wire _02517_;
wire _02518_;
wire _02519_;
wire _02520_;
wire _02521_;
wire _02522_;
wire _02523_;
wire _02524_;
wire _02525_;
wire _02526_;
wire _02527_;
wire _02528_;
wire _02529_;
wire _02530_;
wire _02531_;
wire _02532_;
wire _02533_;
wire _02534_;
wire _02535_;
wire _02536_;
wire _02537_;
wire _02538_;
wire _02539_;
wire _02540_;
wire _02541_;
wire _02542_;
wire _02543_;
wire _02544_;
wire _02545_;
wire _02546_;
wire _02547_;
wire _02548_;
wire _02549_;
wire _02550_;
wire _02551_;
wire _02552_;
wire _02553_;
wire _02554_;
wire _02555_;
wire _02556_;
wire _02557_;
wire _02558_;
wire _02559_;
wire _02560_;
wire _02561_;
wire _02562_;
wire _02563_;
wire _02564_;
wire _02565_;
wire _02566_;
wire _02567_;
wire _02568_;
wire _02569_;
wire _02570_;
wire _02571_;
wire _02572_;
wire _02573_;
wire _02574_;
wire _02575_;
wire _02576_;
wire _02577_;
wire _02578_;
wire _02579_;
wire _02580_;
wire _02581_;
wire _02582_;
wire _02583_;
wire _02584_;
wire _02585_;
wire _02586_;
wire _02587_;
wire _02588_;
wire _02589_;
wire _02590_;
wire _02591_;
wire _02592_;
wire _02593_;
wire _02594_;
wire _02595_;
wire _02596_;
wire _02597_;
wire _02598_;
wire _02599_;
wire _02600_;
wire _02601_;
wire _02602_;
wire _02603_;
wire _02604_;
wire _02605_;
wire _02606_;
wire _02607_;
wire _02608_;
wire _02609_;
wire _02610_;
wire _02611_;
wire _02612_;
wire _02613_;
wire _02614_;
wire _02615_;
wire _02616_;
wire _02617_;
wire _02618_;
wire _02619_;
wire _02620_;
wire _02621_;
wire _02622_;
wire _02623_;
wire _02624_;
wire _02625_;
wire _02626_;
wire _02627_;
wire _02628_;
wire _02629_;
wire _02630_;
wire _02631_;
wire _02632_;
wire _02633_;
wire _02634_;
wire _02635_;
wire _02636_;
wire _02637_;
wire _02638_;
wire _02639_;
wire _02640_;
wire _02641_;
wire _02642_;
wire _02643_;
wire _02644_;
wire _02645_;
wire _02646_;
wire _02647_;
wire _02648_;
wire _02649_;
wire _02650_;
wire _02651_;
wire _02652_;
wire _02653_;
wire _02654_;
wire _02655_;
wire _02656_;
wire _02657_;
wire _02658_;
wire _02659_;
wire _02660_;
wire _02661_;
wire _02662_;
wire _02663_;
wire _02664_;
wire _02665_;
wire _02666_;
wire _02667_;
wire _02668_;
wire _02669_;
wire _02670_;
wire _02671_;
wire _02672_;
wire _02673_;
wire _02674_;
wire _02675_;
wire _02676_;
wire _02677_;
wire _02678_;
wire _02679_;
wire _02680_;
wire _02681_;
wire _02682_;
wire _02683_;
wire _02684_;
wire _02685_;
wire _02686_;
wire _02687_;
wire _02688_;
wire _02689_;
wire _02690_;
wire _02691_;
wire _02692_;
wire _02693_;
wire _02694_;
wire _02695_;
wire _02696_;
wire _02697_;
wire _02698_;
wire _02699_;
wire _02700_;
wire _02701_;
wire _02702_;
wire _02703_;
wire _02704_;
wire _02705_;
wire _02706_;
wire _02707_;
wire _02708_;
wire _02709_;
wire _02710_;
wire _02711_;
wire _02712_;
wire _02713_;
wire _02714_;
wire _02715_;
wire _02716_;
wire _02717_;
wire _02718_;
wire _02719_;
wire _02720_;
wire _02721_;
wire _02722_;
wire _02723_;
wire _02724_;
wire _02725_;
wire _02726_;
wire _02727_;
wire _02728_;
wire _02729_;
wire _02730_;
wire _02731_;
wire _02732_;
wire _02733_;
wire _02734_;
wire _02735_;
wire _02736_;
wire _02737_;
wire _02738_;
wire _02739_;
wire _02740_;
wire _02741_;
wire _02742_;
wire _02743_;
wire _02744_;
wire _02745_;
wire _02746_;
wire _02747_;
wire _02748_;
wire _02749_;
wire _02750_;
wire _02751_;
wire _02752_;
wire _02753_;
wire _02754_;
wire _02755_;
wire _02756_;
wire _02757_;
wire _02758_;
wire _02759_;
wire _02760_;
wire _02761_;
wire _02762_;
wire _02763_;
wire _02764_;
wire _02765_;
wire _02766_;
wire _02767_;
wire _02768_;
wire _02769_;
wire _02770_;
wire _02771_;
wire _02772_;
wire _02773_;
wire _02774_;
wire _02775_;
wire _02776_;
wire _02777_;
wire _02778_;
wire _02779_;
wire _02780_;
wire _02781_;
wire _02782_;
wire _02783_;
wire _02784_;
wire _02785_;
wire _02786_;
wire _02787_;
wire _02788_;
wire _02789_;
wire _02790_;
wire _02791_;
wire _02792_;
wire _02793_;
wire _02794_;
wire _02795_;
wire _02796_;
wire _02797_;
wire _02798_;
wire _02799_;
wire _02800_;
wire _02801_;
wire _02802_;
wire _02803_;
wire _02804_;
wire _02805_;
wire _02806_;
wire _02807_;
wire _02808_;
wire _02809_;
wire _02810_;
wire _02811_;
wire _02812_;
wire _02813_;
wire _02814_;
wire _02815_;
wire _02816_;
wire _02817_;
wire _02818_;
wire _02819_;
wire _02820_;
wire _02821_;
wire _02822_;
wire _02823_;
wire _02824_;
wire _02825_;
wire _02826_;
wire _02827_;
wire _02828_;
wire _02829_;
wire _02830_;
wire _02831_;
wire _02832_;
wire _02833_;
wire _02834_;
wire _02835_;
wire _02836_;
wire _02837_;
wire _02838_;
wire _02839_;
wire _02840_;
wire _02841_;
wire _02842_;
wire _02843_;
wire _02844_;
wire _02845_;
wire _02846_;
wire _02847_;
wire _02848_;
wire _02849_;
wire _02850_;
wire _02851_;
wire _02852_;
wire _02853_;
wire _02854_;
wire _02855_;
wire _02856_;
wire _02857_;
wire _02858_;
wire _02859_;
wire _02860_;
wire _02861_;
wire _02862_;
wire _02863_;
wire _02864_;
wire _02865_;
wire _02866_;
wire _02867_;
wire _02868_;
wire _02869_;
wire _02870_;
wire _02871_;
wire _02872_;
wire _02873_;
wire _02874_;
wire _02875_;
wire _02876_;
wire _02877_;
wire _02878_;
wire _02879_;
wire _02880_;
wire _02881_;
wire _02882_;
wire _02883_;
wire _02884_;
wire _02885_;
wire _02886_;
wire _02887_;
wire _02888_;
wire _02889_;
wire _02890_;
wire _02891_;
wire _02892_;
wire _02893_;
wire _02894_;
wire _02895_;
wire _02896_;
wire _02897_;
wire _02898_;
wire _02899_;
wire _02900_;
wire _02901_;
wire _02902_;
wire _02903_;
wire _02904_;
wire _02905_;
wire _02906_;
wire _02907_;
wire _02908_;
wire _02909_;
wire _02910_;
wire _02911_;
wire _02912_;
wire _02913_;
wire _02914_;
wire _02915_;
wire _02916_;
wire _02917_;
wire _02918_;
wire _02919_;
wire _02920_;
wire _02921_;
wire _02922_;
wire _02923_;
wire _02924_;
wire _02925_;
wire _02926_;
wire _02927_;
wire _02928_;
wire _02929_;
wire _02930_;
wire _02931_;
wire _02932_;
wire _02933_;
wire _02934_;
wire _02935_;
wire _02936_;
wire _02937_;
wire _02938_;
wire _02939_;
wire _02940_;
wire _02941_;
wire _02942_;
wire _02943_;
wire _02944_;
wire _02945_;
wire _02946_;
wire _02947_;
wire _02948_;
wire _02949_;
wire _02950_;
wire _02951_;
wire _02952_;
wire _02953_;
wire _02954_;
wire _02955_;
wire _02956_;
wire _02957_;
wire _02958_;
wire _02959_;
wire _02960_;
wire _02961_;
wire _02962_;
wire _02963_;
wire _02964_;
wire _02965_;
wire _02966_;
wire _02967_;
wire _02968_;
wire _02969_;
wire _02970_;
wire _02971_;
wire _02972_;
wire _02973_;
wire _02974_;
wire _02975_;
wire _02976_;
wire _02977_;
wire _02978_;
wire _02979_;
wire _02980_;
wire _02981_;
wire _02982_;
wire _02983_;
wire _02984_;
wire _02985_;
wire _02986_;
wire _02987_;
wire _02988_;
wire _02989_;
wire _02990_;
wire _02991_;
wire _02992_;
wire _02993_;
wire _02994_;
wire _02995_;
wire _02996_;
wire _02997_;
wire _02998_;
wire _02999_;
wire _03000_;
wire _03001_;
wire _03002_;
wire _03003_;
wire _03004_;
wire _03005_;
wire _03006_;
wire _03007_;
wire _03008_;
wire _03009_;
wire _03010_;
wire _03011_;
wire _03012_;
wire _03013_;
wire _03014_;
wire _03015_;
wire _03016_;
wire _03017_;
wire _03018_;
wire _03019_;
wire _03020_;
wire _03021_;
wire _03022_;
wire _03023_;
wire _03024_;
wire _03025_;
wire _03026_;
wire _03027_;
wire _03028_;
wire _03029_;
wire _03030_;
wire _03031_;
wire _03032_;
wire _03033_;
wire _03034_;
wire _03035_;
wire _03036_;
wire _03037_;
wire _03038_;
wire _03039_;
wire _03040_;
wire _03041_;
wire _03042_;
wire _03043_;
wire _03044_;
wire _03045_;
wire _03046_;
wire _03047_;
wire _03048_;
wire _03049_;
wire _03050_;
wire _03051_;
wire _03052_;
wire _03053_;
wire _03054_;
wire _03055_;
wire _03056_;
wire _03057_;
wire _03058_;
wire _03059_;
wire _03060_;
wire _03061_;
wire _03062_;
wire _03063_;
wire _03064_;
wire _03065_;
wire _03066_;
wire _03067_;
wire _03068_;
wire _03069_;
wire _03070_;
wire _03071_;
wire _03072_;
wire _03073_;
wire _03074_;
wire _03075_;
wire _03076_;
wire _03077_;
wire _03078_;
wire _03079_;
wire _03080_;
wire _03081_;
wire _03082_;
wire _03083_;
wire _03084_;
wire _03085_;
wire _03086_;
wire _03087_;
wire _03088_;
wire _03089_;
wire _03090_;
wire _03091_;
wire _03092_;
wire _03093_;
wire _03094_;
wire _03095_;
wire _03096_;
wire _03097_;
wire _03098_;
wire _03099_;
wire _03100_;
wire _03101_;
wire _03102_;
wire _03103_;
wire _03104_;
wire _03105_;
wire _03106_;
wire _03107_;
wire _03108_;
wire _03109_;
wire _03110_;
wire _03111_;
wire _03112_;
wire _03113_;
wire _03114_;
wire _03115_;
wire _03116_;
wire _03117_;
wire _03118_;
wire _03119_;
wire _03120_;
wire _03121_;
wire _03122_;
wire _03123_;
wire _03124_;
wire _03125_;
wire _03126_;
wire _03127_;
wire _03128_;
wire _03129_;
wire _03130_;
wire _03131_;
wire _03132_;
wire _03133_;
wire _03134_;
wire _03135_;
wire _03136_;
wire _03137_;
wire _03138_;
wire _03139_;
wire _03140_;
wire _03141_;
wire _03142_;
wire _03143_;
wire _03144_;
wire _03145_;
wire _03146_;
wire _03147_;
wire _03148_;
wire _03149_;
wire _03150_;
wire _03151_;
wire _03152_;
wire _03153_;
wire _03154_;
wire _03155_;
wire _03156_;
wire _03157_;
wire _03158_;
wire _03159_;
wire _03160_;
wire _03161_;
wire _03162_;
wire _03163_;
wire _03164_;
wire _03165_;
wire _03166_;
wire _03167_;
wire _03168_;
wire _03169_;
wire _03170_;
wire _03171_;
wire _03172_;
wire _03173_;
wire _03174_;
wire _03175_;
wire _03176_;
wire _03177_;
wire _03178_;
wire _03179_;
wire _03180_;
wire _03181_;
wire _03182_;
wire _03183_;
wire _03184_;
wire _03185_;
wire _03186_;
wire _03187_;
wire _03188_;
wire _03189_;
wire _03190_;
wire _03191_;
wire _03192_;
wire _03193_;
wire _03194_;
wire _03195_;
wire _03196_;
wire _03197_;
wire _03198_;
wire _03199_;
wire _03200_;
wire _03201_;
wire _03202_;
wire _03203_;
wire _03204_;
wire _03205_;
wire _03206_;
wire _03207_;
wire _03208_;
wire _03209_;
wire _03210_;
wire _03211_;
wire _03212_;
wire _03213_;
wire _03214_;
wire _03215_;
wire _03216_;
wire _03217_;
wire _03218_;
wire _03219_;
wire _03220_;
wire _03221_;
wire _03222_;
wire _03223_;
wire _03224_;
wire _03225_;
wire _03226_;
wire _03227_;
wire _03228_;
wire _03229_;
wire _03230_;
wire _03231_;
wire _03232_;
wire _03233_;
wire _03234_;
wire _03235_;
wire _03236_;
wire _03237_;
wire _03238_;
wire _03239_;
wire _03240_;
wire _03241_;
wire _03242_;
wire _03243_;
wire _03244_;
wire _03245_;
wire _03246_;
wire _03247_;
wire _03248_;
wire _03249_;
wire _03250_;
wire _03251_;
wire _03252_;
wire _03253_;
wire _03254_;
wire _03255_;
wire _03256_;
wire _03257_;
wire _03258_;
wire _03259_;
wire _03260_;
wire _03261_;
wire _03262_;
wire _03263_;
wire _03264_;
wire _03265_;
wire _03266_;
wire _03267_;
wire _03268_;
wire _03269_;
wire _03270_;
wire _03271_;
wire _03272_;
wire _03273_;
wire _03274_;
wire _03275_;
wire _03276_;
wire _03277_;
wire _03278_;
wire _03279_;
wire _03280_;
wire _03281_;
wire _03282_;
wire _03283_;
wire _03284_;
wire _03285_;
wire _03286_;
wire _03287_;
wire _03288_;
wire _03289_;
wire _03290_;
wire _03291_;
wire _03292_;
wire _03293_;
wire _03294_;
wire _03295_;
wire _03296_;
wire _03297_;
wire _03298_;
wire _03299_;
wire _03300_;
wire _03301_;
wire _03302_;
wire _03303_;
wire _03304_;
wire _03305_;
wire _03306_;
wire _03307_;
wire _03308_;
wire _03309_;
wire _03310_;
wire _03311_;
wire _03312_;
wire _03313_;
wire _03314_;
wire _03315_;
wire _03316_;
wire _03317_;
wire _03318_;
wire _03319_;
wire _03320_;
wire _03321_;
wire _03322_;
wire _03323_;
wire _03324_;
wire _03325_;
wire _03326_;
wire _03327_;
wire _03328_;
wire _03329_;
wire _03330_;
wire _03331_;
wire _03332_;
wire _03333_;
wire _03334_;
wire _03335_;
wire _03336_;
wire _03337_;
wire _03338_;
wire _03339_;
wire _03340_;
wire _03341_;
wire _03342_;
wire _03343_;
wire _03344_;
wire _03345_;
wire _03346_;
wire _03347_;
wire _03348_;
wire _03349_;
wire _03350_;
wire _03351_;
wire _03352_;
wire _03353_;
wire _03354_;
wire _03355_;
wire _03356_;
wire _03357_;
wire _03358_;
wire _03359_;
wire _03360_;
wire _03361_;
wire _03362_;
wire _03363_;
wire _03364_;
wire _03365_;
wire _03366_;
wire _03367_;
wire _03368_;
wire _03369_;
wire _03370_;
wire _03371_;
wire _03372_;
wire _03373_;
wire _03374_;
wire _03375_;
wire _03376_;
wire _03377_;
wire _03378_;
wire _03379_;
wire _03380_;
wire _03381_;
wire _03382_;
wire _03383_;
wire _03384_;
wire _03385_;
wire _03386_;
wire _03387_;
wire _03388_;
wire _03389_;
wire _03390_;
wire _03391_;
wire _03392_;
wire _03393_;
wire _03394_;
wire _03395_;
wire _03396_;
wire _03397_;
wire _03398_;
wire _03399_;
wire _03400_;
wire _03401_;
wire _03402_;
wire _03403_;
wire _03404_;
wire _03405_;
wire _03406_;
wire _03407_;
wire _03408_;
wire _03409_;
wire _03410_;
wire _03411_;
wire _03412_;
wire _03413_;
wire _03414_;
wire _03415_;
wire _03416_;
wire _03417_;
wire _03418_;
wire _03419_;
wire _03420_;
wire _03421_;
wire _03422_;
wire _03423_;
wire _03424_;
wire _03425_;
wire _03426_;
wire _03427_;
wire _03428_;
wire _03429_;
wire _03430_;
wire _03431_;
wire _03432_;
wire _03433_;
wire _03434_;
wire _03435_;
wire _03436_;
wire _03437_;
wire _03438_;
wire _03439_;
wire _03440_;
wire _03441_;
wire _03442_;
wire _03443_;
wire _03444_;
wire _03445_;
wire _03446_;
wire _03447_;
wire _03448_;
wire _03449_;
wire _03450_;
wire _03451_;
wire _03452_;
wire _03453_;
wire _03454_;
wire _03455_;
wire _03456_;
wire _03457_;
wire _03458_;
wire _03459_;
wire _03460_;
wire _03461_;
wire _03462_;
wire _03463_;
wire _03464_;
wire _03465_;
wire _03466_;
wire _03467_;
wire _03468_;
wire _03469_;
wire _03470_;
wire _03471_;
wire _03472_;
wire _03473_;
wire _03474_;
wire _03475_;
wire _03476_;
wire _03477_;
wire _03478_;
wire _03479_;
wire _03480_;
wire _03481_;
wire _03482_;
wire _03483_;
wire _03484_;
wire _03485_;
wire _03486_;
wire _03487_;
wire _03488_;
wire _03489_;
wire _03490_;
wire _03491_;
wire _03492_;
wire _03493_;
wire _03494_;
wire _03495_;
wire _03496_;
wire _03497_;
wire _03498_;
wire _03499_;
wire _03500_;
wire _03501_;
wire _03502_;
wire _03503_;
wire _03504_;
wire _03505_;
wire _03506_;
wire _03507_;
wire _03508_;
wire _03509_;
wire _03510_;
wire _03511_;
wire _03512_;
wire _03513_;
wire _03514_;
wire _03515_;
wire _03516_;
wire _03517_;
wire _03518_;
wire _03519_;
wire _03520_;
wire _03521_;
wire _03522_;
wire _03523_;
wire _03524_;
wire _03525_;
wire _03526_;
wire _03527_;
wire _03528_;
wire _03529_;
wire _03530_;
wire _03531_;
wire _03532_;
wire _03533_;
wire _03534_;
wire _03535_;
wire _03536_;
wire _03537_;
wire _03538_;
wire _03539_;
wire _03540_;
wire _03541_;
wire _03542_;
wire _03543_;
wire _03544_;
wire _03545_;
wire _03546_;
wire _03547_;
wire _03548_;
wire _03549_;
wire _03550_;
wire _03551_;
wire _03552_;
wire _03553_;
wire _03554_;
wire _03555_;
wire _03556_;
wire _03557_;
wire _03558_;
wire _03559_;
wire _03560_;
wire _03561_;
wire _03562_;
wire _03563_;
wire _03564_;
wire _03565_;
wire _03566_;
wire _03567_;
wire _03568_;
wire _03569_;
wire _03570_;
wire _03571_;
wire _03572_;
wire _03573_;
wire _03574_;
wire _03575_;
wire _03576_;
wire _03577_;
wire _03578_;
wire _03579_;
wire _03580_;
wire _03581_;
wire _03582_;
wire _03583_;
wire _03584_;
wire _03585_;
wire _03586_;
wire _03587_;
wire _03588_;
wire _03589_;
wire _03590_;
wire _03591_;
wire _03592_;
wire _03593_;
wire _03594_;
wire _03595_;
wire _03596_;
wire _03597_;
wire _03598_;
wire _03599_;
wire _03600_;
wire _03601_;
wire _03602_;
wire _03603_;
wire _03604_;
wire _03605_;
wire _03606_;
wire _03607_;
wire _03608_;
wire _03609_;
wire _03610_;
wire _03611_;
wire _03612_;
wire _03613_;
wire _03614_;
wire _03615_;
wire _03616_;
wire _03617_;
wire _03618_;
wire _03619_;
wire _03620_;
wire _03621_;
wire _03622_;
wire _03623_;
wire _03624_;
wire _03625_;
wire _03626_;
wire _03627_;
wire _03628_;
wire _03629_;
wire _03630_;
wire _03631_;
wire _03632_;
wire _03633_;
wire _03634_;
wire _03635_;
wire _03636_;
wire _03637_;
wire _03638_;
wire _03639_;
wire _03640_;
wire _03641_;
wire _03642_;
wire _03643_;
wire _03644_;
wire _03645_;
wire _03646_;
wire _03647_;
wire _03648_;
wire _03649_;
wire _03650_;
wire _03651_;
wire _03652_;
wire _03653_;
wire _03654_;
wire _03655_;
wire _03656_;
wire _03657_;
wire _03658_;
wire _03659_;
wire _03660_;
wire _03661_;
wire _03662_;
wire _03663_;
wire _03664_;
wire _03665_;
wire _03666_;
wire _03667_;
wire _03668_;
wire _03669_;
wire _03670_;
wire _03671_;
wire _03672_;
wire _03673_;
wire _03674_;
wire _03675_;
wire _03676_;
wire _03677_;
wire _03678_;
wire _03679_;
wire _03680_;
wire _03681_;
wire _03682_;
wire _03683_;
wire _03684_;
wire _03685_;
wire _03686_;
wire _03687_;
wire _03688_;
wire _03689_;
wire _03690_;
wire _03691_;
wire _03692_;
wire _03693_;
wire _03694_;
wire _03695_;
wire _03696_;
wire _03697_;
wire _03698_;
wire _03699_;
wire _03700_;
wire _03701_;
wire _03702_;
wire _03703_;
wire _03704_;
wire _03705_;
wire _03706_;
wire _03707_;
wire _03708_;
wire _03709_;
wire _03710_;
wire _03711_;
wire _03712_;
wire _03713_;
wire _03714_;
wire _03715_;
wire _03716_;
wire _03717_;
wire _03718_;
wire _03719_;
wire _03720_;
wire _03721_;
wire _03722_;
wire _03723_;
wire _03724_;
wire _03725_;
wire _03726_;
wire _03727_;
wire _03728_;
wire _03729_;
wire _03730_;
wire _03731_;
wire _03732_;
wire _03733_;
wire _03734_;
wire _03735_;
wire _03736_;
wire _03737_;
wire _03738_;
wire _03739_;
wire _03740_;
wire _03741_;
wire _03742_;
wire _03743_;
wire _03744_;
wire _03745_;
wire _03746_;
wire _03747_;
wire _03748_;
wire _03749_;
wire _03750_;
wire _03751_;
wire _03752_;
wire _03753_;
wire _03754_;
wire _03755_;
wire _03756_;
wire _03757_;
wire _03758_;
wire _03759_;
wire _03760_;
wire _03761_;
wire _03762_;
wire _03763_;
wire _03764_;
wire _03765_;
wire _03766_;
wire _03767_;
wire _03768_;
wire _03769_;
wire _03770_;
wire _03771_;
wire _03772_;
wire _03773_;
wire _03774_;
wire _03775_;
wire _03776_;
wire _03777_;
wire _03778_;
wire _03779_;
wire _03780_;
wire _03781_;
wire _03782_;
wire _03783_;
wire _03784_;
wire _03785_;
wire _03786_;
wire _03787_;
wire _03788_;
wire _03789_;
wire _03790_;
wire _03791_;
wire _03792_;
wire _03793_;
wire _03794_;
wire _03795_;
wire _03796_;
wire _03797_;
wire _03798_;
wire _03799_;
wire _03800_;
wire _03801_;
wire _03802_;
wire _03803_;
wire _03804_;
wire _03805_;
wire _03806_;
wire _03807_;
wire _03808_;
wire _03809_;
wire _03810_;
wire _03811_;
wire _03812_;
wire _03813_;
wire _03814_;
wire _03815_;
wire _03816_;
wire _03817_;
wire _03818_;
wire _03819_;
wire _03820_;
wire _03821_;
wire _03822_;
wire _03823_;
wire _03824_;
wire _03825_;
wire _03826_;
wire _03827_;
wire _03828_;
wire _03829_;
wire _03830_;
wire _03831_;
wire _03832_;
wire _03833_;
wire _03834_;
wire _03835_;
wire _03836_;
wire _03837_;
wire _03838_;
wire _03839_;
wire _03840_;
wire _03841_;
wire _03842_;
wire _03843_;
wire _03844_;
wire _03845_;
wire _03846_;
wire _03847_;
wire _03848_;
wire _03849_;
wire _03850_;
wire _03851_;
wire _03852_;
wire _03853_;
wire _03854_;
wire _03855_;
wire _03856_;
wire _03857_;
wire _03858_;
wire _03859_;
wire _03860_;
wire _03861_;
wire _03862_;
wire _03863_;
wire _03864_;
wire _03865_;
wire _03866_;
wire _03867_;
wire _03868_;
wire _03869_;
wire _03870_;
wire _03871_;
wire _03872_;
wire _03873_;
wire _03874_;
wire _03875_;
wire _03876_;
wire _03877_;
wire _03878_;
wire _03879_;
wire _03880_;
wire _03881_;
wire _03882_;
wire _03883_;
wire _03884_;
wire _03885_;
wire _03886_;
wire _03887_;
wire _03888_;
wire _03889_;
wire _03890_;
wire _03891_;
wire _03892_;
wire _03893_;
wire _03894_;
wire _03895_;
wire _03896_;
wire _03897_;
wire _03898_;
wire _03899_;
wire _03900_;
wire _03901_;
wire _03902_;
wire _03903_;
wire _03904_;
wire _03905_;
wire _03906_;
wire _03907_;
wire _03908_;
wire _03909_;
wire _03910_;
wire _03911_;
wire _03912_;
wire _03913_;
wire _03914_;
wire _03915_;
wire _03916_;
wire _03917_;
wire _03918_;
wire _03919_;
wire _03920_;
wire _03921_;
wire _03922_;
wire _03923_;
wire _03924_;
wire _03925_;
wire _03926_;
wire _03927_;
wire _03928_;
wire _03929_;
wire _03930_;
wire _03931_;
wire _03932_;
wire _03933_;
wire _03934_;
wire _03935_;
wire _03936_;
wire _03937_;
wire _03938_;
wire _03939_;
wire _03940_;
wire _03941_;
wire _03942_;
wire _03943_;
wire _03944_;
wire _03945_;
wire _03946_;
wire _03947_;
wire _03948_;
wire _03949_;
wire _03950_;
wire _03951_;
wire _03952_;
wire _03953_;
wire _03954_;
wire _03955_;
wire _03956_;
wire _03957_;
wire _03958_;
wire _03959_;
wire _03960_;
wire _03961_;
wire _03962_;
wire _03963_;
wire _03964_;
wire _03965_;
wire _03966_;
wire _03967_;
wire _03968_;
wire _03969_;
wire _03970_;
wire _03971_;
wire _03972_;
wire _03973_;
wire _03974_;
wire _03975_;
wire _03976_;
wire _03977_;
wire _03978_;
wire _03979_;
wire _03980_;
wire _03981_;
wire _03982_;
wire _03983_;
wire _03984_;
wire _03985_;
wire _03986_;
wire _03987_;
wire _03988_;
wire _03989_;
wire _03990_;
wire _03991_;
wire _03992_;
wire _03993_;
wire _03994_;
wire _03995_;
wire _03996_;
wire _03997_;
wire _03998_;
wire _03999_;
wire _04000_;
wire _04001_;
wire _04002_;
wire _04003_;
wire _04004_;
wire _04005_;
wire _04006_;
wire _04007_;
wire _04008_;
wire _04009_;
wire _04010_;
wire _04011_;
wire _04012_;
wire _04013_;
wire _04014_;
wire _04015_;
wire _04016_;
wire _04017_;
wire _04018_;
wire _04019_;
wire _04020_;
wire _04021_;
wire _04022_;
wire _04023_;
wire _04024_;
wire _04025_;
wire _04026_;
wire _04027_;
wire _04028_;
wire _04029_;
wire _04030_;
wire _04031_;
wire _04032_;
wire _04033_;
wire _04034_;
wire _04035_;
wire _04036_;
wire _04037_;
wire _04038_;
wire _04039_;
wire _04040_;
wire _04041_;
wire _04042_;
wire _04043_;
wire _04044_;
wire _04045_;
wire _04046_;
wire _04047_;
wire _04048_;
wire _04049_;
wire _04050_;
wire _04051_;
wire _04052_;
wire _04053_;
wire _04054_;
wire _04055_;
wire _04056_;
wire _04057_;
wire _04058_;
wire _04059_;
wire _04060_;
wire _04061_;
wire _04062_;
wire _04063_;
wire _04064_;
wire _04065_;
wire _04066_;
wire _04067_;
wire _04068_;
wire _04069_;
wire _04070_;
wire _04071_;
wire _04072_;
wire _04073_;
wire _04074_;
wire _04075_;
wire _04076_;
wire _04077_;
wire _04078_;
wire _04079_;
wire _04080_;
wire _04081_;
wire _04082_;
wire _04083_;
wire _04084_;
wire _04085_;
wire _04086_;
wire _04087_;
wire _04088_;
wire _04089_;
wire _04090_;
wire _04091_;
wire _04092_;
wire _04093_;
wire _04094_;
wire _04095_;
wire _04096_;
wire _04097_;
wire _04098_;
wire _04099_;
wire _04100_;
wire _04101_;
wire _04102_;
wire _04103_;
wire _04104_;
wire _04105_;
wire _04106_;
wire _04107_;
wire _04108_;
wire _04109_;
wire _04110_;
wire _04111_;
wire _04112_;
wire _04113_;
wire _04114_;
wire _04115_;
wire _04116_;
wire _04117_;
wire _04118_;
wire _04119_;
wire _04120_;
wire _04121_;
wire _04122_;
wire _04123_;
wire _04124_;
wire _04125_;
wire _04126_;
wire _04127_;
wire _04128_;
wire _04129_;
wire _04130_;
wire _04131_;
wire _04132_;
wire _04133_;
wire _04134_;
wire _04135_;
wire _04136_;
wire _04137_;
wire _04138_;
wire _04139_;
wire _04140_;
wire _04141_;
wire _04142_;
wire _04143_;
wire _04144_;
wire _04145_;
wire _04146_;
wire _04147_;
wire _04148_;
wire _04149_;
wire _04150_;
wire _04151_;
wire _04152_;
wire _04153_;
wire _04154_;
wire _04155_;
wire _04156_;
wire _04157_;
wire _04158_;
wire _04159_;
wire _04160_;
wire _04161_;
wire _04162_;
wire _04163_;
wire _04164_;
wire _04165_;
wire _04166_;
wire _04167_;
wire _04168_;
wire _04169_;
wire _04170_;
wire _04171_;
wire _04172_;
wire _04173_;
wire _04174_;
wire _04175_;
wire _04176_;
wire _04177_;
wire _04178_;
wire _04179_;
wire _04180_;
wire _04181_;
wire _04182_;
wire _04183_;
wire _04184_;
wire _04185_;
wire _04186_;
wire _04187_;
wire _04188_;
wire _04189_;
wire _04190_;
wire _04191_;
wire _04192_;
wire _04193_;
wire _04194_;
wire _04195_;
wire _04196_;
wire _04197_;
wire _04198_;
wire _04199_;
wire _04200_;
wire _04201_;
wire _04202_;
wire _04203_;
wire _04204_;
wire _04205_;
wire _04206_;
wire _04207_;
wire _04208_;
wire _04209_;
wire _04210_;
wire _04211_;
wire _04212_;
wire _04213_;
wire _04214_;
wire _04215_;
wire _04216_;
wire _04217_;
wire _04218_;
wire _04219_;
wire _04220_;
wire _04221_;
wire _04222_;
wire _04223_;
wire _04224_;
wire _04225_;
wire _04226_;
wire _04227_;
wire _04228_;
wire _04229_;
wire _04230_;
wire _04231_;
wire _04232_;
wire _04233_;
wire _04234_;
wire _04235_;
wire _04236_;
wire _04237_;
wire _04238_;
wire _04239_;
wire _04240_;
wire _04241_;
wire _04242_;
wire _04243_;
wire _04244_;
wire _04245_;
wire _04246_;
wire _04247_;
wire _04248_;
wire _04249_;
wire _04250_;
wire _04251_;
wire _04252_;
wire _04253_;
wire _04254_;
wire _04255_;
wire _04256_;
wire _04257_;
wire _04258_;
wire _04259_;
wire _04260_;
wire _04261_;
wire _04262_;
wire _04263_;
wire _04264_;
wire _04265_;
wire _04266_;
wire _04267_;
wire _04268_;
wire _04269_;
wire _04270_;
wire _04271_;
wire _04272_;
wire _04273_;
wire _04274_;
wire _04275_;
wire _04276_;
wire _04277_;
wire _04278_;
wire _04279_;
wire _04280_;
wire _04281_;
wire _04282_;
wire _04283_;
wire _04284_;
wire _04285_;
wire _04286_;
wire _04287_;
wire _04288_;
wire _04289_;
wire _04290_;
wire _04291_;
wire _04292_;
wire _04293_;
wire _04294_;
wire _04295_;
wire _04296_;
wire _04297_;
wire _04298_;
wire _04299_;
wire _04300_;
wire _04301_;
wire _04302_;
wire _04303_;
wire _04304_;
wire _04305_;
wire _04306_;
wire _04307_;
wire _04308_;
wire _04309_;
wire _04310_;
wire _04311_;
wire _04312_;
wire _04313_;
wire _04314_;
wire _04315_;
wire _04316_;
wire _04317_;
wire _04318_;
wire _04319_;
wire _04320_;
wire _04321_;
wire _04322_;
wire _04323_;
wire _04324_;
wire _04325_;
wire _04326_;
wire _04327_;
wire _04328_;
wire _04329_;
wire _04330_;
wire _04331_;
wire _04332_;
wire _04333_;
wire _04334_;
wire _04335_;
wire _04336_;
wire _04337_;
wire _04338_;
wire _04339_;
wire _04340_;
wire _04341_;
wire _04342_;
wire _04343_;
wire _04344_;
wire _04345_;
wire _04346_;
wire _04347_;
wire _04348_;
wire _04349_;
wire _04350_;
wire _04351_;
wire _04352_;
wire _04353_;
wire _04354_;
wire _04355_;
wire _04356_;
wire _04357_;
wire _04358_;
wire _04359_;
wire _04360_;
wire _04361_;
wire _04362_;
wire _04363_;
wire _04364_;
wire _04365_;
wire _04366_;
wire _04367_;
wire _04368_;
wire _04369_;
wire _04370_;
wire _04371_;
wire _04372_;
wire _04373_;
wire _04374_;
wire _04375_;
wire _04376_;
wire _04377_;
wire _04378_;
wire _04379_;
wire _04380_;
wire _04381_;
wire _04382_;
wire _04383_;
wire _04384_;
wire _04385_;
wire _04386_;
wire _04387_;
wire _04388_;
wire _04389_;
wire _04390_;
wire _04391_;
wire _04392_;
wire _04393_;
wire _04394_;
wire _04395_;
wire _04396_;
wire _04397_;
wire _04398_;
wire _04399_;
wire _04400_;
wire _04401_;
wire _04402_;
wire _04403_;
wire _04404_;
wire _04405_;
wire _04406_;
wire _04407_;
wire _04408_;
wire _04409_;
wire _04410_;
wire _04411_;
wire _04412_;
wire _04413_;
wire _04414_;
wire _04415_;
wire _04416_;
wire _04417_;
wire _04418_;
wire _04419_;
wire _04420_;
wire _04421_;
wire _04422_;
wire _04423_;
wire _04424_;
wire _04425_;
wire _04426_;
wire _04427_;
wire _04428_;
wire _04429_;
wire _04430_;
wire _04431_;
wire _04432_;
wire _04433_;
wire _04434_;
wire _04435_;
wire _04436_;
wire _04437_;
wire _04438_;
wire _04439_;
wire _04440_;
wire _04441_;
wire _04442_;
wire _04443_;
wire _04444_;
wire _04445_;
wire _04446_;
wire _04447_;
wire _04448_;
wire _04449_;
wire _04450_;
wire _04451_;
wire _04452_;
wire _04453_;
wire _04454_;
wire _04455_;
wire _04456_;
wire _04457_;
wire _04458_;
wire _04459_;
wire _04460_;
wire _04461_;
wire _04462_;
wire _04463_;
wire _04464_;
wire _04465_;
wire _04466_;
wire _04467_;
wire _04468_;
wire _04469_;
wire _04470_;
wire _04471_;
wire _04472_;
wire _04473_;
wire _04474_;
wire _04475_;
wire _04476_;
wire _04477_;
wire _04478_;
wire _04479_;
wire _04480_;
wire _04481_;
wire _04482_;
wire _04483_;
wire _04484_;
wire _04485_;
wire _04486_;
wire _04487_;
wire _04488_;
wire _04489_;
wire _04490_;
wire _04491_;
wire _04492_;
wire _04493_;
wire _04494_;
wire _04495_;
wire _04496_;
wire _04497_;
wire _04498_;
wire _04499_;
wire _04500_;
wire _04501_;
wire _04502_;
wire _04503_;
wire _04504_;
wire _04505_;
wire _04506_;
wire _04507_;
wire _04508_;
wire _04509_;
wire _04510_;
wire _04511_;
wire _04512_;
wire _04513_;
wire _04514_;
wire _04515_;
wire _04516_;
wire _04517_;
wire _04518_;
wire _04519_;
wire _04520_;
wire _04521_;
wire _04522_;
wire _04523_;
wire _04524_;
wire _04525_;
wire _04526_;
wire _04527_;
wire _04528_;
wire _04529_;
wire _04530_;
wire _04531_;
wire _04532_;
wire _04533_;
wire _04534_;
wire _04535_;
wire _04536_;
wire _04537_;
wire _04538_;
wire _04539_;
wire _04540_;
wire _04541_;
wire _04542_;
wire _04543_;
wire _04544_;
wire _04545_;
wire _04546_;
wire _04547_;
wire _04548_;
wire _04549_;
wire _04550_;
wire _04551_;
wire _04552_;
wire _04553_;
wire _04554_;
wire _04555_;
wire _04556_;
wire _04557_;
wire _04558_;
wire _04559_;
wire _04560_;
wire _04561_;
wire _04562_;
wire _04563_;
wire _04564_;
wire _04565_;
wire _04566_;
wire _04567_;
wire _04568_;
wire _04569_;
wire _04570_;
wire _04571_;
wire _04572_;
wire _04573_;
wire _04574_;
wire _04575_;
wire _04576_;
wire _04577_;
wire _04578_;
wire _04579_;
wire _04580_;
wire _04581_;
wire _04582_;
wire _04583_;
wire _04584_;
wire _04585_;
wire _04586_;
wire _04587_;
wire _04588_;
wire _04589_;
wire _04590_;
wire _04591_;
wire _04592_;
wire _04593_;
wire _04594_;
wire _04595_;
wire _04596_;
wire _04597_;
wire _04598_;
wire _04599_;
wire _04600_;
wire _04601_;
wire _04602_;
wire _04603_;
wire _04604_;
wire _04605_;
wire _04606_;
wire _04607_;
wire _04608_;
wire _04609_;
wire _04610_;
wire _04611_;
wire _04612_;
wire _04613_;
wire _04614_;
wire _04615_;
wire _04616_;
wire _04617_;
wire _04618_;
wire _04619_;
wire _04620_;
wire _04621_;
wire _04622_;
wire _04623_;
wire _04624_;
wire _04625_;
wire _04626_;
wire _04627_;
wire _04628_;
wire _04629_;
wire _04630_;
wire _04631_;
wire _04632_;
wire _04633_;
wire _04634_;
wire _04635_;
wire _04636_;
wire _04637_;
wire _04638_;
wire _04639_;
wire _04640_;
wire _04641_;
wire _04642_;
wire _04643_;
wire _04644_;
wire _04645_;
wire _04646_;
wire _04647_;
wire _04648_;
wire _04649_;
wire _04650_;
wire _04651_;
wire _04652_;
wire _04653_;
wire _04654_;
wire _04655_;
wire _04656_;
wire _04657_;
wire _04658_;
wire _04659_;
wire _04660_;
wire _04661_;
wire _04662_;
wire _04663_;
wire _04664_;
wire _04665_;
wire _04666_;
wire _04667_;
wire _04668_;
wire _04669_;
wire _04670_;
wire _04671_;
wire _04672_;
wire _04673_;
wire _04674_;
wire _04675_;
wire _04676_;
wire _04677_;
wire _04678_;
wire _04679_;
wire _04680_;
wire _04681_;
wire _04682_;
wire _04683_;
wire _04684_;
wire _04685_;
wire _04686_;
wire _04687_;
wire _04688_;
wire _04689_;
wire _04690_;
wire _04691_;
wire _04692_;
wire _04693_;
wire _04694_;
wire _04695_;
wire _04696_;
wire _04697_;
wire _04698_;
wire _04699_;
wire _04700_;
wire _04701_;
wire _04702_;
wire _04703_;
wire _04704_;
wire _04705_;
wire _04706_;
wire _04707_;
wire _04708_;
wire _04709_;
wire _04710_;
wire _04711_;
wire _04712_;
wire _04713_;
wire _04714_;
wire _04715_;
wire _04716_;
wire _04717_;
wire _04718_;
wire _04719_;
wire _04720_;
wire _04721_;
wire _04722_;
wire _04723_;
wire _04724_;
wire _04725_;
wire _04726_;
wire _04727_;
wire _04728_;
wire _04729_;
wire _04730_;
wire _04731_;
wire _04732_;
wire _04733_;
wire _04734_;
wire _04735_;
wire _04736_;
wire _04737_;
wire _04738_;
wire _04739_;
wire _04740_;
wire _04741_;
wire _04742_;
wire _04743_;
wire _04744_;
wire _04745_;
wire _04746_;
wire _04747_;
wire _04748_;
wire _04749_;
wire _04750_;
wire _04751_;
wire _04752_;
wire _04753_;
wire _04754_;
wire _04755_;
wire _04756_;
wire _04757_;
wire _04758_;
wire _04759_;
wire _04760_;
wire _04761_;
wire _04762_;
wire _04763_;
wire _04764_;
wire _04765_;
wire _04766_;
wire _04767_;
wire _04768_;
wire _04769_;
wire _04770_;
wire _04771_;
wire _04772_;
wire _04773_;
wire _04774_;
wire _04775_;
wire _04776_;
wire _04777_;
wire _04778_;
wire _04779_;
wire _04780_;
wire _04781_;
wire _04782_;
wire _04783_;
wire _04784_;
wire _04785_;
wire _04786_;
wire _04787_;
wire _04788_;
wire _04789_;
wire _04790_;
wire _04791_;
wire _04792_;
wire _04793_;
wire _04794_;
wire _04795_;
wire _04796_;
wire _04797_;
wire _04798_;
wire _04799_;
wire _04800_;
wire _04801_;
wire _04802_;
wire _04803_;
wire _04804_;
wire _04805_;
wire _04806_;
wire _04807_;
wire _04808_;
wire _04809_;
wire _04810_;
wire _04811_;
wire _04812_;
wire _04813_;
wire _04814_;
wire _04815_;
wire _04816_;
wire _04817_;
wire _04818_;
wire _04819_;
wire _04820_;
wire _04821_;
wire _04822_;
wire _04823_;
wire _04824_;
wire _04825_;
wire _04826_;
wire _04827_;
wire _04828_;
wire _04829_;
wire _04830_;
wire _04831_;
wire _04832_;
wire _04833_;
wire _04834_;
wire _04835_;
wire _04836_;
wire _04837_;
wire _04838_;
wire _04839_;
wire _04840_;
wire _04841_;
wire _04842_;
wire _04843_;
wire _04844_;
wire _04845_;
wire _04846_;
wire _04847_;
wire _04848_;
wire _04849_;
wire _04850_;
wire _04851_;
wire _04852_;
wire _04853_;
wire _04854_;
wire _04855_;
wire _04856_;
wire _04857_;
wire _04858_;
wire _04859_;
wire _04860_;
wire _04861_;
wire _04862_;
wire _04863_;
wire _04864_;
wire _04865_;
wire _04866_;
wire _04867_;
wire _04868_;
wire _04869_;
wire _04870_;
wire _04871_;
wire _04872_;
wire _04873_;
wire _04874_;
wire _04875_;
wire _04876_;
wire _04877_;
wire _04878_;
wire _04879_;
wire _04880_;
wire _04881_;
wire _04882_;
wire _04883_;
wire _04884_;
wire _04885_;
wire _04886_;
wire _04887_;
wire _04888_;
wire _04889_;
wire _04890_;
wire _04891_;
wire _04892_;
wire _04893_;
wire _04894_;
wire _04895_;
wire _04896_;
wire _04897_;
wire _04898_;
wire _04899_;
wire _04900_;
wire _04901_;
wire _04902_;
wire _04903_;
wire _04904_;
wire _04905_;
wire _04906_;
wire _04907_;
wire _04908_;
wire _04909_;
wire _04910_;
wire _04911_;
wire _04912_;
wire _04913_;
wire _04914_;
wire _04915_;
wire _04916_;
wire _04917_;
wire _04918_;
wire _04919_;
wire _04920_;
wire _04921_;
wire _04922_;
wire _04923_;
wire _04924_;
wire _04925_;
wire _04926_;
wire _04927_;
wire _04928_;
wire _04929_;
wire _04930_;
wire _04931_;
wire _04932_;
wire _04933_;
wire _04934_;
wire _04935_;
wire _04936_;
wire _04937_;
wire _04938_;
wire _04939_;
wire _04940_;
wire _04941_;
wire _04942_;
wire _04943_;
wire _04944_;
wire _04945_;
wire _04946_;
wire _04947_;
wire _04948_;
wire _04949_;
wire _04950_;
wire _04951_;
wire _04952_;
wire _04953_;
wire _04954_;
wire _04955_;
wire _04956_;
wire _04957_;
wire _04958_;
wire _04959_;
wire _04960_;
wire _04961_;
wire _04962_;
wire _04963_;
wire _04964_;
wire _04965_;
wire _04966_;
wire _04967_;
wire _04968_;
wire _04969_;
wire _04970_;
wire _04971_;
wire _04972_;
wire _04973_;
wire _04974_;
wire _04975_;
wire _04976_;
wire _04977_;
wire _04978_;
wire _04979_;
wire _04980_;
wire _04981_;
wire _04982_;
wire _04983_;
wire _04984_;
wire _04985_;
wire _04986_;
wire _04987_;
wire _04988_;
wire _04989_;
wire _04990_;
wire _04991_;
wire _04992_;
wire _04993_;
wire _04994_;
wire _04995_;
wire _04996_;
wire _04997_;
wire _04998_;
wire _04999_;
wire _05000_;
wire _05001_;
wire _05002_;
wire _05003_;
wire _05004_;
wire _05005_;
wire _05006_;
wire _05007_;
wire _05008_;
wire _05009_;
wire _05010_;
wire _05011_;
wire _05012_;
wire _05013_;
wire _05014_;
wire _05015_;
wire _05016_;
wire _05017_;
wire _05018_;
wire _05019_;
wire _05020_;
wire _05021_;
wire _05022_;
wire _05023_;
wire _05024_;
wire _05025_;
wire _05026_;
wire _05027_;
wire _05028_;
wire _05029_;
wire _05030_;
wire _05031_;
wire _05032_;
wire _05033_;
wire _05034_;
wire _05035_;
wire _05036_;
wire _05037_;
wire _05038_;
wire _05039_;
wire _05040_;
wire _05041_;
wire _05042_;
wire _05043_;
wire _05044_;
wire _05045_;
wire _05046_;
wire _05047_;
wire _05048_;
wire _05049_;
wire _05050_;
wire _05051_;
wire _05052_;
wire _05053_;
wire _05054_;
wire _05055_;
wire _05056_;
wire _05057_;
wire _05058_;
wire _05059_;
wire _05060_;
wire _05061_;
wire _05062_;
wire _05063_;
wire _05064_;
wire _05065_;
wire _05066_;
wire _05067_;
wire _05068_;
wire _05069_;
wire _05070_;
wire _05071_;
wire _05072_;
wire _05073_;
wire _05074_;
wire _05075_;
wire _05076_;
wire _05077_;
wire _05078_;
wire _05079_;
wire _05080_;
wire _05081_;
wire _05082_;
wire _05083_;
wire _05084_;
wire _05085_;
wire _05086_;
wire _05087_;
wire _05088_;
wire _05089_;
wire _05090_;
wire _05091_;
wire _05092_;
wire _05093_;
wire _05094_;
wire _05095_;
wire _05096_;
wire _05097_;
wire _05098_;
wire _05099_;
wire _05100_;
wire _05101_;
wire _05102_;
wire _05103_;
wire _05104_;
wire _05105_;
wire _05106_;
wire _05107_;
wire _05108_;
wire _05109_;
wire _05110_;
wire _05111_;
wire _05112_;
wire _05113_;
wire _05114_;
wire _05115_;
wire _05116_;
wire _05117_;
wire _05118_;
wire _05119_;
wire _05120_;
wire _05121_;
wire _05122_;
wire _05123_;
wire _05124_;
wire _05125_;
wire _05126_;
wire _05127_;
wire _05128_;
wire _05129_;
wire _05130_;
wire _05131_;
wire _05132_;
wire _05133_;
wire _05134_;
wire _05135_;
wire _05136_;
wire _05137_;
wire _05138_;
wire _05139_;
wire _05140_;
wire _05141_;
wire _05142_;
wire _05143_;
wire _05144_;
wire _05145_;
wire _05146_;
wire _05147_;
wire _05148_;
wire _05149_;
wire _05150_;
wire _05151_;
wire _05152_;
wire _05153_;
wire _05154_;
wire _05155_;
wire _05156_;
wire _05157_;
wire _05158_;
wire _05159_;
wire _05160_;
wire _05161_;
wire _05162_;
wire _05163_;
wire _05164_;
wire _05165_;
wire _05166_;
wire _05167_;
wire _05168_;
wire _05169_;
wire _05170_;
wire _05171_;
wire _05172_;
wire _05173_;
wire _05174_;
wire _05175_;
wire _05176_;
wire _05177_;
wire _05178_;
wire _05179_;
wire _05180_;
wire _05181_;
wire _05182_;
wire _05183_;
wire _05184_;
wire _05185_;
wire _05186_;
wire _05187_;
wire _05188_;
wire _05189_;
wire _05190_;
wire _05191_;
wire _05192_;
wire _05193_;
wire _05194_;
wire _05195_;
wire _05196_;
wire _05197_;
wire _05198_;
wire _05199_;
wire _05200_;
wire _05201_;
wire _05202_;
wire _05203_;
wire _05204_;
wire _05205_;
wire _05206_;
wire _05207_;
wire _05208_;
wire _05209_;
wire _05210_;
wire _05211_;
wire _05212_;
wire _05213_;
wire _05214_;
wire _05215_;
wire _05216_;
wire _05217_;
wire _05218_;
wire _05219_;
wire _05220_;
wire _05221_;
wire _05222_;
wire _05223_;
wire _05224_;
wire _05225_;
wire _05226_;
wire _05227_;
wire _05228_;
wire _05229_;
wire _05230_;
wire _05231_;
wire _05232_;
wire _05233_;
wire _05234_;
wire _05235_;
wire _05236_;
wire _05237_;
wire _05238_;
wire _05239_;
wire _05240_;
wire _05241_;
wire _05242_;
wire _05243_;
wire _05244_;
wire _05245_;
wire _05246_;
wire _05247_;
wire _05248_;
wire _05249_;
wire _05250_;
wire _05251_;
wire _05252_;
wire _05253_;
wire _05254_;
wire _05255_;
wire _05256_;
wire _05257_;
wire _05258_;
wire _05259_;
wire _05260_;
wire _05261_;
wire _05262_;
wire _05263_;
wire _05264_;
wire _05265_;
wire _05266_;
wire _05267_;
wire _05268_;
wire _05269_;
wire _05270_;
wire _05271_;
wire _05272_;
wire _05273_;
wire _05274_;
wire _05275_;
wire _05276_;
wire _05277_;
wire _05278_;
wire _05279_;
wire _05280_;
wire _05281_;
wire _05282_;
wire _05283_;
wire _05284_;
wire _05285_;
wire _05286_;
wire _05287_;
wire _05288_;
wire _05289_;
wire _05290_;
wire _05291_;
wire _05292_;
wire _05293_;
wire _05294_;
wire _05295_;
wire _05296_;
wire _05297_;
wire _05298_;
wire _05299_;
wire _05300_;
wire _05301_;
wire _05302_;
wire _05303_;
wire _05304_;
wire _05305_;
wire _05306_;
wire _05307_;
wire _05308_;
wire _05309_;
wire _05310_;
wire _05311_;
wire _05312_;
wire _05313_;
wire _05314_;
wire _05315_;
wire _05316_;
wire _05317_;
wire _05318_;
wire _05319_;
wire _05320_;
wire _05321_;
wire _05322_;
wire _05323_;
wire _05324_;
wire _05325_;
wire _05326_;
wire _05327_;
wire _05328_;
wire _05329_;
wire _05330_;
wire _05331_;
wire _05332_;
wire _05333_;
wire _05334_;
wire _05335_;
wire _05336_;
wire _05337_;
wire _05338_;
wire _05339_;
wire _05340_;
wire _05341_;
wire _05342_;
wire _05343_;
wire _05344_;
wire _05345_;
wire _05346_;
wire _05347_;
wire _05348_;
wire _05349_;
wire _05350_;
wire _05351_;
wire _05352_;
wire _05353_;
wire _05354_;
wire _05355_;
wire _05356_;
wire _05357_;
wire _05358_;
wire _05359_;
wire _05360_;
wire _05361_;
wire _05362_;
wire _05363_;
wire _05364_;
wire _05365_;
wire _05366_;
wire _05367_;
wire _05368_;
wire _05369_;
wire _05370_;
wire _05371_;
wire _05372_;
wire _05373_;
wire _05374_;
wire _05375_;
wire _05376_;
wire _05377_;
wire _05378_;
wire _05379_;
wire _05380_;
wire _05381_;
wire _05382_;
wire _05383_;
wire _05384_;
wire _05385_;
wire _05386_;
wire _05387_;
wire _05388_;
wire _05389_;
wire _05390_;
wire _05391_;
wire _05392_;
wire _05393_;
wire _05394_;
wire _05395_;
wire _05396_;
wire _05397_;
wire _05398_;
wire _05399_;
wire _05400_;
wire _05401_;
wire _05402_;
wire _05403_;
wire _05404_;
wire _05405_;
wire _05406_;
wire _05407_;
wire _05408_;
wire _05409_;
wire _05410_;
wire _05411_;
wire _05412_;
wire _05413_;
wire _05414_;
wire _05415_;
wire _05416_;
wire _05417_;
wire _05418_;
wire _05419_;
wire _05420_;
wire _05421_;
wire _05422_;
wire _05423_;
wire _05424_;
wire _05425_;
wire _05426_;
wire _05427_;
wire _05428_;
wire _05429_;
wire _05430_;
wire _05431_;
wire _05432_;
wire _05433_;
wire _05434_;
wire _05435_;
wire _05436_;
wire _05437_;
wire _05438_;
wire _05439_;
wire _05440_;
wire _05441_;
wire _05442_;
wire _05443_;
wire _05444_;
wire _05445_;
wire _05446_;
wire _05447_;
wire _05448_;
wire _05449_;
wire _05450_;
wire _05451_;
wire _05452_;
wire _05453_;
wire _05454_;
wire _05455_;
wire _05456_;
wire _05457_;
wire _05458_;
wire _05459_;
wire _05460_;
wire _05461_;
wire _05462_;
wire _05463_;
wire _05464_;
wire _05465_;
wire _05466_;
wire _05467_;
wire _05468_;
wire _05469_;
wire _05470_;
wire _05471_;
wire _05472_;
wire _05473_;
wire _05474_;
wire _05475_;
wire _05476_;
wire _05477_;
wire _05478_;
wire _05479_;
wire _05480_;
wire _05481_;
wire _05482_;
wire _05483_;
wire _05484_;
wire _05485_;
wire _05486_;
wire _05487_;
wire _05488_;
wire _05489_;
wire _05490_;
wire _05491_;
wire _05492_;
wire _05493_;
wire _05494_;
wire _05495_;
wire _05496_;
wire _05497_;
wire _05498_;
wire _05499_;
wire _05500_;
wire _05501_;
wire _05502_;
wire _05503_;
wire _05504_;
wire _05505_;
wire _05506_;
wire _05507_;
wire _05508_;
wire _05509_;
wire _05510_;
wire _05511_;
wire _05512_;
wire _05513_;
wire _05514_;
wire _05515_;
wire _05516_;
wire _05517_;
wire _05518_;
wire _05519_;
wire _05520_;
wire _05521_;
wire _05522_;
wire _05523_;
wire _05524_;
wire _05525_;
wire _05526_;
wire _05527_;
wire _05528_;
wire _05529_;
wire _05530_;
wire _05531_;
wire _05532_;
wire _05533_;
wire _05534_;
wire _05535_;
wire _05536_;
wire _05537_;
wire _05538_;
wire _05539_;
wire _05540_;
wire _05541_;
wire _05542_;
wire _05543_;
wire _05544_;
wire _05545_;
wire _05546_;
wire _05547_;
wire _05548_;
wire _05549_;
wire _05550_;
wire _05551_;
wire _05552_;
wire _05553_;
wire _05554_;
wire _05555_;
wire _05556_;
wire _05557_;
wire _05558_;
wire _05559_;
wire _05560_;
wire _05561_;
wire _05562_;
wire _05563_;
wire _05564_;
wire _05565_;
wire _05566_;
wire _05567_;
wire _05568_;
wire _05569_;
wire _05570_;
wire _05571_;
wire _05572_;
wire _05573_;
wire _05574_;
wire _05575_;
wire _05576_;
wire _05577_;
wire _05578_;
wire _05579_;
wire _05580_;
wire _05581_;
wire _05582_;
wire _05583_;
wire _05584_;
wire _05585_;
wire _05586_;
wire _05587_;
wire _05588_;
wire _05589_;
wire _05590_;
wire _05591_;
wire _05592_;
wire _05593_;
wire _05594_;
wire _05595_;
wire _05596_;
wire _05597_;
wire _05598_;
wire _05599_;
wire _05600_;
wire _05601_;
wire _05602_;
wire _05603_;
wire _05604_;
wire _05605_;
wire _05606_;
wire _05607_;
wire _05608_;
wire _05609_;
wire _05610_;
wire _05611_;
wire _05612_;
wire _05613_;
wire _05614_;
wire _05615_;
wire _05616_;
wire _05617_;
wire _05618_;
wire _05619_;
wire _05620_;
wire _05621_;
wire _05622_;
wire _05623_;
wire _05624_;
wire _05625_;
wire _05626_;
wire _05627_;
wire _05628_;
wire _05629_;
wire _05630_;
wire _05631_;
wire _05632_;
wire _05633_;
wire _05634_;
wire _05635_;
wire _05636_;
wire _05637_;
wire _05638_;
wire _05639_;
wire _05640_;
wire _05641_;
wire _05642_;
wire _05643_;
wire _05644_;
wire _05645_;
wire _05646_;
wire _05647_;
wire _05648_;
wire _05649_;
wire _05650_;
wire _05651_;
wire _05652_;
wire _05653_;
wire _05654_;
wire _05655_;
wire _05656_;
wire _05657_;
wire _05658_;
wire _05659_;
wire _05660_;
wire _05661_;
wire _05662_;
wire _05663_;
wire _05664_;
wire _05665_;
wire _05666_;
wire _05667_;
wire _05668_;
wire _05669_;
wire _05670_;
wire _05671_;
wire _05672_;
wire _05673_;
wire _05674_;
wire _05675_;
wire _05676_;
wire _05677_;
wire _05678_;
wire _05679_;
wire _05680_;
wire _05681_;
wire _05682_;
wire _05683_;
wire _05684_;
wire _05685_;
wire _05686_;
wire _05687_;
wire _05688_;
wire _05689_;
wire _05690_;
wire _05691_;
wire _05692_;
wire _05693_;
wire _05694_;
wire _05695_;
wire _05696_;
wire _05697_;
wire _05698_;
wire _05699_;
wire _05700_;
wire _05701_;
wire _05702_;
wire _05703_;
wire _05704_;
wire _05705_;
wire _05706_;
wire _05707_;
wire _05708_;
wire _05709_;
wire _05710_;
wire _05711_;
wire _05712_;
wire _05713_;
wire _05714_;
wire _05715_;
wire _05716_;
wire _05717_;
wire _05718_;
wire _05719_;
wire _05720_;
wire _05721_;
wire _05722_;
wire _05723_;
wire _05724_;
wire _05725_;
wire _05726_;
wire _05727_;
wire _05728_;
wire _05729_;
wire _05730_;
wire _05731_;
wire _05732_;
wire _05733_;
wire _05734_;
wire _05735_;
wire _05736_;
wire _05737_;
wire _05738_;
wire _05739_;
wire _05740_;
wire _05741_;
wire _05742_;
wire _05743_;
wire _05744_;
wire _05745_;
wire _05746_;
wire _05747_;
wire _05748_;
wire _05749_;
wire _05750_;
wire _05751_;
wire _05752_;
wire _05753_;
wire _05754_;
wire _05755_;
wire _05756_;
wire _05757_;
wire _05758_;
wire _05759_;
wire _05760_;
wire _05761_;
wire _05762_;
wire _05763_;
wire _05764_;
wire _05765_;
wire _05766_;
wire _05767_;
wire _05768_;
wire _05769_;
wire _05770_;
wire _05771_;
wire _05772_;
wire _05773_;
wire _05774_;
wire _05775_;
wire _05776_;
wire _05777_;
wire _05778_;
wire _05779_;
wire _05780_;
wire _05781_;
wire _05782_;
wire _05783_;
wire _05784_;
wire _05785_;
wire _05786_;
wire _05787_;
wire _05788_;
wire _05789_;
wire _05790_;
wire _05791_;
wire _05792_;
wire _05793_;
wire _05794_;
wire _05795_;
wire _05796_;
wire _05797_;
wire _05798_;
wire _05799_;
wire _05800_;
wire _05801_;
wire _05802_;
wire _05803_;
wire _05804_;
wire _05805_;
wire _05806_;
wire _05807_;
wire _05808_;
wire _05809_;
wire _05810_;
wire _05811_;
wire _05812_;
wire _05813_;
wire _05814_;
wire _05815_;
wire _05816_;
wire _05817_;
wire _05818_;
wire _05819_;
wire _05820_;
wire _05821_;
wire _05822_;
wire _05823_;
wire _05824_;
wire _05825_;
wire _05826_;
wire _05827_;
wire _05828_;
wire _05829_;
wire _05830_;
wire _05831_;
wire _05832_;
wire _05833_;
wire _05834_;
wire _05835_;
wire _05836_;
wire _05837_;
wire _05838_;
wire _05839_;
wire _05840_;
wire _05841_;
wire _05842_;
wire _05843_;
wire _05844_;
wire _05845_;
wire _05846_;
wire _05847_;
wire _05848_;
wire _05849_;
wire _05850_;
wire _05851_;
wire _05852_;
wire _05853_;
wire _05854_;
wire _05855_;
wire _05856_;
wire _05857_;
wire _05858_;
wire _05859_;
wire _05860_;
wire _05861_;
wire _05862_;
wire _05863_;
wire _05864_;
wire _05865_;
wire _05866_;
wire _05867_;
wire _05868_;
wire _05869_;
wire _05870_;
wire _05871_;
wire _05872_;
wire _05873_;
wire _05874_;
wire _05875_;
wire _05876_;
wire _05877_;
wire _05878_;
wire _05879_;
wire _05880_;
wire _05881_;
wire _05882_;
wire _05883_;
wire _05884_;
wire _05885_;
wire _05886_;
wire _05887_;
wire _05888_;
wire _05889_;
wire _05890_;
wire _05891_;
wire _05892_;
wire _05893_;
wire _05894_;
wire _05895_;
wire _05896_;
wire _05897_;
wire _05898_;
wire _05899_;
wire _05900_;
wire _05901_;
wire _05902_;
wire _05903_;
wire _05904_;
wire _05905_;
wire _05906_;
wire _05907_;
wire _05908_;
wire _05909_;
wire _05910_;
wire _05911_;
wire _05912_;
wire _05913_;
wire _05914_;
wire _05915_;
wire _05916_;
wire _05917_;
wire _05918_;
wire _05919_;
wire _05920_;
wire _05921_;
wire _05922_;
wire _05923_;
wire _05924_;
wire _05925_;
wire _05926_;
wire _05927_;
wire _05928_;
wire _05929_;
wire _05930_;
wire _05931_;
wire _05932_;
wire _05933_;
wire _05934_;
wire _05935_;
wire _05936_;
wire _05937_;
wire _05938_;
wire _05939_;
wire _05940_;
wire _05941_;
wire _05942_;
wire _05943_;
wire _05944_;
wire _05945_;
wire _05946_;
wire _05947_;
wire _05948_;
wire _05949_;
wire _05950_;
wire _05951_;
wire _05952_;
wire _05953_;
wire _05954_;
wire _05955_;
wire _05956_;
wire _05957_;
wire _05958_;
wire _05959_;
wire _05960_;
wire _05961_;
wire _05962_;
wire _05963_;
wire _05964_;
wire _05965_;
wire _05966_;
wire _05967_;
wire _05968_;
wire _05969_;
wire _05970_;
wire _05971_;
wire _05972_;
wire _05973_;
wire _05974_;
wire _05975_;
wire _05976_;
wire _05977_;
wire _05978_;
wire _05979_;
wire _05980_;
wire _05981_;
wire _05982_;
wire _05983_;
wire _05984_;
wire _05985_;
wire _05986_;
wire _05987_;
wire _05988_;
wire _05989_;
wire _05990_;
wire _05991_;
wire _05992_;
wire _05993_;
wire _05994_;
wire _05995_;
wire _05996_;
wire _05997_;
wire _05998_;
wire _05999_;
wire _06000_;
wire _06001_;
wire _06002_;
wire _06003_;
wire _06004_;
wire _06005_;
wire _06006_;
wire _06007_;
wire _06008_;
wire _06009_;
wire _06010_;
wire _06011_;
wire _06012_;
wire _06013_;
wire _06014_;
wire _06015_;
wire _06016_;
wire _06017_;
wire _06018_;
wire _06019_;
wire _06020_;
wire _06021_;
wire _06022_;
wire _06023_;
wire _06024_;
wire _06025_;
wire _06026_;
wire _06027_;
wire _06028_;
wire _06029_;
wire _06030_;
wire _06031_;
wire _06032_;
wire _06033_;
wire _06034_;
wire _06035_;
wire _06036_;
wire _06037_;
wire _06038_;
wire _06039_;
wire _06040_;
wire _06041_;
wire _06042_;
wire _06043_;
wire _06044_;
wire _06045_;
wire _06046_;
wire _06047_;
wire _06048_;
wire _06049_;
wire _06050_;
wire _06051_;
wire _06052_;
wire _06053_;
wire _06054_;
wire _06055_;
wire _06056_;
wire _06057_;
wire _06058_;
wire _06059_;
wire _06060_;
wire _06061_;
wire _06062_;
wire _06063_;
wire _06064_;
wire _06065_;
wire _06066_;
wire _06067_;
wire _06068_;
wire _06069_;
wire _06070_;
wire _06071_;
wire _06072_;
wire _06073_;
wire _06074_;
wire _06075_;
wire _06076_;
wire _06077_;
wire _06078_;
wire _06079_;
wire _06080_;
wire _06081_;
wire _06082_;
wire _06083_;
wire _06084_;
wire _06085_;
wire _06086_;
wire _06087_;
wire _06088_;
wire _06089_;
wire _06090_;
wire _06091_;
wire _06092_;
wire _06093_;
wire _06094_;
wire _06095_;
wire _06096_;
wire _06097_;
wire _06098_;
wire _06099_;
wire _06100_;
wire _06101_;
wire _06102_;
wire _06103_;
wire _06104_;
wire _06105_;
wire _06106_;
wire _06107_;
wire _06108_;
wire _06109_;
wire _06110_;
wire _06111_;
wire _06112_;
wire _06113_;
wire _06114_;
wire _06115_;
wire _06116_;
wire _06117_;
wire _06118_;
wire _06119_;
wire _06120_;
wire _06121_;
wire _06122_;
wire _06123_;
wire _06124_;
wire _06125_;
wire _06126_;
wire _06127_;
wire _06128_;
wire _06129_;
wire _06130_;
wire _06131_;
wire _06132_;
wire _06133_;
wire _06134_;
wire _06135_;
wire _06136_;
wire _06137_;
wire _06138_;
wire _06139_;
wire _06140_;
wire _06141_;
wire _06142_;
wire _06143_;
wire _06144_;
wire _06145_;
wire _06146_;
wire _06147_;
wire _06148_;
wire _06149_;
wire _06150_;
wire _06151_;
wire _06152_;
wire _06153_;
wire _06154_;
wire _06155_;
wire _06156_;
wire _06157_;
wire _06158_;
wire _06159_;
wire _06160_;
wire _06161_;
wire _06162_;
wire _06163_;
wire _06164_;
wire _06165_;
wire _06166_;
wire _06167_;
wire _06168_;
wire _06169_;
wire _06170_;
wire _06171_;
wire _06172_;
wire _06173_;
wire _06174_;
wire _06175_;
wire _06176_;
wire _06177_;
wire _06178_;
wire _06179_;
wire _06180_;
wire _06181_;
wire _06182_;
wire _06183_;
wire _06184_;
wire _06185_;
wire _06186_;
wire _06187_;
wire _06188_;
wire _06189_;
wire _06190_;
wire _06191_;
wire _06192_;
wire _06193_;
wire _06194_;
wire _06195_;
wire _06196_;
wire _06197_;
wire _06198_;
wire _06199_;
wire _06200_;
wire _06201_;
wire _06202_;
wire _06203_;
wire _06204_;
wire _06205_;
wire _06206_;
wire _06207_;
wire _06208_;
wire _06209_;
wire _06210_;
wire _06211_;
wire _06212_;
wire _06213_;
wire _06214_;
wire _06215_;
wire _06216_;
wire _06217_;
wire _06218_;
wire _06219_;
wire _06220_;
wire _06221_;
wire _06222_;
wire _06223_;
wire _06224_;
wire _06225_;
wire _06226_;
wire _06227_;
wire _06228_;
wire _06229_;
wire _06230_;
wire _06231_;
wire _06232_;
wire _06233_;
wire _06234_;
wire _06235_;
wire _06236_;
wire _06237_;
wire _06238_;
wire _06239_;
wire _06240_;
wire _06241_;
wire _06242_;
wire _06243_;
wire _06244_;
wire _06245_;
wire _06246_;
wire _06247_;
wire _06248_;
wire _06249_;
wire _06250_;
wire _06251_;
wire _06252_;
wire _06253_;
wire _06254_;
wire _06255_;
wire _06256_;
wire _06257_;
wire _06258_;
wire _06259_;
wire _06260_;
wire _06261_;
wire _06262_;
wire _06263_;
wire _06264_;
wire _06265_;
wire _06266_;
wire _06267_;
wire _06268_;
wire _06269_;
wire _06270_;
wire _06271_;
wire _06272_;
wire _06273_;
wire _06274_;
wire _06275_;
wire _06276_;
wire _06277_;
wire _06278_;
wire _06279_;
wire _06280_;
wire _06281_;
wire _06282_;
wire _06283_;
wire _06284_;
wire _06285_;
wire _06286_;
wire _06287_;
wire _06288_;
wire _06289_;
wire _06290_;
wire _06291_;
wire _06292_;
wire _06293_;
wire _06294_;
wire _06295_;
wire _06296_;
wire _06297_;
wire _06298_;
wire _06299_;
wire _06300_;
wire _06301_;
wire _06302_;
wire _06303_;
wire _06304_;
wire _06305_;
wire _06306_;
wire _06307_;
wire _06308_;
wire _06309_;
wire _06310_;
wire _06311_;
wire _06312_;
wire _06313_;
wire _06314_;
wire _06315_;
wire _06316_;
wire _06317_;
wire _06318_;
wire _06319_;
wire _06320_;
wire _06321_;
wire _06322_;
wire _06323_;
wire _06324_;
wire _06325_;
wire _06326_;
wire _06327_;
wire _06328_;
wire _06329_;
wire _06330_;
wire _06331_;
wire _06332_;
wire _06333_;
wire _06334_;
wire _06335_;
wire _06336_;
wire _06337_;
wire _06338_;
wire _06339_;
wire _06340_;
wire _06341_;
wire _06342_;
wire _06343_;
wire _06344_;
wire _06345_;
wire _06346_;
wire _06347_;
wire _06348_;
wire _06349_;
wire _06350_;
wire _06351_;
wire _06352_;
wire _06353_;
wire _06354_;
wire _06355_;
wire _06356_;
wire _06357_;
wire _06358_;
wire _06359_;
wire _06360_;
wire _06361_;
wire _06362_;
wire _06363_;
wire _06364_;
wire _06365_;
wire _06366_;
wire _06367_;
wire _06368_;
wire _06369_;
wire _06370_;
wire _06371_;
wire _06372_;
wire _06373_;
wire _06374_;
wire _06375_;
wire _06376_;
wire _06377_;
wire _06378_;
wire _06379_;
wire _06380_;
wire _06381_;
wire _06382_;
wire _06383_;
wire _06384_;
wire _06385_;
wire _06386_;
wire _06387_;
wire _06388_;
wire _06389_;
wire _06390_;
wire _06391_;
wire _06392_;
wire _06393_;
wire _06394_;
wire _06395_;
wire _06396_;
wire _06397_;
wire _06398_;
wire _06399_;
wire _06400_;
wire _06401_;
wire _06402_;
wire _06403_;
wire _06404_;
wire _06405_;
wire _06406_;
wire _06407_;
wire _06408_;
wire _06409_;
wire _06410_;
wire _06411_;
wire _06412_;
wire _06413_;
wire _06414_;
wire _06415_;
wire _06416_;
wire _06417_;
wire _06418_;
wire _06419_;
wire _06420_;
wire _06421_;
wire _06422_;
wire _06423_;
wire _06424_;
wire _06425_;
wire _06426_;
wire _06427_;
wire _06428_;
wire _06429_;
wire _06430_;
wire _06431_;
wire _06432_;
wire _06433_;
wire _06434_;
wire _06435_;
wire _06436_;
wire _06437_;
wire _06438_;
wire _06439_;
wire _06440_;
wire _06441_;
wire _06442_;
wire _06443_;
wire _06444_;
wire _06445_;
wire _06446_;
wire _06447_;
wire _06448_;
wire _06449_;
wire _06450_;
wire _06451_;
wire _06452_;
wire _06453_;
wire _06454_;
wire _06455_;
wire _06456_;
wire _06457_;
wire _06458_;
wire _06459_;
wire _06460_;
wire _06461_;
wire _06462_;
wire _06463_;
wire _06464_;
wire _06465_;
wire _06466_;
wire _06467_;
wire _06468_;
wire _06469_;
wire _06470_;
wire _06471_;
wire _06472_;
wire _06473_;
wire _06474_;
wire _06475_;
wire _06476_;
wire _06477_;
wire _06478_;
wire _06479_;
wire _06480_;
wire _06481_;
wire _06482_;
wire _06483_;
wire _06484_;
wire _06485_;
wire _06486_;
wire _06487_;
wire _06488_;
wire _06489_;
wire _06490_;
wire _06491_;
wire _06492_;
wire _06493_;
wire _06494_;
wire _06495_;
wire _06496_;
wire _06497_;
wire _06498_;
wire _06499_;
wire _06500_;
wire _06501_;
wire _06502_;
wire _06503_;
wire _06504_;
wire _06505_;
wire _06506_;
wire _06507_;
wire _06508_;
wire _06509_;
wire _06510_;
wire _06511_;
wire _06512_;
wire _06513_;
wire _06514_;
wire _06515_;
wire _06516_;
wire _06517_;
wire _06518_;
wire _06519_;
wire _06520_;
wire _06521_;
wire _06522_;
wire _06523_;
wire _06524_;
wire _06525_;
wire _06526_;
wire _06527_;
wire _06528_;
wire _06529_;
wire _06530_;
wire _06531_;
wire _06532_;
wire _06533_;
wire _06534_;
wire _06535_;
wire _06536_;
wire _06537_;
wire _06538_;
wire _06539_;
wire _06540_;
wire _06541_;
wire _06542_;
wire _06543_;
wire _06544_;
wire _06545_;
wire _06546_;
wire _06547_;
wire _06548_;
wire _06549_;
wire _06550_;
wire _06551_;
wire _06552_;
wire _06553_;
wire _06554_;
wire _06555_;
wire _06556_;
wire _06557_;
wire _06558_;
wire _06559_;
wire _06560_;
wire _06561_;
wire _06562_;
wire _06563_;
wire _06564_;
wire _06565_;
wire _06566_;
wire _06567_;
wire _06568_;
wire _06569_;
wire _06570_;
wire _06571_;
wire _06572_;
wire _06573_;
wire _06574_;
wire _06575_;
wire _06576_;
wire _06577_;
wire _06578_;
wire _06579_;
wire _06580_;
wire _06581_;
wire _06582_;
wire _06583_;
wire _06584_;
wire _06585_;
wire _06586_;
wire _06587_;
wire _06588_;
wire _06589_;
wire _06590_;
wire _06591_;
wire _06592_;
wire _06593_;
wire _06594_;
wire _06595_;
wire _06596_;
wire _06597_;
wire _06598_;
wire _06599_;
wire _06600_;
wire _06601_;
wire _06602_;
wire _06603_;
wire _06604_;
wire _06605_;
wire _06606_;
wire _06607_;
wire _06608_;
wire _06609_;
wire _06610_;
wire _06611_;
wire _06612_;
wire _06613_;
wire _06614_;
wire _06615_;
wire _06616_;
wire _06617_;
wire _06618_;
wire _06619_;
wire _06620_;
wire _06621_;
wire _06622_;
wire _06623_;
wire _06624_;
wire _06625_;
wire _06626_;
wire _06627_;
wire _06628_;
wire _06629_;
wire _06630_;
wire _06631_;
wire _06632_;
wire _06633_;
wire _06634_;
wire _06635_;
wire _06636_;
wire _06637_;
wire _06638_;
wire _06639_;
wire _06640_;
wire _06641_;
wire _06642_;
wire _06643_;
wire _06644_;
wire _06645_;
wire _06646_;
wire _06647_;
wire _06648_;
wire _06649_;
wire _06650_;
wire _06651_;
wire _06652_;
wire _06653_;
wire _06654_;
wire _06655_;
wire _06656_;
wire _06657_;
wire _06658_;
wire _06659_;
wire _06660_;
wire _06661_;
wire _06662_;
wire _06663_;
wire _06664_;
wire _06665_;
wire _06666_;
wire _06667_;
wire _06668_;
wire _06669_;
wire _06670_;
wire _06671_;
wire _06672_;
wire _06673_;
wire _06674_;
wire _06675_;
wire _06676_;
wire _06677_;
wire _06678_;
wire _06679_;
wire _06680_;
wire _06681_;
wire _06682_;
wire _06683_;
wire _06684_;
wire _06685_;
wire _06686_;
wire _06687_;
wire _06688_;
wire _06689_;
wire _06690_;
wire _06691_;
wire _06692_;
wire _06693_;
wire _06694_;
wire _06695_;
wire _06696_;
wire _06697_;
wire _06698_;
wire _06699_;
wire _06700_;
wire _06701_;
wire _06702_;
wire _06703_;
wire _06704_;
wire _06705_;
wire _06706_;
wire _06707_;
wire _06708_;
wire _06709_;
wire _06710_;
wire _06711_;
wire _06712_;
wire _06713_;
wire _06714_;
wire _06715_;
wire _06716_;
wire _06717_;
wire _06718_;
wire _06719_;
wire _06720_;
wire _06721_;
wire _06722_;
wire _06723_;
wire _06724_;
wire _06725_;
wire _06726_;
wire _06727_;
wire _06728_;
wire _06729_;
wire _06730_;
wire _06731_;
wire _06732_;
wire _06733_;
wire _06734_;
wire _06735_;
wire _06736_;
wire _06737_;
wire _06738_;
wire _06739_;
wire _06740_;
wire _06741_;
wire _06742_;
wire _06743_;
wire _06744_;
wire _06745_;
wire _06746_;
wire _06747_;
wire _06748_;
wire _06749_;
wire _06750_;
wire _06751_;
wire _06752_;
wire _06753_;
wire _06754_;
wire _06755_;
wire _06756_;
wire _06757_;
wire _06758_;
wire _06759_;
wire _06760_;
wire _06761_;
wire _06762_;
wire _06763_;
wire _06764_;
wire _06765_;
wire _06766_;
wire _06767_;
wire _06768_;
wire _06769_;
wire _06770_;
wire _06771_;
wire _06772_;
wire _06773_;
wire _06774_;
wire _06775_;
wire _06776_;
wire _06777_;
wire _06778_;
wire _06779_;
wire _06780_;
wire _06781_;
wire _06782_;
wire _06783_;
wire _06784_;
wire _06785_;
wire _06786_;
wire _06787_;
wire _06788_;
wire _06789_;
wire _06790_;
wire _06791_;
wire _06792_;
wire _06793_;
wire _06794_;
wire _06795_;
wire _06796_;
wire _06797_;
wire _06798_;
wire _06799_;
wire _06800_;
wire _06801_;
wire _06802_;
wire _06803_;
wire _06804_;
wire _06805_;
wire _06806_;
wire _06807_;
wire _06808_;
wire _06809_;
wire _06810_;
wire _06811_;
wire _06812_;
wire _06813_;
wire _06814_;
wire _06815_;
wire _06816_;
wire _06817_;
wire _06818_;
wire _06819_;
wire _06820_;
wire _06821_;
wire _06822_;
wire _06823_;
wire _06824_;
wire _06825_;
wire _06826_;
wire _06827_;
wire _06828_;
wire _06829_;
wire _06830_;
wire _06831_;
wire _06832_;
wire _06833_;
wire _06834_;
wire _06835_;
wire _06836_;
wire _06837_;
wire _06838_;
wire _06839_;
wire _06840_;
wire _06841_;
wire _06842_;
wire _06843_;
wire _06844_;
wire _06845_;
wire _06846_;
wire _06847_;
wire _06848_;
wire _06849_;
wire _06850_;
wire _06851_;
wire _06852_;
wire _06853_;
wire _06854_;
wire _06855_;
wire _06856_;
wire _06857_;
wire _06858_;
wire _06859_;
wire _06860_;
wire _06861_;
wire _06862_;
wire _06863_;
wire _06864_;
wire _06865_;
wire _06866_;
wire _06867_;
wire _06868_;
wire _06869_;
wire _06870_;
wire _06871_;
wire _06872_;
wire _06873_;
wire _06874_;
wire _06875_;
wire _06876_;
wire _06877_;
wire _06878_;
wire _06879_;
wire _06880_;
wire _06881_;
wire _06882_;
wire _06883_;
wire _06884_;
wire _06885_;
wire _06886_;
wire _06887_;
wire _06888_;
wire _06889_;
wire _06890_;
wire _06891_;
wire _06892_;
wire _06893_;
wire _06894_;
wire _06895_;
wire _06896_;
wire _06897_;
wire _06898_;
wire _06899_;
wire _06900_;
wire _06901_;
wire _06902_;
wire _06903_;
wire _06904_;
wire _06905_;
wire _06906_;
wire _06907_;
wire _06908_;
wire _06909_;
wire _06910_;
wire _06911_;
wire _06912_;
wire _06913_;
wire _06914_;
wire _06915_;
wire _06916_;
wire _06917_;
wire _06918_;
wire _06919_;
wire _06920_;
wire _06921_;
wire _06922_;
wire _06923_;
wire _06924_;
wire _06925_;
wire _06926_;
wire _06927_;
wire _06928_;
wire _06929_;
wire _06930_;
wire _06931_;
wire _06932_;
wire _06933_;
wire _06934_;
wire _06935_;
wire _06936_;
wire _06937_;
wire _06938_;
wire _06939_;
wire _06940_;
wire _06941_;
wire _06942_;
wire _06943_;
wire _06944_;
wire _06945_;
wire _06946_;
wire _06947_;
wire _06948_;
wire _06949_;
wire _06950_;
wire _06951_;
wire _06952_;
wire _06953_;
wire _06954_;
wire _06955_;
wire _06956_;
wire _06957_;
wire _06958_;
wire _06959_;
wire _06960_;
wire _06961_;
wire _06962_;
wire _06963_;
wire _06964_;
wire _06965_;
wire _06966_;
wire _06967_;
wire _06968_;
wire _06969_;
wire _06970_;
wire _06971_;
wire _06972_;
wire _06973_;
wire _06974_;
wire _06975_;
wire _06976_;
wire _06977_;
wire _06978_;
wire _06979_;
wire _06980_;
wire _06981_;
wire _06982_;
wire _06983_;
wire _06984_;
wire _06985_;
wire _06986_;
wire _06987_;
wire _06988_;
wire _06989_;
wire _06990_;
wire _06991_;
wire _06992_;
wire _06993_;
wire _06994_;
wire _06995_;
wire _06996_;
wire _06997_;
wire _06998_;
wire _06999_;
wire _07000_;
wire _07001_;
wire _07002_;
wire _07003_;
wire _07004_;
wire _07005_;
wire _07006_;
wire _07007_;
wire _07008_;
wire _07009_;
wire _07010_;
wire _07011_;
wire _07012_;
wire _07013_;
wire _07014_;
wire _07015_;
wire _07016_;
wire _07017_;
wire _07018_;
wire _07019_;
wire _07020_;
wire _07021_;
wire _07022_;
wire _07023_;
wire _07024_;
wire _07025_;
wire _07026_;
wire _07027_;
wire _07028_;
wire _07029_;
wire _07030_;
wire _07031_;
wire _07032_;
wire _07033_;
wire _07034_;
wire _07035_;
wire _07036_;
wire _07037_;
wire _07038_;
wire _07039_;
wire _07040_;
wire _07041_;
wire _07042_;
wire _07043_;
wire _07044_;
wire _07045_;
wire _07046_;
wire _07047_;
wire _07048_;
wire _07049_;
wire _07050_;
wire _07051_;
wire _07052_;
wire _07053_;
wire _07054_;
wire _07055_;
wire _07056_;
wire _07057_;
wire _07058_;
wire _07059_;
wire _07060_;
wire _07061_;
wire _07062_;
wire _07063_;
wire _07064_;
wire _07065_;
wire _07066_;
wire _07067_;
wire _07068_;
wire _07069_;
wire _07070_;
wire _07071_;
wire _07072_;
wire _07073_;
wire _07074_;
wire _07075_;
wire _07076_;
wire _07077_;
wire _07078_;
wire _07079_;
wire _07080_;
wire _07081_;
wire _07082_;
wire _07083_;
wire _07084_;
wire _07085_;
wire _07086_;
wire _07087_;
wire _07088_;
wire _07089_;
wire _07090_;
wire _07091_;
wire _07092_;
wire _07093_;
wire _07094_;
wire _07095_;
wire _07096_;
wire _07097_;
wire _07098_;
wire _07099_;
wire _07100_;
wire _07101_;
wire _07102_;
wire _07103_;
wire _07104_;
wire _07105_;
wire _07106_;
wire _07107_;
wire _07108_;
wire _07109_;
wire _07110_;
wire _07111_;
wire _07112_;
wire _07113_;
wire _07114_;
wire _07115_;
wire _07116_;
wire _07117_;
wire _07118_;
wire _07119_;
wire _07120_;
wire _07121_;
wire _07122_;
wire _07123_;
wire _07124_;
wire _07125_;
wire _07126_;
wire _07127_;
wire _07128_;
wire _07129_;
wire _07130_;
wire _07131_;
wire _07132_;
wire _07133_;
wire _07134_;
wire _07135_;
wire _07136_;
wire _07137_;
wire _07138_;
wire _07139_;
wire _07140_;
wire _07141_;
wire _07142_;
wire _07143_;
wire _07144_;
wire _07145_;
wire _07146_;
wire _07147_;
wire _07148_;
wire _07149_;
wire _07150_;
wire _07151_;
wire _07152_;
wire _07153_;
wire _07154_;
wire _07155_;
wire _07156_;
wire _07157_;
wire _07158_;
wire _07159_;
wire _07160_;
wire _07161_;
wire _07162_;
wire _07163_;
wire _07164_;
wire _07165_;
wire _07166_;
wire _07167_;
wire _07168_;
wire _07169_;
wire _07170_;
wire _07171_;
wire _07172_;
wire _07173_;
wire _07174_;
wire _07175_;
wire _07176_;
wire _07177_;
wire _07178_;
wire _07179_;
wire _07180_;
wire _07181_;
wire _07182_;
wire _07183_;
wire _07184_;
wire _07185_;
wire _07186_;
wire _07187_;
wire _07188_;
wire _07189_;
wire _07190_;
wire _07191_;
wire _07192_;
wire _07193_;
wire _07194_;
wire _07195_;
wire _07196_;
wire _07197_;
wire _07198_;
wire _07199_;
wire _07200_;
wire _07201_;
wire _07202_;
wire _07203_;
wire _07204_;
wire _07205_;
wire _07206_;
wire _07207_;
wire _07208_;
wire _07209_;
wire _07210_;
wire _07211_;
wire _07212_;
wire _07213_;
wire _07214_;
wire _07215_;
wire _07216_;
wire _07217_;
wire _07218_;
wire _07219_;
wire _07220_;
wire _07221_;
wire _07222_;
wire _07223_;
wire _07224_;
wire _07225_;
wire _07226_;
wire _07227_;
wire _07228_;
wire _07229_;
wire _07230_;
wire _07231_;
wire _07232_;
wire _07233_;
wire _07234_;
wire _07235_;
wire _07236_;
wire _07237_;
wire _07238_;
wire _07239_;
wire _07240_;
wire _07241_;
wire _07242_;
wire _07243_;
wire _07244_;
wire _07245_;
wire _07246_;
wire _07247_;
wire _07248_;
wire _07249_;
wire _07250_;
wire _07251_;
wire _07252_;
wire _07253_;
wire _07254_;
wire _07255_;
wire _07256_;
wire _07257_;
wire _07258_;
wire _07259_;
wire _07260_;
wire _07261_;
wire _07262_;
wire _07263_;
wire _07264_;
wire _07265_;
wire _07266_;
wire _07267_;
wire _07268_;
wire _07269_;
wire _07270_;
wire _07271_;
wire _07272_;
wire _07273_;
wire _07274_;
wire _07275_;
wire _07276_;
wire _07277_;
wire _07278_;
wire _07279_;
wire _07280_;
wire _07281_;
wire _07282_;
wire _07283_;
wire _07284_;
wire _07285_;
wire _07286_;
wire _07287_;
wire _07288_;
wire _07289_;
wire _07290_;
wire _07291_;
wire _07292_;
wire _07293_;
wire _07294_;
wire _07295_;
wire _07296_;
wire _07297_;
wire _07298_;
wire _07299_;
wire _07300_;
wire _07301_;
wire _07302_;
wire _07303_;
wire _07304_;
wire _07305_;
wire _07306_;
wire _07307_;
wire _07308_;
wire _07309_;
wire _07310_;
wire _07311_;
wire _07312_;
wire _07313_;
wire _07314_;
wire _07315_;
wire _07316_;
wire _07317_;
wire _07318_;
wire _07319_;
wire _07320_;
wire _07321_;
wire _07322_;
wire _07323_;
wire _07324_;
wire _07325_;
wire _07326_;
wire _07327_;
wire _07328_;
wire _07329_;
wire _07330_;
wire _07331_;
wire _07332_;
wire _07333_;
wire _07334_;
wire _07335_;
wire _07336_;
wire _07337_;
wire _07338_;
wire _07339_;
wire _07340_;
wire _07341_;
wire _07342_;
wire _07343_;
wire _07344_;
wire _07345_;
wire _07346_;
wire _07347_;
wire _07348_;
wire _07349_;
wire _07350_;
wire _07351_;
wire _07352_;
wire _07353_;
wire _07354_;
wire _07355_;
wire _07356_;
wire _07357_;
wire _07358_;
wire _07359_;
wire _07360_;
wire _07361_;
wire _07362_;
wire _07363_;
wire _07364_;
wire _07365_;
wire _07366_;
wire _07367_;
wire _07368_;
wire _07369_;
wire _07370_;
wire _07371_;
wire _07372_;
wire _07373_;
wire _07374_;
wire _07375_;
wire _07376_;
wire _07377_;
wire _07378_;
wire _07379_;
wire _07380_;
wire _07381_;
wire _07382_;
wire _07383_;
wire _07384_;
wire _07385_;
wire _07386_;
wire _07387_;
wire _07388_;
wire _07389_;
wire _07390_;
wire _07391_;
wire _07392_;
wire _07393_;
wire _07394_;
wire _07395_;
wire _07396_;
wire _07397_;
wire _07398_;
wire _07399_;
wire _07400_;
wire _07401_;
wire _07402_;
wire _07403_;
wire _07404_;
wire _07405_;
wire _07406_;
wire _07407_;
wire _07408_;
wire _07409_;
wire _07410_;
wire _07411_;
wire _07412_;
wire _07413_;
wire _07414_;
wire _07415_;
wire _07416_;
wire _07417_;
wire _07418_;
wire _07419_;
wire _07420_;
wire _07421_;
wire _07422_;
wire _07423_;
wire _07424_;
wire _07425_;
wire _07426_;
wire _07427_;
wire _07428_;
wire _07429_;
wire _07430_;
wire _07431_;
wire _07432_;
wire _07433_;
wire _07434_;
wire _07435_;
wire _07436_;
wire _07437_;
wire _07438_;
wire _07439_;
wire _07440_;
wire _07441_;
wire _07442_;
wire _07443_;
wire _07444_;
wire _07445_;
wire _07446_;
wire _07447_;
wire _07448_;
wire _07449_;
wire _07450_;
wire _07451_;
wire _07452_;
wire _07453_;
wire _07454_;
wire _07455_;
wire _07456_;
wire _07457_;
wire _07458_;
wire _07459_;
wire _07460_;
wire _07461_;
wire _07462_;
wire _07463_;
wire _07464_;
wire _07465_;
wire _07466_;
wire _07467_;
wire _07468_;
wire _07469_;
wire _07470_;
wire _07471_;
wire _07472_;
wire _07473_;
wire _07474_;
wire _07475_;
wire _07476_;
wire _07477_;
wire _07478_;
wire _07479_;
wire _07480_;
wire _07481_;
wire _07482_;
wire _07483_;
wire _07484_;
wire _07485_;
wire _07486_;
wire _07487_;
wire _07488_;
wire _07489_;
wire _07490_;
wire _07491_;
wire _07492_;
wire _07493_;
wire _07494_;
wire _07495_;
wire _07496_;
wire _07497_;
wire _07498_;
wire _07499_;
wire _07500_;
wire _07501_;
wire _07502_;
wire _07503_;
wire _07504_;
wire _07505_;
wire _07506_;
wire _07507_;
wire _07508_;
wire _07509_;
wire _07510_;
wire _07511_;
wire _07512_;
wire _07513_;
wire _07514_;
wire _07515_;
wire _07516_;
wire _07517_;
wire _07518_;
wire _07519_;
wire _07520_;
wire _07521_;
wire _07522_;
wire _07523_;
wire _07524_;
wire _07525_;
wire _07526_;
wire _07527_;
wire _07528_;
wire _07529_;
wire _07530_;
wire _07531_;
wire _07532_;
wire _07533_;
wire _07534_;
wire _07535_;
wire _07536_;
wire _07537_;
wire _07538_;
wire _07539_;
wire _07540_;
wire _07541_;
wire _07542_;
wire _07543_;
wire _07544_;
wire _07545_;
wire _07546_;
wire _07547_;
wire _07548_;
wire _07549_;
wire _07550_;
wire _07551_;
wire _07552_;
wire _07553_;
wire _07554_;
wire _07555_;
wire _07556_;
wire _07557_;
wire _07558_;
wire _07559_;
wire _07560_;
wire _07561_;
wire _07562_;
wire _07563_;
wire _07564_;
wire _07565_;
wire _07566_;
wire _07567_;
wire _07568_;
wire _07569_;
wire _07570_;
wire _07571_;
wire _07572_;
wire _07573_;
wire _07574_;
wire _07575_;
wire _07576_;
wire _07577_;
wire _07578_;
wire _07579_;
wire _07580_;
wire _07581_;
wire _07582_;
wire _07583_;
wire _07584_;
wire _07585_;
wire _07586_;
wire _07587_;
wire _07588_;
wire _07589_;
wire _07590_;
wire _07591_;
wire _07592_;
wire _07593_;
wire _07594_;
wire _07595_;
wire _07596_;
wire _07597_;
wire _07598_;
wire _07599_;
wire _07600_;
wire _07601_;
wire _07602_;
wire _07603_;
wire _07604_;
wire _07605_;
wire _07606_;
wire _07607_;
wire _07608_;
wire _07609_;
wire _07610_;
wire _07611_;
wire _07612_;
wire _07613_;
wire _07614_;
wire _07615_;
wire _07616_;
wire _07617_;
wire _07618_;
wire _07619_;
wire _07620_;
wire _07621_;
wire _07622_;
wire _07623_;
wire _07624_;
wire _07625_;
wire _07626_;
wire _07627_;
wire _07628_;
wire _07629_;
wire _07630_;
wire _07631_;
wire _07632_;
wire _07633_;
wire _07634_;
wire _07635_;
wire _07636_;
wire _07637_;
wire _07638_;
wire _07639_;
wire _07640_;
wire _07641_;
wire _07642_;
wire _07643_;
wire _07644_;
wire _07645_;
wire _07646_;
wire _07647_;
wire _07648_;
wire _07649_;
wire _07650_;
wire _07651_;
wire _07652_;
wire _07653_;
wire _07654_;
wire _07655_;
wire _07656_;
wire _07657_;
wire _07658_;
wire _07659_;
wire _07660_;
wire _07661_;
wire _07662_;
wire _07663_;
wire _07664_;
wire _07665_;
wire _07666_;
wire _07667_;
wire _07668_;
wire _07669_;
wire _07670_;
wire _07671_;
wire _07672_;
wire _07673_;
wire _07674_;
wire _07675_;
wire _07676_;
wire _07677_;
wire _07678_;
wire _07679_;
wire _07680_;
wire _07681_;
wire _07682_;
wire _07683_;
wire _07684_;
wire _07685_;
wire _07686_;
wire _07687_;
wire _07688_;
wire _07689_;
wire _07690_;
wire _07691_;
wire _07692_;
wire _07693_;
wire _07694_;
wire _07695_;
wire _07696_;
wire _07697_;
wire _07698_;
wire _07699_;
wire _07700_;
wire _07701_;
wire _07702_;
wire _07703_;
wire _07704_;
wire _07705_;
wire _07706_;
wire _07707_;
wire _07708_;
wire _07709_;
wire _07710_;
wire _07711_;
wire _07712_;
wire _07713_;
wire _07714_;
wire _07715_;
wire _07716_;
wire _07717_;
wire _07718_;
wire _07719_;
wire _07720_;
wire _07721_;
wire _07722_;
wire _07723_;
wire _07724_;
wire _07725_;
wire _07726_;
wire _07727_;
wire _07728_;
wire _07729_;
wire _07730_;
wire _07731_;
wire _07732_;
wire _07733_;
wire _07734_;
wire _07735_;
wire _07736_;
wire _07737_;
wire _07738_;
wire _07739_;
wire _07740_;
wire _07741_;
wire _07742_;
wire _07743_;
wire _07744_;
wire _07745_;
wire _07746_;
wire _07747_;
wire _07748_;
wire _07749_;
wire _07750_;
wire _07751_;
wire _07752_;
wire _07753_;
wire _07754_;
wire _07755_;
wire _07756_;
wire _07757_;
wire _07758_;
wire _07759_;
wire _07760_;
wire _07761_;
wire _07762_;
wire _07763_;
wire _07764_;
wire _07765_;
wire _07766_;
wire _07767_;
wire _07768_;
wire _07769_;
wire _07770_;
wire _07771_;
wire _07772_;
wire _07773_;
wire _07774_;
wire _07775_;
wire _07776_;
wire _07777_;
wire _07778_;
wire _07779_;
wire _07780_;
wire _07781_;
wire _07782_;
wire _07783_;
wire _07784_;
wire _07785_;
wire _07786_;
wire _07787_;
wire _07788_;
wire _07789_;
wire _07790_;
wire _07791_;
wire _07792_;
wire _07793_;
wire _07794_;
wire _07795_;
wire _07796_;
wire _07797_;
wire _07798_;
wire _07799_;
wire _07800_;
wire _07801_;
wire _07802_;
wire _07803_;
wire _07804_;
wire _07805_;
wire _07806_;
wire _07807_;
wire _07808_;
wire _07809_;
wire _07810_;
wire _07811_;
wire _07812_;
wire _07813_;
wire _07814_;
wire _07815_;
wire _07816_;
wire _07817_;
wire _07818_;
wire _07819_;
wire _07820_;
wire _07821_;
wire _07822_;
wire _07823_;
wire _07824_;
wire _07825_;
wire _07826_;
wire _07827_;
wire _07828_;
wire _07829_;
wire _07830_;
wire _07831_;
wire _07832_;
wire _07833_;
wire _07834_;
wire _07835_;
wire _07836_;
wire _07837_;
wire _07838_;
wire _07839_;
wire _07840_;
wire _07841_;
wire _07842_;
wire _07843_;
wire _07844_;
wire _07845_;
wire _07846_;
wire _07847_;
wire _07848_;
wire _07849_;
wire _07850_;
wire _07851_;
wire _07852_;
wire _07853_;
wire _07854_;
wire _07855_;
wire _07856_;
wire _07857_;
wire _07858_;
wire _07859_;
wire _07860_;
wire _07861_;
wire _07862_;
wire _07863_;
wire _07864_;
wire _07865_;
wire _07866_;
wire _07867_;
wire _07868_;
wire _07869_;
wire _07870_;
wire _07871_;
wire _07872_;
wire _07873_;
wire _07874_;
wire _07875_;
wire _07876_;
wire _07877_;
wire _07878_;
wire _07879_;
wire _07880_;
wire _07881_;
wire _07882_;
wire _07883_;
wire _07884_;
wire _07885_;
wire _07886_;
wire _07887_;
wire _07888_;
wire _07889_;
wire _07890_;
wire _07891_;
wire _07892_;
wire _07893_;
wire _07894_;
wire _07895_;
wire _07896_;
wire _07897_;
wire _07898_;
wire _07899_;
wire _07900_;
wire _07901_;
wire _07902_;
wire _07903_;
wire _07904_;
wire _07905_;
wire _07906_;
wire _07907_;
wire _07908_;
wire _07909_;
wire _07910_;
wire _07911_;
wire _07912_;
wire _07913_;
wire _07914_;
wire _07915_;
wire _07916_;
wire _07917_;
wire _07918_;
wire _07919_;
wire _07920_;
wire _07921_;
wire _07922_;
wire _07923_;
wire _07924_;
wire _07925_;
wire _07926_;
wire _07927_;
wire _07928_;
wire _07929_;
wire _07930_;
wire _07931_;
wire _07932_;
wire _07933_;
wire _07934_;
wire _07935_;
wire _07936_;
wire _07937_;
wire _07938_;
wire _07939_;
wire _07940_;
wire _07941_;
wire _07942_;
wire _07943_;
wire _07944_;
wire _07945_;
wire _07946_;
wire _07947_;
wire _07948_;
wire _07949_;
wire _07950_;
wire _07951_;
wire _07952_;
wire _07953_;
wire _07954_;
wire _07955_;
wire _07956_;
wire _07957_;
wire _07958_;
wire _07959_;
wire _07960_;
wire _07961_;
wire _07962_;
wire _07963_;
wire _07964_;
wire _07965_;
wire _07966_;
wire _07967_;
wire _07968_;
wire _07969_;
wire _07970_;
wire _07971_;
wire _07972_;
wire _07973_;
wire _07974_;
wire _07975_;
wire _07976_;
wire _07977_;
wire _07978_;
wire _07979_;
wire _07980_;
wire _07981_;
wire _07982_;
wire _07983_;
wire _07984_;
wire _07985_;
wire _07986_;
wire _07987_;
wire _07988_;
wire _07989_;
wire _07990_;
wire _07991_;
wire _07992_;
wire _07993_;
wire _07994_;
wire _07995_;
wire _07996_;
wire _07997_;
wire _07998_;
wire _07999_;
wire _08000_;
wire _08001_;
wire _08002_;
wire _08003_;
wire _08004_;
wire _08005_;
wire _08006_;
wire _08007_;
wire _08008_;
wire _08009_;
wire _08010_;
wire _08011_;
wire _08012_;
wire _08013_;
wire _08014_;
wire _08015_;
wire _08016_;
wire _08017_;
wire _08018_;
wire _08019_;
wire _08020_;
wire _08021_;
wire _08022_;
wire _08023_;
wire _08024_;
wire _08025_;
wire _08026_;
wire _08027_;
wire _08028_;
wire _08029_;
wire _08030_;
wire _08031_;
wire _08032_;
wire _08033_;
wire _08034_;
wire _08035_;
wire _08036_;
wire _08037_;
wire _08038_;
wire _08039_;
wire _08040_;
wire _08041_;
wire _08042_;
wire _08043_;
wire _08044_;
wire _08045_;
wire _08046_;
wire _08047_;
wire _08048_;
wire _08049_;
wire _08050_;
wire _08051_;
wire _08052_;
wire _08053_;
wire _08054_;
wire _08055_;
wire _08056_;
wire _08057_;
wire _08058_;
wire _08059_;
wire _08060_;
wire _08061_;
wire _08062_;
wire _08063_;
wire _08064_;
wire _08065_;
wire _08066_;
wire _08067_;
wire _08068_;
wire _08069_;
wire _08070_;
wire _08071_;
wire _08072_;
wire _08073_;
wire _08074_;
wire _08075_;
wire _08076_;
wire _08077_;
wire _08078_;
wire _08079_;
wire _08080_;
wire _08081_;
wire _08082_;
wire _08083_;
wire _08084_;
wire _08085_;
wire _08086_;
wire _08087_;
wire _08088_;
wire _08089_;
wire _08090_;
wire _08091_;
wire _08092_;
wire _08093_;
wire _08094_;
wire _08095_;
wire _08096_;
wire _08097_;
wire _08098_;
wire _08099_;
wire _08100_;
wire _08101_;
wire _08102_;
wire _08103_;
wire _08104_;
wire _08105_;
wire _08106_;
wire _08107_;
wire _08108_;
wire _08109_;
wire _08110_;
wire _08111_;
wire _08112_;
wire _08113_;
wire _08114_;
wire _08115_;
wire _08116_;
wire _08117_;
wire _08118_;
wire _08119_;
wire _08120_;
wire _08121_;
wire _08122_;
wire _08123_;
wire _08124_;
wire _08125_;
wire _08126_;
wire _08127_;
wire _08128_;
wire _08129_;
wire _08130_;
wire _08131_;
wire _08132_;
wire _08133_;
wire _08134_;
wire _08135_;
wire _08136_;
wire _08137_;
wire _08138_;
wire _08139_;
wire _08140_;
wire _08141_;
wire _08142_;
wire _08143_;
wire _08144_;
wire _08145_;
wire _08146_;
wire _08147_;
wire _08148_;
wire _08149_;
wire _08150_;
wire _08151_;
wire _08152_;
wire _08153_;
wire _08154_;
wire _08155_;
wire _08156_;
wire _08157_;
wire _08158_;
wire _08159_;
wire _08160_;
wire _08161_;
wire _08162_;
wire _08163_;
wire _08164_;
wire _08165_;
wire _08166_;
wire _08167_;
wire _08168_;
wire _08169_;
wire _08170_;
wire _08171_;
wire _08172_;
wire _08173_;
wire _08174_;
wire _08175_;
wire _08176_;
wire _08177_;
wire _08178_;
wire _08179_;
wire _08180_;
wire _08181_;
wire _08182_;
wire _08183_;
wire _08184_;
wire _08185_;
wire _08186_;
wire _08187_;
wire _08188_;
wire _08189_;
wire _08190_;
wire _08191_;
wire _08192_;
wire _08193_;
wire _08194_;
wire _08195_;
wire _08196_;
wire _08197_;
wire _08198_;
wire _08199_;
wire _08200_;
wire _08201_;
wire _08202_;
wire _08203_;
wire _08204_;
wire _08205_;
wire _08206_;
wire _08207_;
wire _08208_;
wire _08209_;
wire _08210_;
wire _08211_;
wire _08212_;
wire _08213_;
wire _08214_;
wire _08215_;
wire _08216_;
wire _08217_;
wire _08218_;
wire _08219_;
wire _08220_;
wire _08221_;
wire _08222_;
wire _08223_;
wire _08224_;
wire _08225_;
wire _08226_;
wire _08227_;
wire _08228_;
wire _08229_;
wire _08230_;
wire _08231_;
wire _08232_;
wire _08233_;
wire _08234_;
wire _08235_;
wire _08236_;
wire _08237_;
wire _08238_;
wire _08239_;
wire _08240_;
wire _08241_;
wire _08242_;
wire _08243_;
wire _08244_;
wire _08245_;
wire _08246_;
wire _08247_;
wire _08248_;
wire _08249_;
wire _08250_;
wire _08251_;
wire _08252_;
wire _08253_;
wire _08254_;
wire _08255_;
wire _08256_;
wire _08257_;
wire _08258_;
wire _08259_;
wire _08260_;
wire _08261_;
wire _08262_;
wire _08263_;
wire _08264_;
wire _08265_;
wire _08266_;
wire _08267_;
wire _08268_;
wire _08269_;
wire _08270_;
wire _08271_;
wire _08272_;
wire _08273_;
wire _08274_;
wire _08275_;
wire _08276_;
wire _08277_;
wire _08278_;
wire _08279_;
wire _08280_;
wire _08281_;
wire _08282_;
wire _08283_;
wire _08284_;
wire _08285_;
wire _08286_;
wire _08287_;
wire _08288_;
wire _08289_;
wire _08290_;
wire _08291_;
wire _08292_;
wire _08293_;
wire _08294_;
wire _08295_;
wire _08296_;
wire _08297_;
wire _08298_;
wire _08299_;
wire _08300_;
wire _08301_;
wire _08302_;
wire _08303_;
wire _08304_;
wire _08305_;
wire _08306_;
wire _08307_;
wire _08308_;
wire _08309_;
wire _08310_;
wire _08311_;
wire _08312_;
wire _08313_;
wire _08314_;
wire _08315_;
wire _08316_;
wire _08317_;
wire _08318_;
wire _08319_;
wire _08320_;
wire _08321_;
wire _08322_;
wire _08323_;
wire _08324_;
wire _08325_;
wire _08326_;
wire _08327_;
wire _08328_;
wire _08329_;
wire _08330_;
wire _08331_;
wire _08332_;
wire _08333_;
wire _08334_;
wire _08335_;
wire _08336_;
wire _08337_;
wire _08338_;
wire _08339_;
wire _08340_;
wire _08341_;
wire _08342_;
wire _08343_;
wire _08344_;
wire _08345_;
wire _08346_;
wire _08347_;
wire _08348_;
wire _08349_;
wire _08350_;
wire _08351_;
wire _08352_;
wire _08353_;
wire _08354_;
wire _08355_;
wire _08356_;
wire _08357_;
wire _08358_;
wire _08359_;
wire _08360_;
wire _08361_;
wire _08362_;
wire _08363_;
wire _08364_;
wire _08365_;
wire _08366_;
wire _08367_;
wire _08368_;
wire _08369_;
wire _08370_;
wire _08371_;
wire _08372_;
wire _08373_;
wire _08374_;
wire _08375_;
wire _08376_;
wire _08377_;
wire _08378_;
wire _08379_;
wire _08380_;
wire _08381_;
wire _08382_;
wire _08383_;
wire _08384_;
wire _08385_;
wire _08386_;
wire _08387_;
wire _08388_;
wire _08389_;
wire _08390_;
wire _08391_;
wire _08392_;
wire _08393_;
wire _08394_;
wire _08395_;
wire _08396_;
wire _08397_;
wire _08398_;
wire _08399_;
wire _08400_;
wire _08401_;
wire _08402_;
wire _08403_;
wire _08404_;
wire _08405_;
wire _08406_;
wire _08407_;
wire _08408_;
wire _08409_;
wire _08410_;
wire _08411_;
wire _08412_;
wire _08413_;
wire _08414_;
wire _08415_;
wire _08416_;
wire _08417_;
wire _08418_;
wire _08419_;
wire _08420_;
wire _08421_;
wire _08422_;
wire _08423_;
wire _08424_;
wire _08425_;
wire _08426_;
wire _08427_;
wire _08428_;
wire _08429_;
wire _08430_;
wire _08431_;
wire _08432_;
wire _08433_;
wire _08434_;
wire _08435_;
wire _08436_;
wire _08437_;
wire _08438_;
wire _08439_;
wire _08440_;
wire _08441_;
wire _08442_;
wire _08443_;
wire _08444_;
wire _08445_;
wire _08446_;
wire _08447_;
wire _08448_;
wire _08449_;
wire _08450_;
wire _08451_;
wire _08452_;
wire _08453_;
wire _08454_;
wire _08455_;
wire _08456_;
wire _08457_;
wire _08458_;
wire _08459_;
wire _08460_;
wire _08461_;
wire _08462_;
wire _08463_;
wire _08464_;
wire _08465_;
wire _08466_;
wire _08467_;
wire _08468_;
wire _08469_;
wire _08470_;
wire _08471_;
wire _08472_;
wire _08473_;
wire _08474_;
wire _08475_;
wire _08476_;
wire _08477_;
wire _08478_;
wire _08479_;
wire _08480_;
wire _08481_;
wire _08482_;
wire _08483_;
wire _08484_;
wire _08485_;
wire _08486_;
wire _08487_;
wire _08488_;
wire _08489_;
wire _08490_;
wire _08491_;
wire _08492_;
wire _08493_;
wire _08494_;
wire _08495_;
wire _08496_;
wire _08497_;
wire _08498_;
wire _08499_;
wire _08500_;
wire _08501_;
wire _08502_;
wire _08503_;
wire _08504_;
wire _08505_;
wire _08506_;
wire _08507_;
wire _08508_;
wire _08509_;
wire _08510_;
wire _08511_;
wire _08512_;
wire _08513_;
wire _08514_;
wire _08515_;
wire _08516_;
wire _08517_;
wire _08518_;
wire _08519_;
wire _08520_;
wire _08521_;
wire _08522_;
wire _08523_;
wire _08524_;
wire _08525_;
wire _08526_;
wire _08527_;
wire _08528_;
wire _08529_;
wire _08530_;
wire _08531_;
wire _08532_;
wire _08533_;
wire _08534_;
wire _08535_;
wire _08536_;
wire _08537_;
wire _08538_;
wire _08539_;
wire _08540_;
wire _08541_;
wire _08542_;
wire _08543_;
wire _08544_;
wire _08545_;
wire _08546_;
wire _08547_;
wire _08548_;
wire _08549_;
wire _08550_;
wire _08551_;
wire _08552_;
wire _08553_;
wire _08554_;
wire _08555_;
wire _08556_;
wire _08557_;
wire _08558_;
wire _08559_;
wire _08560_;
wire _08561_;
wire _08562_;
wire _08563_;
wire _08564_;
wire _08565_;
wire _08566_;
wire _08567_;
wire _08568_;
wire _08569_;
wire _08570_;
wire _08571_;
wire _08572_;
wire _08573_;
wire _08574_;
wire _08575_;
wire _08576_;
wire _08577_;
wire _08578_;
wire _08579_;
wire _08580_;
wire _08581_;
wire _08582_;
wire _08583_;
wire _08584_;
wire _08585_;
wire _08586_;
wire _08587_;
wire _08588_;
wire _08589_;
wire _08590_;
wire _08591_;
wire _08592_;
wire _08593_;
wire _08594_;
wire _08595_;
wire _08596_;
wire _08597_;
wire _08598_;
wire _08599_;
wire _08600_;
wire _08601_;
wire _08602_;
wire _08603_;
wire _08604_;
wire _08605_;
wire _08606_;
wire _08607_;
wire _08608_;
wire _08609_;
wire _08610_;
wire _08611_;
wire _08612_;
wire _08613_;
wire _08614_;
wire _08615_;
wire _08616_;
wire _08617_;
wire _08618_;
wire _08619_;
wire _08620_;
wire _08621_;
wire _08622_;
wire _08623_;
wire _08624_;
wire _08625_;
wire _08626_;
wire _08627_;
wire _08628_;
wire _08629_;
wire _08630_;
wire _08631_;
wire _08632_;
wire _08633_;
wire _08634_;
wire _08635_;
wire _08636_;
wire _08637_;
wire _08638_;
wire _08639_;
wire _08640_;
wire _08641_;
wire _08642_;
wire _08643_;
wire _08644_;
wire _08645_;
wire _08646_;
wire _08647_;
wire _08648_;
wire _08649_;
wire _08650_;
wire _08651_;
wire _08652_;
wire _08653_;
wire _08654_;
wire _08655_;
wire _08656_;
wire _08657_;
wire _08658_;
wire _08659_;
wire _08660_;
wire _08661_;
wire _08662_;
wire _08663_;
wire _08664_;
wire _08665_;
wire _08666_;
wire _08667_;
wire _08668_;
wire _08669_;
wire _08670_;
wire _08671_;
wire _08672_;
wire _08673_;
wire _08674_;
wire _08675_;
wire _08676_;
wire _08677_;
wire _08678_;
wire _08679_;
wire _08680_;
wire _08681_;
wire _08682_;
wire _08683_;
wire _08684_;
wire _08685_;
wire _08686_;
wire _08687_;
wire _08688_;
wire _08689_;
wire _08690_;
wire _08691_;
wire _08692_;
wire _08693_;
wire _08694_;
wire _08695_;
wire _08696_;
wire _08697_;
wire _08698_;
wire _08699_;
wire _08700_;
wire _08701_;
wire _08702_;
wire _08703_;
wire _08704_;
wire _08705_;
wire _08706_;
wire _08707_;
wire _08708_;
wire _08709_;
wire _08710_;
wire _08711_;
wire _08712_;
wire _08713_;
wire _08714_;
wire _08715_;
wire _08716_;
wire _08717_;
wire _08718_;
wire _08719_;
wire _08720_;
wire _08721_;
wire _08722_;
wire _08723_;
wire _08724_;
wire _08725_;
wire _08726_;
wire _08727_;
wire _08728_;
wire _08729_;
wire _08730_;
wire _08731_;
wire _08732_;
wire _08733_;
wire _08734_;
wire _08735_;
wire _08736_;
wire _08737_;
wire _08738_;
wire _08739_;
wire _08740_;
wire _08741_;
wire _08742_;
wire _08743_;
wire _08744_;
wire _08745_;
wire _08746_;
wire _08747_;
wire _08748_;
wire _08749_;
wire _08750_;
wire _08751_;
wire _08752_;
wire _08753_;
wire _08754_;
wire _08755_;
wire _08756_;
wire _08757_;
wire _08758_;
wire _08759_;
wire _08760_;
wire _08761_;
wire _08762_;
wire _08763_;
wire _08764_;
wire _08765_;
wire _08766_;
wire _08767_;
wire _08768_;
wire _08769_;
wire _08770_;
wire _08771_;
wire _08772_;
wire _08773_;
wire _08774_;
wire _08775_;
wire _08776_;
wire _08777_;
wire _08778_;
wire _08779_;
wire _08780_;
wire _08781_;
wire _08782_;
wire _08783_;
wire _08784_;
wire _08785_;
wire _08786_;
wire _08787_;
wire _08788_;
wire _08789_;
wire _08790_;
wire _08791_;
wire _08792_;
wire _08793_;
wire _08794_;
wire _08795_;
wire _08796_;
wire _08797_;
wire _08798_;
wire _08799_;
wire _08800_;
wire _08801_;
wire _08802_;
wire _08803_;
wire _08804_;
wire _08805_;
wire _08806_;
wire _08807_;
wire _08808_;
wire _08809_;
wire _08810_;
wire _08811_;
wire _08812_;
wire _08813_;
wire _08814_;
wire _08815_;
wire _08816_;
wire _08817_;
wire _08818_;
wire _08819_;
wire _08820_;
wire _08821_;
wire _08822_;
wire _08823_;
wire _08824_;
wire _08825_;
wire _08826_;
wire _08827_;
wire _08828_;
wire _08829_;
wire _08830_;
wire _08831_;
wire _08832_;
wire _08833_;
wire _08834_;
wire _08835_;
wire _08836_;
wire _08837_;
wire _08838_;
wire _08839_;
wire _08840_;
wire _08841_;
wire _08842_;
wire _08843_;
wire _08844_;
wire _08845_;
wire _08846_;
wire _08847_;
wire _08848_;
wire _08849_;
wire _08850_;
wire _08851_;
wire _08852_;
wire _08853_;
wire _08854_;
wire _08855_;
wire _08856_;
wire _08857_;
wire _08858_;
wire _08859_;
wire _08860_;
wire _08861_;
wire _08862_;
wire _08863_;
wire _08864_;
wire _08865_;
wire _08866_;
wire _08867_;
wire _08868_;
wire _08869_;
wire _08870_;
wire _08871_;
wire _08872_;
wire _08873_;
wire _08874_;
wire _08875_;
wire _08876_;
wire _08877_;
wire _08878_;
wire _08879_;
wire _08880_;
wire _08881_;
wire _08882_;
wire _08883_;
wire _08884_;
wire _08885_;
wire _08886_;
wire _08887_;
wire _08888_;
wire _08889_;
wire _08890_;
wire _08891_;
wire _08892_;
wire _08893_;
wire _08894_;
wire _08895_;
wire _08896_;
wire _08897_;
wire _08898_;
wire _08899_;
wire _08900_;
wire _08901_;
wire _08902_;
wire _08903_;
wire _08904_;
wire _08905_;
wire _08906_;
wire _08907_;
wire _08908_;
wire _08909_;
wire _08910_;
wire _08911_;
wire _08912_;
wire _08913_;
wire _08914_;
wire _08915_;
wire _08916_;
wire _08917_;
wire _08918_;
wire _08919_;
wire _08920_;
wire _08921_;
wire _08922_;
wire _08923_;
wire _08924_;
wire _08925_;
wire _08926_;
wire _08927_;
wire _08928_;
wire _08929_;
wire _08930_;
wire _08931_;
wire _08932_;
wire _08933_;
wire _08934_;
wire _08935_;
wire _08936_;
wire _08937_;
wire _08938_;
wire _08939_;
wire _08940_;
wire _08941_;
wire _08942_;
wire _08943_;
wire _08944_;
wire _08945_;
wire _08946_;
wire _08947_;
wire _08948_;
wire _08949_;
wire _08950_;
wire _08951_;
wire _08952_;
wire _08953_;
wire _08954_;
wire _08955_;
wire _08956_;
wire _08957_;
wire _08958_;
wire _08959_;
wire _08960_;
wire _08961_;
wire _08962_;
wire _08963_;
wire _08964_;
wire _08965_;
wire _08966_;
wire _08967_;
wire _08968_;
wire _08969_;
wire _08970_;
wire _08971_;
wire _08972_;
wire _08973_;
wire _08974_;
wire _08975_;
wire _08976_;
wire _08977_;
wire _08978_;
wire _08979_;
wire _08980_;
wire _08981_;
wire _08982_;
wire _08983_;
wire _08984_;
wire _08985_;
wire _08986_;
wire _08987_;
wire _08988_;
wire _08989_;
wire _08990_;
wire _08991_;
wire _08992_;
wire _08993_;
wire _08994_;
wire _08995_;
wire _08996_;
wire _08997_;
wire _08998_;
wire _08999_;
wire _09000_;
wire _09001_;
wire _09002_;
wire _09003_;
wire _09004_;
wire _09005_;
wire _09006_;
wire _09007_;
wire _09008_;
wire _09009_;
wire _09010_;
wire _09011_;
wire _09012_;
wire _09013_;
wire _09014_;
wire _09015_;
wire _09016_;
wire _09017_;
wire _09018_;
wire _09019_;
wire _09020_;
wire _09021_;
wire _09022_;
wire _09023_;
wire _09024_;
wire _09025_;
wire _09026_;
wire _09027_;
wire _09028_;
wire _09029_;
wire _09030_;
wire _09031_;
wire _09032_;
wire _09033_;
wire _09034_;
wire _09035_;
wire _09036_;
wire _09037_;
wire _09038_;
wire _09039_;
wire _09040_;
wire _09041_;
wire _09042_;
wire _09043_;
wire _09044_;
wire _09045_;
wire _09046_;
wire _09047_;
wire _09048_;
wire _09049_;
wire _09050_;
wire _09051_;
wire _09052_;
wire _09053_;
wire _09054_;
wire _09055_;
wire _09056_;
wire _09057_;
wire _09058_;
wire _09059_;
wire _09060_;
wire _09061_;
wire _09062_;
wire _09063_;
wire _09064_;
wire _09065_;
wire _09066_;
wire _09067_;
wire _09068_;
wire _09069_;
wire _09070_;
wire _09071_;
wire _09072_;
wire _09073_;
wire _09074_;
wire _09075_;
wire _09076_;
wire _09077_;
wire _09078_;
wire _09079_;
wire _09080_;
wire _09081_;
wire _09082_;
wire _09083_;
wire _09084_;
wire _09085_;
wire _09086_;
wire _09087_;
wire _09088_;
wire _09089_;
wire _09090_;
wire _09091_;
wire _09092_;
wire _09093_;
wire _09094_;
wire _09095_;
wire _09096_;
wire _09097_;
wire _09098_;
wire _09099_;
wire _09100_;
wire _09101_;
wire _09102_;
wire _09103_;
wire _09104_;
wire _09105_;
wire _09106_;
wire _09107_;
wire _09108_;
wire _09109_;
wire _09110_;
wire _09111_;
wire _09112_;
wire _09113_;
wire _09114_;
wire _09115_;
wire _09116_;
wire _09117_;
wire _09118_;
wire _09119_;
wire _09120_;
wire _09121_;
wire _09122_;
wire _09123_;
wire _09124_;
wire _09125_;
wire _09126_;
wire _09127_;
wire _09128_;
wire _09129_;
wire _09130_;
wire _09131_;
wire _09132_;
wire _09133_;
wire _09134_;
wire _09135_;
wire _09136_;
wire _09137_;
wire _09138_;
wire _09139_;
wire _09140_;
wire _09141_;
wire _09142_;
wire _09143_;
wire _09144_;
wire _09145_;
wire _09146_;
wire _09147_;
wire _09148_;
wire _09149_;
wire _09150_;
wire _09151_;
wire _09152_;
wire _09153_;
wire _09154_;
wire _09155_;
wire _09156_;
wire _09157_;
wire _09158_;
wire _09159_;
wire _09160_;
wire _09161_;
wire _09162_;
wire _09163_;
wire _09164_;
wire _09165_;
wire _09166_;
wire _09167_;
wire _09168_;
wire _09169_;
wire _09170_;
wire _09171_;
wire _09172_;
wire _09173_;
wire _09174_;
wire _09175_;
wire _09176_;
wire _09177_;
wire _09178_;
wire _09179_;
wire _09180_;
wire _09181_;
wire _09182_;
wire _09183_;
wire _09184_;
wire _09185_;
wire _09186_;
wire _09187_;
wire _09188_;
wire _09189_;
wire _09190_;
wire _09191_;
wire _09192_;
wire _09193_;
wire _09194_;
wire _09195_;
wire _09196_;
wire _09197_;
wire _09198_;
wire _09199_;
wire _09200_;
wire _09201_;
wire _09202_;
wire _09203_;
wire _09204_;
wire _09205_;
wire _09206_;
wire _09207_;
wire _09208_;
wire _09209_;
wire _09210_;
wire _09211_;
wire _09212_;
wire _09213_;
wire _09214_;
wire _09215_;
wire _09216_;
wire _09217_;
wire _09218_;
wire _09219_;
wire _09220_;
wire _09221_;
wire _09222_;
wire _09223_;
wire _09224_;
wire _09225_;
wire _09226_;
wire _09227_;
wire _09228_;
wire _09229_;
wire _09230_;
wire _09231_;
wire _09232_;
wire _09233_;
wire _09234_;
wire _09235_;
wire _09236_;
wire _09237_;
wire _09238_;
wire _09239_;
wire _09240_;
wire _09241_;
wire _09242_;
wire _09243_;
wire _09244_;
wire _09245_;
wire _09246_;
wire _09247_;
wire _09248_;
wire _09249_;
wire _09250_;
wire _09251_;
wire _09252_;
wire _09253_;
wire _09254_;
wire _09255_;
wire _09256_;
wire _09257_;
wire _09258_;
wire _09259_;
wire _09260_;
wire _09261_;
wire _09262_;
wire _09263_;
wire _09264_;
wire _09265_;
wire _09266_;
wire _09267_;
wire _09268_;
wire _09269_;
wire _09270_;
wire _09271_;
wire _09272_;
wire _09273_;
wire _09274_;
wire _09275_;
wire _09276_;
wire _09277_;
wire _09278_;
wire _09279_;
wire _09280_;
wire _09281_;
wire _09282_;
wire _09283_;
wire _09284_;
wire _09285_;
wire _09286_;
wire _09287_;
wire _09288_;
wire _09289_;
wire _09290_;
wire _09291_;
wire _09292_;
wire _09293_;
wire _09294_;
wire _09295_;
wire _09296_;
wire _09297_;
wire _09298_;
wire _09299_;
wire _09300_;
wire _09301_;
wire _09302_;
wire _09303_;
wire _09304_;
wire _09305_;
wire _09306_;
wire _09307_;
wire _09308_;
wire _09309_;
wire _09310_;
wire _09311_;
wire _09312_;
wire _09313_;
wire _09314_;
wire _09315_;
wire _09316_;
wire _09317_;
wire _09318_;
wire _09319_;
wire _09320_;
wire _09321_;
wire _09322_;
wire _09323_;
wire _09324_;
wire _09325_;
wire _09326_;
wire _09327_;
wire _09328_;
wire _09329_;
wire _09330_;
wire _09331_;
wire _09332_;
wire _09333_;
wire _09334_;
wire _09335_;
wire _09336_;
wire _09337_;
wire _09338_;
wire _09339_;
wire _09340_;
wire _09341_;
wire _09342_;
wire _09343_;
wire _09344_;
wire _09345_;
wire _09346_;
wire _09347_;
wire _09348_;
wire _09349_;
wire _09350_;
wire _09351_;
wire _09352_;
wire _09353_;
wire _09354_;
wire _09355_;
wire _09356_;
wire _09357_;
wire _09358_;
wire _09359_;
wire _09360_;
wire _09361_;
wire _09362_;
wire _09363_;
wire _09364_;
wire _09365_;
wire _09366_;
wire _09367_;
wire _09368_;
wire _09369_;
wire _09370_;
wire _09371_;
wire _09372_;
wire _09373_;
wire _09374_;
wire _09375_;
wire _09376_;
wire _09377_;
wire _09378_;
wire _09379_;
wire _09380_;
wire _09381_;
wire _09382_;
wire _09383_;
wire _09384_;
wire _09385_;
wire _09386_;
wire _09387_;
wire _09388_;
wire _09389_;
wire _09390_;
wire _09391_;
wire _09392_;
wire _09393_;
wire _09394_;
wire _09395_;
wire _09396_;
wire _09397_;
wire _09398_;
wire _09399_;
wire _09400_;
wire _09401_;
wire _09402_;
wire _09403_;
wire _09404_;
wire _09405_;
wire _09406_;
wire _09407_;
wire _09408_;
wire _09409_;
wire _09410_;
wire _09411_;
wire _09412_;
wire _09413_;
wire _09414_;
wire _09415_;
wire _09416_;
wire _09417_;
wire _09418_;
wire _09419_;
wire _09420_;
wire _09421_;
wire _09422_;
wire _09423_;
wire _09424_;
wire _09425_;
wire _09426_;
wire _09427_;
wire _09428_;
wire _09429_;
wire _09430_;
wire _09431_;
wire _09432_;
wire _09433_;
wire _09434_;
wire _09435_;
wire _09436_;
wire _09437_;
wire _09438_;
wire _09439_;
wire _09440_;
wire _09441_;
wire _09442_;
wire _09443_;
wire _09444_;
wire _09445_;
wire _09446_;
wire _09447_;
wire _09448_;
wire _09449_;
wire _09450_;
wire _09451_;
wire _09452_;
wire _09453_;
wire _09454_;
wire _09455_;
wire _09456_;
wire _09457_;
wire _09458_;
wire _09459_;
wire _09460_;
wire _09461_;
wire _09462_;
wire _09463_;
wire _09464_;
wire _09465_;
wire _09466_;
wire _09467_;
wire _09468_;
wire _09469_;
wire _09470_;
wire _09471_;
wire _09472_;
wire _09473_;
wire _09474_;
wire _09475_;
wire _09476_;
wire _09477_;
wire _09478_;
wire _09479_;
wire _09480_;
wire _09481_;
wire _09482_;
wire _09483_;
wire _09484_;
wire _09485_;
wire _09486_;
wire _09487_;
wire _09488_;
wire _09489_;
wire _09490_;
wire _09491_;
wire _09492_;
wire _09493_;
wire _09494_;
wire _09495_;
wire _09496_;
wire _09497_;
wire _09498_;
wire _09499_;
wire _09500_;
wire _09501_;
wire _09502_;
wire _09503_;
wire _09504_;
wire _09505_;
wire _09506_;
wire _09507_;
wire _09508_;
wire _09509_;
wire _09510_;
wire _09511_;
wire _09512_;
wire _09513_;
wire _09514_;
wire _09515_;
wire _09516_;
wire _09517_;
wire _09518_;
wire _09519_;
wire _09520_;
wire _09521_;
wire _09522_;
wire _09523_;
wire _09524_;
wire _09525_;
wire _09526_;
wire _09527_;
wire _09528_;
wire _09529_;
wire _09530_;
wire _09531_;
wire _09532_;
wire _09533_;
wire _09534_;
wire _09535_;
wire _09536_;
wire _09537_;
wire _09538_;
wire _09539_;
wire _09540_;
wire _09541_;
wire _09542_;
wire _09543_;
wire _09544_;
wire _09545_;
wire _09546_;
wire _09547_;
wire _09548_;
wire _09549_;
wire _09550_;
wire _09551_;
wire _09552_;
wire _09553_;
wire _09554_;
wire _09555_;
wire _09556_;
wire _09557_;
wire _09558_;
wire _09559_;
wire _09560_;
wire _09561_;
wire _09562_;
wire _09563_;
wire _09564_;
wire _09565_;
wire _09566_;
wire _09567_;
wire _09568_;
wire _09569_;
wire _09570_;
wire _09571_;
wire _09572_;
wire _09573_;
wire _09574_;
wire _09575_;
wire _09576_;
wire _09577_;
wire _09578_;
wire _09579_;
wire _09580_;
wire _09581_;
wire _09582_;
wire _09583_;
wire _09584_;
wire _09585_;
wire _09586_;
wire _09587_;
wire _09588_;
wire _09589_;
wire _09590_;
wire _09591_;
wire _09592_;
wire _09593_;
wire _09594_;
wire _09595_;
wire _09596_;
wire _09597_;
wire _09598_;
wire _09599_;
wire _09600_;
wire _09601_;
wire _09602_;
wire _09603_;
wire _09604_;
wire _09605_;
wire _09606_;
wire _09607_;
wire _09608_;
wire _09609_;
wire _09610_;
wire _09611_;
wire _09612_;
wire _09613_;
wire _09614_;
wire _09615_;
wire _09616_;
wire _09617_;
wire _09618_;
wire _09619_;
wire _09620_;
wire _09621_;
wire _09622_;
wire _09623_;
wire _09624_;
wire _09625_;
wire _09626_;
wire _09627_;
wire _09628_;
wire _09629_;
wire _09630_;
wire _09631_;
wire _09632_;
wire _09633_;
wire _09634_;
wire _09635_;
wire _09636_;
wire _09637_;
wire _09638_;
wire _09639_;
wire _09640_;
wire _09641_;
wire _09642_;
wire _09643_;
wire _09644_;
wire _09645_;
wire _09646_;
wire _09647_;
wire _09648_;
wire _09649_;
wire _09650_;
wire _09651_;
wire _09652_;
wire _09653_;
wire _09654_;
wire _09655_;
wire _09656_;
wire _09657_;
wire _09658_;
wire _09659_;
wire _09660_;
wire _09661_;
wire _09662_;
wire _09663_;
wire _09664_;
wire _09665_;
wire _09666_;
wire _09667_;
wire _09668_;
wire _09669_;
wire _09670_;
wire _09671_;
wire _09672_;
wire _09673_;
wire _09674_;
wire _09675_;
wire _09676_;
wire _09677_;
wire _09678_;
wire _09679_;
wire _09680_;
wire _09681_;
wire _09682_;
wire _09683_;
wire _09684_;
wire _09685_;
wire _09686_;
wire _09687_;
wire _09688_;
wire _09689_;
wire _09690_;
wire _09691_;
wire _09692_;
wire _09693_;
wire _09694_;
wire _09695_;
wire _09696_;
wire _09697_;
wire _09698_;
wire _09699_;
wire _09700_;
wire _09701_;
wire _09702_;
wire _09703_;
wire _09704_;
wire _09705_;
wire _09706_;
wire _09707_;
wire _09708_;
wire _09709_;
wire _09710_;
wire _09711_;
wire _09712_;
wire _09713_;
wire _09714_;
wire _09715_;
wire _09716_;
wire _09717_;
wire _09718_;
wire _09719_;
wire _09720_;
wire _09721_;
wire _09722_;
wire _09723_;
wire _09724_;
wire _09725_;
wire _09726_;
wire _09727_;
wire _09728_;
wire _09729_;
wire _09730_;
wire _09731_;
wire _09732_;
wire _09733_;
wire _09734_;
wire _09735_;
wire _09736_;
wire _09737_;
wire _09738_;
wire _09739_;
wire _09740_;
wire _09741_;
wire _09742_;
wire _09743_;
wire _09744_;
wire _09745_;
wire _09746_;
wire _09747_;
wire _09748_;
wire _09749_;
wire _09750_;
wire _09751_;
wire _09752_;
wire _09753_;
wire _09754_;
wire _09755_;
wire _09756_;
wire _09757_;
wire _09758_;
wire _09759_;
wire _09760_;
wire _09761_;
wire _09762_;
wire _09763_;
wire _09764_;
wire _09765_;
wire _09766_;
wire _09767_;
wire _09768_;
wire _09769_;
wire _09770_;
wire _09771_;
wire _09772_;
wire _09773_;
wire _09774_;
wire _09775_;
wire _09776_;
wire _09777_;
wire _09778_;
wire _09779_;
wire _09780_;
wire _09781_;
wire _09782_;
wire _09783_;
wire _09784_;
wire _09785_;
wire _09786_;
wire _09787_;
wire _09788_;
wire _09789_;
wire _09790_;
wire _09791_;
wire _09792_;
wire _09793_;
wire _09794_;
wire _09795_;
wire _09796_;
wire _09797_;
wire _09798_;
wire _09799_;
wire _09800_;
wire _09801_;
wire _09802_;
wire _09803_;
wire _09804_;
wire _09805_;
wire _09806_;
wire _09807_;
wire _09808_;
wire _09809_;
wire _09810_;
wire _09811_;
wire _09812_;
wire _09813_;
wire _09814_;
wire _09815_;
wire _09816_;
wire _09817_;
wire _09818_;
wire _09819_;
wire _09820_;
wire _09821_;
wire _09822_;
wire _09823_;
wire _09824_;
wire _09825_;
wire _09826_;
wire _09827_;
wire _09828_;
wire _09829_;
wire _09830_;
wire _09831_;
wire _09832_;
wire _09833_;
wire _09834_;
wire _09835_;
wire _09836_;
wire _09837_;
wire _09838_;
wire _09839_;
wire _09840_;
wire _09841_;
wire _09842_;
wire _09843_;
wire _09844_;
wire _09845_;
wire _09846_;
wire _09847_;
wire _09848_;
wire _09849_;
wire _09850_;
wire _09851_;
wire _09852_;
wire _09853_;
wire _09854_;
wire _09855_;
wire _09856_;
wire _09857_;
wire _09858_;
wire _09859_;
wire _09860_;
wire _09861_;
wire _09862_;
wire _09863_;
wire _09864_;
wire _09865_;
wire _09866_;
wire _09867_;
wire _09868_;
wire _09869_;
wire _09870_;
wire _09871_;
wire _09872_;
wire _09873_;
wire _09874_;
wire _09875_;
wire _09876_;
wire _09877_;
wire _09878_;
wire _09879_;
wire _09880_;
wire _09881_;
wire _09882_;
wire _09883_;
wire _09884_;
wire _09885_;
wire _09886_;
wire _09887_;
wire _09888_;
wire _09889_;
wire _09890_;
wire _09891_;
wire _09892_;
wire _09893_;
wire _09894_;
wire _09895_;
wire _09896_;
wire _09897_;
wire _09898_;
wire _09899_;
wire _09900_;
wire _09901_;
wire _09902_;
wire _09903_;
wire _09904_;
wire _09905_;
wire _09906_;
wire _09907_;
wire _09908_;
wire _09909_;
wire _09910_;
wire _09911_;
wire _09912_;
wire _09913_;
wire _09914_;
wire _09915_;
wire _09916_;
wire _09917_;
wire _09918_;
wire _09919_;
wire _09920_;
wire _09921_;
wire _09922_;
wire _09923_;
wire _09924_;
wire _09925_;
wire _09926_;
wire _09927_;
wire _09928_;
wire _09929_;
wire _09930_;
wire _09931_;
wire _09932_;
wire _09933_;
wire _09934_;
wire _09935_;
wire _09936_;
wire _09937_;
wire _09938_;
wire _09939_;
wire _09940_;
wire _09941_;
wire _09942_;
wire _09943_;
wire _09944_;
wire _09945_;
wire _09946_;
wire _09947_;
wire _09948_;
wire _09949_;
wire _09950_;
wire _09951_;
wire _09952_;
wire _09953_;
wire _09954_;
wire _09955_;
wire _09956_;
wire _09957_;
wire _09958_;
wire _09959_;
wire _09960_;
wire _09961_;
wire _09962_;
wire _09963_;
wire _09964_;
wire _09965_;
wire _09966_;
wire _09967_;
wire _09968_;
wire _09969_;
wire _09970_;
wire _09971_;
wire _09972_;
wire _09973_;
wire _09974_;
wire _09975_;
wire _09976_;
wire _09977_;
wire _09978_;
wire _09979_;
wire _09980_;
wire _09981_;
wire _09982_;
wire _09983_;
wire _09984_;
wire _09985_;
wire _09986_;
wire _09987_;
wire _09988_;
wire _09989_;
wire _09990_;
wire _09991_;
wire _09992_;
wire _09993_;
wire _09994_;
wire _09995_;
wire _09996_;
wire _09997_;
wire _09998_;
wire _09999_;
wire _10000_;
wire _10001_;
wire _10002_;
wire _10003_;
wire _10004_;
wire _10005_;
wire _10006_;
wire _10007_;
wire _10008_;
wire _10009_;
wire _10010_;
wire _10011_;
wire _10012_;
wire _10013_;
wire _10014_;
wire _10015_;
wire _10016_;
wire _10017_;
wire _10018_;
wire _10019_;
wire _10020_;
wire _10021_;
wire _10022_;
wire _10023_;
wire _10024_;
wire _10025_;
wire _10026_;
wire _10027_;
wire _10028_;
wire _10029_;
wire _10030_;
wire _10031_;
wire _10032_;
wire _10033_;
wire _10034_;
wire _10035_;
wire _10036_;
wire _10037_;
wire _10038_;
wire _10039_;
wire _10040_;
wire _10041_;
wire _10042_;
wire _10043_;
wire _10044_;
wire _10045_;
wire _10046_;
wire _10047_;
wire _10048_;
wire _10049_;
wire _10050_;
wire _10051_;
wire _10052_;
wire _10053_;
wire _10054_;
wire _10055_;
wire _10056_;
wire _10057_;
wire _10058_;
wire _10059_;
wire _10060_;
wire _10061_;
wire _10062_;
wire _10063_;
wire _10064_;
wire _10065_;
wire _10066_;
wire _10067_;
wire _10068_;
wire _10069_;
wire _10070_;
wire _10071_;
wire _10072_;
wire _10073_;
wire _10074_;
wire _10075_;
wire _10076_;
wire _10077_;
wire _10078_;
wire _10079_;
wire _10080_;
wire _10081_;
wire _10082_;
wire _10083_;
wire _10084_;
wire _10085_;
wire _10086_;
wire _10087_;
wire _10088_;
wire _10089_;
wire _10090_;
wire _10091_;
wire _10092_;
wire _10093_;
wire _10094_;
wire _10095_;
wire _10096_;
wire _10097_;
wire _10098_;
wire _10099_;
wire _10100_;
wire _10101_;
wire _10102_;
wire _10103_;
wire _10104_;
wire _10105_;
wire _10106_;
wire _10107_;
wire _10108_;
wire _10109_;
wire _10110_;
wire _10111_;
wire _10112_;
wire _10113_;
wire _10114_;
wire _10115_;
wire _10116_;
wire _10117_;
wire _10118_;
wire _10119_;
wire _10120_;
wire _10121_;
wire _10122_;
wire _10123_;
wire _10124_;
wire _10125_;
wire _10126_;
wire _10127_;
wire _10128_;
wire _10129_;
wire _10130_;
wire _10131_;
wire _10132_;
wire _10133_;
wire _10134_;
wire _10135_;
wire _10136_;
wire _10137_;
wire _10138_;
wire _10139_;
wire _10140_;
wire _10141_;
wire _10142_;
wire _10143_;
wire _10144_;
wire _10145_;
wire _10146_;
wire _10147_;
wire _10148_;
wire _10149_;
wire _10150_;
wire _10151_;
wire _10152_;
wire _10153_;
wire _10154_;
wire _10155_;
wire _10156_;
wire _10157_;
wire _10158_;
wire _10159_;
wire _10160_;
wire _10161_;
wire _10162_;
wire _10163_;
wire _10164_;
wire _10165_;
wire _10166_;
wire _10167_;
wire _10168_;
wire _10169_;
wire _10170_;
wire _10171_;
wire _10172_;
wire _10173_;
wire _10174_;
wire _10175_;
wire _10176_;
wire _10177_;
wire _10178_;
wire _10179_;
wire _10180_;
wire _10181_;
wire _10182_;
wire _10183_;
wire _10184_;
wire _10185_;
wire _10186_;
wire _10187_;
wire _10188_;
wire _10189_;
wire _10190_;
wire _10191_;
wire _10192_;
wire _10193_;
wire _10194_;
wire _10195_;
wire _10196_;
wire _10197_;
wire _10198_;
wire _10199_;
wire _10200_;
wire _10201_;
wire _10202_;
wire _10203_;
wire _10204_;
wire _10205_;
wire _10206_;
wire _10207_;
wire _10208_;
wire _10209_;
wire _10210_;
wire _10211_;
wire _10212_;
wire _10213_;
wire _10214_;
wire _10215_;
wire _10216_;
wire _10217_;
wire _10218_;
wire _10219_;
wire _10220_;
wire _10221_;
wire _10222_;
wire _10223_;
wire _10224_;
wire _10225_;
wire _10226_;
wire _10227_;
wire _10228_;
wire _10229_;
wire _10230_;
wire _10231_;
wire _10232_;
wire _10233_;
wire _10234_;
wire _10235_;
wire _10236_;
wire _10237_;
wire _10238_;
wire _10239_;
wire _10240_;
wire _10241_;
wire _10242_;
wire _10243_;
wire _10244_;
wire _10245_;
wire _10246_;
wire _10247_;
wire _10248_;
wire _10249_;
wire _10250_;
wire _10251_;
wire _10252_;
wire _10253_;
wire _10254_;
wire _10255_;
wire _10256_;
wire _10257_;
wire _10258_;
wire _10259_;
wire _10260_;
wire _10261_;
wire _10262_;
wire _10263_;
wire _10264_;
wire _10265_;
wire _10266_;
wire _10267_;
wire _10268_;
wire _10269_;
wire _10270_;
wire _10271_;
wire _10272_;
wire _10273_;
wire _10274_;
wire _10275_;
wire _10276_;
wire _10277_;
wire _10278_;
wire _10279_;
wire _10280_;
wire _10281_;
wire _10282_;
wire _10283_;
wire _10284_;
wire _10285_;
wire _10286_;
wire _10287_;
wire _10288_;
wire _10289_;
wire _10290_;
wire _10291_;
wire _10292_;
wire _10293_;
wire _10294_;
wire _10295_;
wire _10296_;
wire _10297_;
wire _10298_;
wire _10299_;
wire _10300_;
wire _10301_;
wire _10302_;
wire _10303_;
wire _10304_;
wire _10305_;
wire _10306_;
wire _10307_;
wire _10308_;
wire _10309_;
wire _10310_;
wire _10311_;
wire _10312_;
wire _10313_;
wire _10314_;
wire _10315_;
wire _10316_;
wire _10317_;
wire _10318_;
wire _10319_;
wire _10320_;
wire _10321_;
wire _10322_;
wire _10323_;
wire _10324_;
wire _10325_;
wire _10326_;
wire _10327_;
wire _10328_;
wire _10329_;
wire _10330_;
wire _10331_;
wire _10332_;
wire _10333_;
wire _10334_;
wire _10335_;
wire _10336_;
wire _10337_;
wire _10338_;
wire _10339_;
wire _10340_;
wire _10341_;
wire _10342_;
wire _10343_;
wire _10344_;
wire _10345_;
wire _10346_;
wire _10347_;
wire _10348_;
wire _10349_;
wire _10350_;
wire _10351_;
wire _10352_;
wire _10353_;
wire _10354_;
wire _10355_;
wire _10356_;
wire _10357_;
wire _10358_;
wire _10359_;
wire _10360_;
wire _10361_;
wire _10362_;
wire _10363_;
wire _10364_;
wire _10365_;
wire _10366_;
wire _10367_;
wire _10368_;
wire _10369_;
wire _10370_;
wire _10371_;
wire _10372_;
wire _10373_;
wire _10374_;
wire _10375_;
wire _10376_;
wire _10377_;
wire _10378_;
wire _10379_;
wire _10380_;
wire _10381_;
wire _10382_;
wire _10383_;
wire _10384_;
wire _10385_;
wire _10386_;
wire _10387_;
wire _10388_;
wire _10389_;
wire _10390_;
wire _10391_;
wire _10392_;
wire _10393_;
wire _10394_;
wire _10395_;
wire _10396_;
wire _10397_;
wire _10398_;
wire _10399_;
wire _10400_;
wire _10401_;
wire _10402_;
wire _10403_;
wire _10404_;
wire _10405_;
wire _10406_;
wire _10407_;
wire _10408_;
wire _10409_;
wire _10410_;
wire _10411_;
wire _10412_;
wire _10413_;
wire _10414_;
wire _10415_;
wire _10416_;
wire _10417_;
wire _10418_;
wire _10419_;
wire _10420_;
wire _10421_;
wire _10422_;
wire _10423_;
wire _10424_;
wire _10425_;
wire _10426_;
wire _10427_;
wire _10428_;
wire _10429_;
wire _10430_;
wire _10431_;
wire _10432_;
wire _10433_;
wire _10434_;
wire _10435_;
wire _10436_;
wire _10437_;
wire _10438_;
wire _10439_;
wire _10440_;
wire _10441_;
wire _10442_;
wire _10443_;
wire _10444_;
wire _10445_;
wire _10446_;
wire _10447_;
wire _10448_;
wire _10449_;
wire _10450_;
wire _10451_;
wire _10452_;
wire _10453_;
wire _10454_;
wire _10455_;
wire _10456_;
wire _10457_;
wire _10458_;
wire _10459_;
wire _10460_;
wire _10461_;
wire _10462_;
wire _10463_;
wire _10464_;
wire _10465_;
wire _10466_;
wire _10467_;
wire _10468_;
wire _10469_;
wire _10470_;
wire _10471_;
wire _10472_;
wire _10473_;
wire _10474_;
wire _10475_;
wire _10476_;
wire _10477_;
wire _10478_;
wire _10479_;
wire _10480_;
wire _10481_;
wire _10482_;
wire _10483_;
wire _10484_;
wire _10485_;
wire _10486_;
wire _10487_;
wire _10488_;
wire _10489_;
wire _10490_;
wire _10491_;
wire _10492_;
wire _10493_;
wire _10494_;
wire _10495_;
wire _10496_;
wire _10497_;
wire _10498_;
wire _10499_;
wire _10500_;
wire _10501_;
wire _10502_;
wire _10503_;
wire _10504_;
wire _10505_;
wire _10506_;
wire _10507_;
wire _10508_;
wire _10509_;
wire _10510_;
wire _10511_;
wire _10512_;
wire _10513_;
wire _10514_;
wire _10515_;
wire _10516_;
wire _10517_;
wire _10518_;
wire _10519_;
wire _10520_;
wire _10521_;
wire _10522_;
wire _10523_;
wire _10524_;
wire _10525_;
wire _10526_;
wire _10527_;
wire _10528_;
wire _10529_;
wire _10530_;
wire _10531_;
wire _10532_;
wire _10533_;
wire _10534_;
wire _10535_;
wire _10536_;
wire _10537_;
wire _10538_;
wire _10539_;
wire _10540_;
wire _10541_;
wire _10542_;
wire _10543_;
wire _10544_;
wire _10545_;
wire _10546_;
wire _10547_;
wire _10548_;
wire _10549_;
wire _10550_;
wire _10551_;
wire _10552_;
wire _10553_;
wire _10554_;
wire _10555_;
wire _10556_;
wire _10557_;
wire _10558_;
wire _10559_;
wire _10560_;
wire _10561_;
wire _10562_;
wire _10563_;
wire _10564_;
wire _10565_;
wire _10566_;
wire _10567_;
wire _10568_;
wire _10569_;
wire _10570_;
wire _10571_;
wire _10572_;
wire _10573_;
wire _10574_;
wire _10575_;
wire _10576_;
wire _10577_;
wire _10578_;
wire _10579_;
wire _10580_;
wire _10581_;
wire _10582_;
wire _10583_;
wire _10584_;
wire _10585_;
wire _10586_;
wire _10587_;
wire _10588_;
wire _10589_;
wire _10590_;
wire _10591_;
wire _10592_;
wire _10593_;
wire _10594_;
wire _10595_;
wire _10596_;
wire _10597_;
wire _10598_;
wire _10599_;
wire _10600_;
wire _10601_;
wire _10602_;
wire _10603_;
wire _10604_;
wire _10605_;
wire _10606_;
wire _10607_;
wire _10608_;
wire _10609_;
wire _10610_;
wire _10611_;
wire _10612_;
wire _10613_;
wire _10614_;
wire _10615_;
wire _10616_;
wire _10617_;
wire _10618_;
wire _10619_;
wire _10620_;
wire _10621_;
wire _10622_;
wire _10623_;
wire _10624_;
wire _10625_;
wire _10626_;
wire _10627_;
wire _10628_;
wire _10629_;
wire _10630_;
wire _10631_;
wire _10632_;
wire _10633_;
wire _10634_;
wire _10635_;
wire _10636_;
wire _10637_;
wire _10638_;
wire _10639_;
wire _10640_;
wire _10641_;
wire _10642_;
wire _10643_;
wire _10644_;
wire _10645_;
wire _10646_;
wire _10647_;
wire _10648_;
wire _10649_;
wire _10650_;
wire _10651_;
wire _10652_;
wire _10653_;
wire _10654_;
wire _10655_;
wire _10656_;
wire _10657_;
wire _10658_;
wire _10659_;
wire _10660_;
wire _10661_;
wire _10662_;
wire _10663_;
wire _10664_;
wire _10665_;
wire _10666_;
wire _10667_;
wire _10668_;
wire _10669_;
wire _10670_;
wire _10671_;
wire _10672_;
wire _10673_;
wire _10674_;
wire _10675_;
wire _10676_;
wire _10677_;
wire _10678_;
wire _10679_;
wire _10680_;
wire _10681_;
wire _10682_;
wire _10683_;
wire _10684_;
wire _10685_;
wire _10686_;
wire _10687_;
wire _10688_;
wire _10689_;
wire _10690_;
wire _10691_;
wire _10692_;
wire _10693_;
wire _10694_;
wire _10695_;
wire _10696_;
wire _10697_;
wire _10698_;
wire _10699_;
wire _10700_;
wire _10701_;
wire _10702_;
wire _10703_;
wire _10704_;
wire _10705_;
wire _10706_;
wire _10707_;
wire _10708_;
wire _10709_;
wire _10710_;
wire _10711_;
wire _10712_;
wire _10713_;
wire _10714_;
wire _10715_;
wire _10716_;
wire _10717_;
wire _10718_;
wire _10719_;
wire _10720_;
wire _10721_;
wire _10722_;
wire _10723_;
wire _10724_;
wire _10725_;
wire _10726_;
wire _10727_;
wire _10728_;
wire _10729_;
wire _10730_;
wire _10731_;
wire _10732_;
wire _10733_;
wire _10734_;
wire _10735_;
wire _10736_;
wire _10737_;
wire _10738_;
wire _10739_;
wire _10740_;
wire _10741_;
wire _10742_;
wire _10743_;
wire _10744_;
wire _10745_;
wire _10746_;
wire _10747_;
wire _10748_;
wire _10749_;
wire _10750_;
wire _10751_;
wire _10752_;
wire _10753_;
wire _10754_;
wire _10755_;
wire _10756_;
wire _10757_;
wire _10758_;
wire _10759_;
wire _10760_;
wire _10761_;
wire _10762_;
wire _10763_;
wire _10764_;
wire _10765_;
wire _10766_;
wire _10767_;
wire _10768_;
wire _10769_;
wire _10770_;
wire _10771_;
wire _10772_;
wire _10773_;
wire _10774_;
wire _10775_;
wire _10776_;
wire _10777_;
wire _10778_;
wire _10779_;
wire _10780_;
wire _10781_;
wire _10782_;
wire _10783_;
wire _10784_;
wire _10785_;
wire _10786_;
wire _10787_;
wire _10788_;
wire _10789_;
wire _10790_;
wire _10791_;
wire _10792_;
wire _10793_;
wire _10794_;
wire _10795_;
wire _10796_;
wire _10797_;
wire _10798_;
wire _10799_;
wire _10800_;
wire _10801_;
wire _10802_;
wire _10803_;
wire _10804_;
wire _10805_;
wire _10806_;
wire _10807_;
wire _10808_;
wire _10809_;
wire _10810_;
wire _10811_;
wire _10812_;
wire _10813_;
wire _10814_;
wire _10815_;
wire _10816_;
wire _10817_;
wire _10818_;
wire _10819_;
wire _10820_;
wire _10821_;
wire _10822_;
wire _10823_;
wire _10824_;
wire _10825_;
wire _10826_;
wire _10827_;
wire _10828_;
wire _10829_;
wire _10830_;
wire _10831_;
wire _10832_;
wire _10833_;
wire _10834_;
wire _10835_;
wire _10836_;
wire _10837_;
wire _10838_;
wire _10839_;
wire _10840_;
wire _10841_;
wire _10842_;
wire _10843_;
wire _10844_;
wire _10845_;
wire _10846_;
wire _10847_;
wire _10848_;
wire _10849_;
wire _10850_;
wire _10851_;
wire _10852_;
wire _10853_;
wire _10854_;
wire _10855_;
wire _10856_;
wire _10857_;
wire _10858_;
wire _10859_;
wire _10860_;
wire _10861_;
wire _10862_;
wire _10863_;
wire _10864_;
wire _10865_;
wire _10866_;
wire _10867_;
wire _10868_;
wire _10869_;
wire _10870_;
wire _10871_;
wire _10872_;
wire _10873_;
wire _10874_;
wire _10875_;
wire _10876_;
wire _10877_;
wire _10878_;
wire _10879_;
wire _10880_;
wire _10881_;
wire _10882_;
wire _10883_;
wire _10884_;
wire _10885_;
wire _10886_;
wire _10887_;
wire _10888_;
wire _10889_;
wire _10890_;
wire _10891_;
wire _10892_;
wire _10893_;
wire _10894_;
wire _10895_;
wire _10896_;
wire _10897_;
wire _10898_;
wire _10899_;
wire _10900_;
wire _10901_;
wire _10902_;
wire _10903_;
wire _10904_;
wire _10905_;
wire _10906_;
wire _10907_;
wire _10908_;
wire _10909_;
wire _10910_;
wire _10911_;
wire _10912_;
wire _10913_;
wire _10914_;
wire _10915_;
wire _10916_;
wire _10917_;
wire _10918_;
wire _10919_;
wire _10920_;
wire _10921_;
wire _10922_;
wire _10923_;
wire _10924_;
wire _10925_;
wire _10926_;
wire _10927_;
wire _10928_;
wire _10929_;
wire _10930_;
wire _10931_;
wire _10932_;
wire _10933_;
wire _10934_;
wire _10935_;
wire _10936_;
wire _10937_;
wire _10938_;
wire _10939_;
wire _10940_;
wire _10941_;
wire _10942_;
wire _10943_;
wire _10944_;
wire _10945_;
wire _10946_;
wire _10947_;
wire _10948_;
wire _10949_;
wire _10950_;
wire _10951_;
wire _10952_;
wire _10953_;
wire _10954_;
wire _10955_;
wire _10956_;
wire _10957_;
wire _10958_;
wire _10959_;
wire _10960_;
wire _10961_;
wire _10962_;
wire _10963_;
wire _10964_;
wire _10965_;
wire _10966_;
wire _10967_;
wire _10968_;
wire _10969_;
wire _10970_;
wire _10971_;
wire _10972_;
wire _10973_;
wire _10974_;
wire _10975_;
wire _10976_;
wire _10977_;
wire _10978_;
wire _10979_;
wire _10980_;
wire _10981_;
wire _10982_;
wire _10983_;
wire _10984_;
wire _10985_;
wire _10986_;
wire _10987_;
wire _10988_;
wire _10989_;
wire _10990_;
wire _10991_;
wire _10992_;
wire _10993_;
wire _10994_;
wire _10995_;
wire _10996_;
wire _10997_;
wire _10998_;
wire _10999_;
wire _11000_;
wire _11001_;
wire _11002_;
wire _11003_;
wire _11004_;
wire _11005_;
wire _11006_;
wire _11007_;
wire _11008_;
wire _11009_;
wire _11010_;
wire _11011_;
wire _11012_;
wire _11013_;
wire _11014_;
wire _11015_;
wire _11016_;
wire _11017_;
wire _11018_;
wire _11019_;
wire _11020_;
wire _11021_;
wire _11022_;
wire _11023_;
wire _11024_;
wire _11025_;
wire _11026_;
wire _11027_;
wire _11028_;
wire _11029_;
wire _11030_;
wire _11031_;
wire _11032_;
wire _11033_;
wire _11034_;
wire _11035_;
wire _11036_;
wire _11037_;
wire _11038_;
wire _11039_;
wire _11040_;
wire _11041_;
wire _11042_;
wire _11043_;
wire _11044_;
wire _11045_;
wire _11046_;
wire _11047_;
wire _11048_;
wire _11049_;
wire _11050_;
wire _11051_;
wire _11052_;
wire _11053_;
wire _11054_;
wire _11055_;
wire _11056_;
wire _11057_;
wire _11058_;
wire _11059_;
wire _11060_;
wire _11061_;
wire _11062_;
wire _11063_;
wire _11064_;
wire _11065_;
wire _11066_;
wire _11067_;
wire _11068_;
wire _11069_;
wire _11070_;
wire _11071_;
wire _11072_;
wire _11073_;
wire _11074_;
wire _11075_;
wire _11076_;
wire _11077_;
wire _11078_;
wire _11079_;
wire _11080_;
wire _11081_;
wire _11082_;
wire _11083_;
wire _11084_;
wire _11085_;
wire _11086_;
wire _11087_;
wire _11088_;
wire _11089_;
wire _11090_;
wire _11091_;
wire _11092_;
wire _11093_;
wire _11094_;
wire _11095_;
wire _11096_;
wire _11097_;
wire _11098_;
wire _11099_;
wire _11100_;
wire _11101_;
wire _11102_;
wire _11103_;
wire _11104_;
wire _11105_;
wire _11106_;
wire _11107_;
wire _11108_;
wire _11109_;
wire _11110_;
wire _11111_;
wire _11112_;
wire _11113_;
wire _11114_;
wire _11115_;
wire _11116_;
wire _11117_;
wire _11118_;
wire _11119_;
wire _11120_;
wire _11121_;
wire _11122_;
wire _11123_;
wire _11124_;
wire _11125_;
wire _11126_;
wire _11127_;
wire _11128_;
wire _11129_;
wire _11130_;
wire _11131_;
wire _11132_;
wire _11133_;
wire _11134_;
wire _11135_;
wire _11136_;
wire _11137_;
wire _11138_;
wire _11139_;
wire _11140_;
wire _11141_;
wire _11142_;
wire _11143_;
wire _11144_;
wire _11145_;
wire _11146_;
wire _11147_;
wire _11148_;
wire _11149_;
wire _11150_;
wire _11151_;
wire _11152_;
wire _11153_;
wire _11154_;
wire _11155_;
wire _11156_;
wire _11157_;
wire _11158_;
wire _11159_;
wire _11160_;
wire _11161_;
wire _11162_;
wire _11163_;
wire _11164_;
wire _11165_;
wire _11166_;
wire _11167_;
wire _11168_;
wire _11169_;
wire _11170_;
wire _11171_;
wire _11172_;
wire _11173_;
wire _11174_;
wire _11175_;
wire _11176_;
wire _11177_;
wire _11178_;
wire _11179_;
wire _11180_;
wire _11181_;
wire _11182_;
wire _11183_;
wire _11184_;
wire _11185_;
wire _11186_;
wire _11187_;
wire _11188_;
wire _11189_;
wire _11190_;
wire _11191_;
wire _11192_;
wire _11193_;
wire _11194_;
wire _11195_;
wire _11196_;
wire _11197_;
wire _11198_;
wire _11199_;
wire _11200_;
wire _11201_;
wire _11202_;
wire _11203_;
wire _11204_;
wire _11205_;
wire _11206_;
wire _11207_;
wire _11208_;
wire _11209_;
wire _11210_;
wire _11211_;
wire _11212_;
wire _11213_;
wire _11214_;
wire _11215_;
wire _11216_;
wire _11217_;
wire _11218_;
wire _11219_;
wire _11220_;
wire _11221_;
wire _11222_;
wire _11223_;
wire _11224_;
wire _11225_;
wire _11226_;
wire _11227_;
wire _11228_;
wire _11229_;
wire _11230_;
wire _11231_;
wire _11232_;
wire _11233_;
wire _11234_;
wire _11235_;
wire _11236_;
wire _11237_;
wire _11238_;
wire _11239_;
wire _11240_;
wire _11241_;
wire _11242_;
wire _11243_;
wire _11244_;
wire _11245_;
wire _11246_;
wire _11247_;
wire _11248_;
wire _11249_;
wire _11250_;
wire _11251_;
wire _11252_;
wire _11253_;
wire _11254_;
wire _11255_;
wire _11256_;
wire _11257_;
wire _11258_;
wire _11259_;
wire _11260_;
wire _11261_;
wire _11262_;
wire _11263_;
wire _11264_;
wire _11265_;
wire _11266_;
wire _11267_;
wire _11268_;
wire _11269_;
wire _11270_;
wire _11271_;
wire _11272_;
wire _11273_;
wire _11274_;
wire _11275_;
wire _11276_;
wire _11277_;
wire _11278_;
wire _11279_;
wire _11280_;
wire _11281_;
wire _11282_;
wire _11283_;
wire _11284_;
wire _11285_;
wire _11286_;
wire _11287_;
wire _11288_;
wire _11289_;
wire _11290_;
wire _11291_;
wire _11292_;
wire _11293_;
wire _11294_;
wire _11295_;
wire _11296_;
wire _11297_;
wire _11298_;
wire _11299_;
wire _11300_;
wire _11301_;
wire _11302_;
wire _11303_;
wire _11304_;
wire _11305_;
wire _11306_;
wire _11307_;
wire _11308_;
wire _11309_;
wire _11310_;
wire _11311_;
wire _11312_;
wire _11313_;
wire _11314_;
wire _11315_;
wire _11316_;
wire _11317_;
wire _11318_;
wire _11319_;
wire _11320_;
wire _11321_;
wire _11322_;
wire _11323_;
wire _11324_;
wire _11325_;
wire _11326_;
wire _11327_;
wire _11328_;
wire _11329_;
wire _11330_;
wire _11331_;
wire _11332_;
wire _11333_;
wire _11334_;
wire _11335_;
wire _11336_;
wire _11337_;
wire _11338_;
wire _11339_;
wire _11340_;
wire _11341_;
wire _11342_;
wire _11343_;
wire _11344_;
wire _11345_;
wire _11346_;
wire _11347_;
wire _11348_;
wire _11349_;
wire _11350_;
wire _11351_;
wire _11352_;
wire _11353_;
wire _11354_;
wire _11355_;
wire _11356_;
wire _11357_;
wire _11358_;
wire _11359_;
wire _11360_;
wire _11361_;
wire _11362_;
wire _11363_;
wire _11364_;
wire _11365_;
wire _11366_;
wire _11367_;
wire _11368_;
wire _11369_;
wire _11370_;
wire _11371_;
wire _11372_;
wire _11373_;
wire _11374_;
wire _11375_;
wire _11376_;
wire _11377_;
wire _11378_;
wire _11379_;
wire _11380_;
wire _11381_;
wire _11382_;
wire _11383_;
wire _11384_;
wire _11385_;
wire _11386_;
wire _11387_;
wire _11388_;
wire _11389_;
wire _11390_;
wire _11391_;
wire _11392_;
wire _11393_;
wire _11394_;
wire _11395_;
wire _11396_;
wire _11397_;
wire _11398_;
wire _11399_;
wire _11400_;
wire _11401_;
wire _11402_;
wire _11403_;
wire _11404_;
wire _11405_;
wire _11406_;
wire _11407_;
wire _11408_;
wire _11409_;
wire _11410_;
wire _11411_;
wire _11412_;
wire _11413_;
wire _11414_;
wire _11415_;
wire _11416_;
wire _11417_;
wire _11418_;
wire _11419_;
wire _11420_;
wire _11421_;
wire _11422_;
wire _11423_;
wire _11424_;
wire _11425_;
wire _11426_;
wire _11427_;
wire _11428_;
wire _11429_;
wire _11430_;
wire _11431_;
wire _11432_;
wire _11433_;
wire _11434_;
wire _11435_;
wire _11436_;
wire _11437_;
wire _11438_;
wire _11439_;
wire _11440_;
wire _11441_;
wire _11442_;
wire _11443_;
wire _11444_;
wire _11445_;
wire _11446_;
wire _11447_;
wire _11448_;
wire _11449_;
wire _11450_;
wire _11451_;
wire _11452_;
wire _11453_;
wire _11454_;
wire _11455_;
wire _11456_;
wire _11457_;
wire _11458_;
wire _11459_;
wire _11460_;
wire _11461_;
wire _11462_;
wire _11463_;
wire _11464_;
wire _11465_;
wire _11466_;
wire _11467_;
wire _11468_;
wire _11469_;
wire _11470_;
wire _11471_;
wire _11472_;
wire _11473_;
wire _11474_;
wire _11475_;
wire _11476_;
wire _11477_;
wire _11478_;
wire _11479_;
wire _11480_;
wire _11481_;
wire _11482_;
wire _11483_;
wire _11484_;
wire _11485_;
wire _11486_;
wire _11487_;
wire _11488_;
wire _11489_;
wire _11490_;
wire _11491_;
wire _11492_;
wire _11493_;
wire _11494_;
wire _11495_;
wire _11496_;
wire _11497_;
wire _11498_;
wire _11499_;
wire _11500_;
wire _11501_;
wire _11502_;
wire _11503_;
wire _11504_;
wire _11505_;
wire _11506_;
wire _11507_;
wire _11508_;
wire _11509_;
wire _11510_;
wire _11511_;
wire _11512_;
wire _11513_;
wire _11514_;
wire _11515_;
wire _11516_;
wire _11517_;
wire _11518_;
wire _11519_;
wire _11520_;
wire _11521_;
wire _11522_;
wire _11523_;
wire _11524_;
wire _11525_;
wire _11526_;
wire _11527_;
wire _11528_;
wire _11529_;
wire _11530_;
wire _11531_;
wire _11532_;
wire _11533_;
wire _11534_;
wire _11535_;
wire _11536_;
wire _11537_;
wire _11538_;
wire _11539_;
wire _11540_;
wire _11541_;
wire _11542_;
wire _11543_;
wire _11544_;
wire _11545_;
wire _11546_;
wire _11547_;
wire _11548_;
wire _11549_;
wire _11550_;
wire _11551_;
wire _11552_;
wire _11553_;
wire _11554_;
wire _11555_;
wire _11556_;
wire _11557_;
wire _11558_;
wire _11559_;
wire _11560_;
wire _11561_;
wire _11562_;
wire _11563_;
wire _11564_;
wire _11565_;
wire _11566_;
wire _11567_;
wire _11568_;
wire _11569_;
wire _11570_;
wire _11571_;
wire _11572_;
wire _11573_;
wire _11574_;
wire _11575_;
wire _11576_;
wire _11577_;
wire _11578_;
wire _11579_;
wire _11580_;
wire _11581_;
wire _11582_;
wire _11583_;
wire _11584_;
wire _11585_;
wire _11586_;
wire _11587_;
wire _11588_;
wire _11589_;
wire _11590_;
wire _11591_;
wire _11592_;
wire _11593_;
wire _11594_;
wire _11595_;
wire _11596_;
wire _11597_;
wire _11598_;
wire _11599_;
wire _11600_;
wire _11601_;
wire _11602_;
wire _11603_;
wire _11604_;
wire _11605_;
wire _11606_;
wire _11607_;
wire _11608_;
wire _11609_;
wire _11610_;
wire _11611_;
wire _11612_;
wire _11613_;
wire _11614_;
wire _11615_;
wire _11616_;
wire _11617_;
wire _11618_;
wire _11619_;
wire _11620_;
wire _11621_;
wire _11622_;
wire _11623_;
wire _11624_;
wire _11625_;
wire _11626_;
wire _11627_;
wire _11628_;
wire _11629_;
wire _11630_;
wire _11631_;
wire _11632_;
wire _11633_;
wire _11634_;
wire _11635_;
wire _11636_;
wire _11637_;
wire _11638_;
wire _11639_;
wire _11640_;
wire _11641_;
wire _11642_;
wire _11643_;
wire _11644_;
wire _11645_;
wire _11646_;
wire _11647_;
wire _11648_;
wire _11649_;
wire _11650_;
wire _11651_;
wire _11652_;
wire _11653_;
wire _11654_;
wire _11655_;
wire _11656_;
wire _11657_;
wire _11658_;
wire _11659_;
wire _11660_;
wire _11661_;
wire _11662_;
wire _11663_;
wire _11664_;
wire _11665_;
wire _11666_;
wire _11667_;
wire _11668_;
wire _11669_;
wire _11670_;
wire _11671_;
wire _11672_;
wire _11673_;
wire _11674_;
wire _11675_;
wire _11676_;
wire _11677_;
wire _11678_;
wire _11679_;
wire _11680_;
wire _11681_;
wire _11682_;
wire _11683_;
wire _11684_;
wire _11685_;
wire _11686_;
wire _11687_;
wire _11688_;
wire _11689_;
wire _11690_;
wire _11691_;
wire _11692_;
wire _11693_;
wire _11694_;
wire _11695_;
wire _11696_;
wire _11697_;
wire _11698_;
wire _11699_;
wire _11700_;
wire _11701_;
wire _11702_;
wire _11703_;
wire _11704_;
wire _11705_;
wire _11706_;
wire _11707_;
wire _11708_;
wire _11709_;
wire _11710_;
wire _11711_;
wire _11712_;
wire _11713_;
wire _11714_;
wire _11715_;
wire _11716_;
wire _11717_;
wire _11718_;
wire _11719_;
wire _11720_;
wire _11721_;
wire _11722_;
wire _11723_;
wire _11724_;
wire _11725_;
wire _11726_;
wire _11727_;
wire _11728_;
wire _11729_;
wire _11730_;
wire _11731_;
wire _11732_;
wire _11733_;
wire _11734_;
wire _11735_;
wire _11736_;
wire _11737_;
wire _11738_;
wire _11739_;
wire _11740_;
wire _11741_;
wire _11742_;
wire _11743_;
wire _11744_;
wire _11745_;
wire _11746_;
wire _11747_;
wire _11748_;
wire _11749_;
wire _11750_;
wire _11751_;
wire _11752_;
wire _11753_;
wire _11754_;
wire _11755_;
wire _11756_;
wire _11757_;
wire _11758_;
wire _11759_;
wire _11760_;
wire _11761_;
wire _11762_;
wire _11763_;
wire _11764_;
wire _11765_;
wire _11766_;
wire _11767_;
wire _11768_;
wire _11769_;
wire _11770_;
wire _11771_;
wire _11772_;
wire _11773_;
wire _11774_;
wire _11775_;
wire _11776_;
wire _11777_;
wire _11778_;
wire _11779_;
wire _11780_;
wire _11781_;
wire _11782_;
wire _11783_;
wire _11784_;
wire _11785_;
wire _11786_;
wire _11787_;
wire _11788_;
wire _11789_;
wire _11790_;
wire _11791_;
wire _11792_;
wire _11793_;
wire _11794_;
wire _11795_;
wire _11796_;
wire _11797_;
wire _11798_;
wire _11799_;
wire _11800_;
wire _11801_;
wire _11802_;
wire _11803_;
wire _11804_;
wire _11805_;
wire _11806_;
wire _11807_;
wire _11808_;
wire _11809_;
wire _11810_;
wire _11811_;
wire _11812_;
wire _11813_;
wire _11814_;
wire _11815_;
wire _11816_;
wire _11817_;
wire _11818_;
wire _11819_;
wire _11820_;
wire _11821_;
wire _11822_;
wire _11823_;
wire _11824_;
wire _11825_;
wire _11826_;
wire _11827_;
wire _11828_;
wire _11829_;
wire _11830_;
wire _11831_;
wire _11832_;
wire _11833_;
wire _11834_;
wire _11835_;
wire _11836_;
wire _11837_;
wire _11838_;
wire _11839_;
wire _11840_;
wire _11841_;
wire _11842_;
wire _11843_;
wire _11844_;
wire _11845_;
wire _11846_;
wire _11847_;
wire _11848_;
wire _11849_;
wire _11850_;
wire _11851_;
wire _11852_;
wire _11853_;
wire _11854_;
wire _11855_;
wire _11856_;
wire _11857_;
wire _11858_;
wire _11859_;
wire _11860_;
wire _11861_;
wire _11862_;
wire _11863_;
wire _11864_;
wire _11865_;
wire _11866_;
wire _11867_;
wire _11868_;
wire _11869_;
wire _11870_;
wire _11871_;
wire _11872_;
wire _11873_;
wire _11874_;
wire _11875_;
wire _11876_;
wire _11877_;
wire _11878_;
wire _11879_;
wire _11880_;
wire _11881_;
wire _11882_;
wire _11883_;
wire _11884_;
wire _11885_;
wire _11886_;
wire _11887_;
wire _11888_;
wire _11889_;
wire _11890_;
wire _11891_;
wire _11892_;
wire _11893_;
wire _11894_;
wire _11895_;
wire _11896_;
wire _11897_;
wire _11898_;
wire _11899_;
wire _11900_;
wire _11901_;
wire _11902_;
wire _11903_;
wire _11904_;
wire _11905_;
wire _11906_;
wire _11907_;
wire _11908_;
wire _11909_;
wire _11910_;
wire _11911_;
wire _11912_;
wire _11913_;
wire _11914_;
wire _11915_;
wire _11916_;
wire _11917_;
wire _11918_;
wire _11919_;
wire _11920_;
wire _11921_;
wire _11922_;
wire _11923_;
wire _11924_;
wire _11925_;
wire _11926_;
wire _11927_;
wire _11928_;
wire _11929_;
wire _11930_;
wire _11931_;
wire _11932_;
wire _11933_;
wire _11934_;
wire _11935_;
wire _11936_;
wire _11937_;
wire _11938_;
wire _11939_;
wire _11940_;
wire _11941_;
wire _11942_;
wire _11943_;
wire _11944_;
wire _11945_;
wire _11946_;
wire _11947_;
wire _11948_;
wire _11949_;
wire _11950_;
wire _11951_;
wire _11952_;
wire _11953_;
wire _11954_;
wire _11955_;
wire _11956_;
wire _11957_;
wire _11958_;
wire _11959_;
wire _11960_;
wire _11961_;
wire _11962_;
wire _11963_;
wire _11964_;
wire _11965_;
wire _11966_;
wire _11967_;
wire _11968_;
wire _11969_;
wire _11970_;
wire _11971_;
wire _11972_;
wire _11973_;
wire _11974_;
wire _11975_;
wire _11976_;
wire _11977_;
wire _11978_;
wire _11979_;
wire _11980_;
wire _11981_;
wire _11982_;
wire _11983_;
wire _11984_;
wire _11985_;
wire _11986_;
wire _11987_;
wire _11988_;
wire _11989_;
wire _11990_;
wire _11991_;
wire _11992_;
wire _11993_;
wire _11994_;
wire _11995_;
wire _11996_;
wire _11997_;
wire _11998_;
wire _11999_;
wire _12000_;
wire _12001_;
wire _12002_;
wire _12003_;
wire _12004_;
wire _12005_;
wire _12006_;
wire _12007_;
wire _12008_;
wire _12009_;
wire _12010_;
wire _12011_;
wire _12012_;
wire _12013_;
wire _12014_;
wire _12015_;
wire _12016_;
wire _12017_;
wire _12018_;
wire _12019_;
wire _12020_;
wire _12021_;
wire _12022_;
wire _12023_;
wire _12024_;
wire _12025_;
wire _12026_;
wire _12027_;
wire _12028_;
wire _12029_;
wire _12030_;
wire _12031_;
wire _12032_;
wire _12033_;
wire _12034_;
wire _12035_;
wire _12036_;
wire _12037_;
wire _12038_;
wire _12039_;
wire _12040_;
wire _12041_;
wire _12042_;
wire _12043_;
wire _12044_;
wire _12045_;
wire _12046_;
wire _12047_;
wire _12048_;
wire _12049_;
wire _12050_;
wire _12051_;
wire _12052_;
wire _12053_;
wire _12054_;
wire _12055_;
wire _12056_;
wire _12057_;
wire _12058_;
wire _12059_;
wire _12060_;
wire _12061_;
wire _12062_;
wire _12063_;
wire _12064_;
wire _12065_;
wire _12066_;
wire _12067_;
wire _12068_;
wire _12069_;
wire _12070_;
wire _12071_;
wire _12072_;
wire _12073_;
wire _12074_;
wire _12075_;
wire _12076_;
wire _12077_;
wire _12078_;
wire _12079_;
wire _12080_;
wire _12081_;
wire _12082_;
wire _12083_;
wire _12084_;
wire _12085_;
wire _12086_;
wire _12087_;
wire _12088_;
wire _12089_;
wire _12090_;
wire _12091_;
wire _12092_;
wire _12093_;
wire _12094_;
wire _12095_;
wire _12096_;
wire _12097_;
wire _12098_;
wire _12099_;
wire _12100_;
wire _12101_;
wire _12102_;
wire _12103_;
wire _12104_;
wire _12105_;
wire _12106_;
wire _12107_;
wire _12108_;
wire _12109_;
wire _12110_;
wire _12111_;
wire _12112_;
wire _12113_;
wire _12114_;
wire _12115_;
wire _12116_;
wire _12117_;
wire _12118_;
wire _12119_;
wire _12120_;
wire _12121_;
wire _12122_;
wire _12123_;
wire _12124_;
wire _12125_;
wire _12126_;
wire _12127_;
wire _12128_;
wire _12129_;
wire _12130_;
wire _12131_;
wire _12132_;
wire _12133_;
wire _12134_;
wire _12135_;
wire _12136_;
wire _12137_;
wire _12138_;
wire _12139_;
wire _12140_;
wire _12141_;
wire _12142_;
wire _12143_;
wire _12144_;
wire _12145_;
wire _12146_;
wire _12147_;
wire _12148_;
wire _12149_;
wire _12150_;
wire _12151_;
wire _12152_;
wire _12153_;
wire _12154_;
wire _12155_;
wire _12156_;
wire _12157_;
wire _12158_;
wire _12159_;
wire _12160_;
wire _12161_;
wire _12162_;
wire _12163_;
wire _12164_;
wire _12165_;
wire _12166_;
wire _12167_;
wire _12168_;
wire _12169_;
wire _12170_;
wire _12171_;
wire _12172_;
wire _12173_;
wire _12174_;
wire _12175_;
wire _12176_;
wire _12177_;
wire _12178_;
wire _12179_;
wire _12180_;
wire _12181_;
wire _12182_;
wire _12183_;
wire _12184_;
wire _12185_;
wire _12186_;
wire _12187_;
wire _12188_;
wire _12189_;
wire _12190_;
wire _12191_;
wire _12192_;
wire _12193_;
wire _12194_;
wire _12195_;
wire _12196_;
wire _12197_;
wire _12198_;
wire _12199_;
wire _12200_;
wire _12201_;
wire _12202_;
wire _12203_;
wire _12204_;
wire _12205_;
wire _12206_;
wire _12207_;
wire _12208_;
wire _12209_;
wire _12210_;
wire _12211_;
wire _12212_;
wire _12213_;
wire _12214_;
wire _12215_;
wire _12216_;
wire _12217_;
wire _12218_;
wire _12219_;
wire _12220_;
wire _12221_;
wire _12222_;
wire _12223_;
wire _12224_;
wire _12225_;
wire _12226_;
wire _12227_;
wire _12228_;
wire _12229_;
wire _12230_;
wire _12231_;
wire _12232_;
wire _12233_;
wire _12234_;
wire _12235_;
wire _12236_;
wire _12237_;
wire _12238_;
wire _12239_;
wire _12240_;
wire _12241_;
wire _12242_;
wire _12243_;
wire _12244_;
wire _12245_;
wire _12246_;
wire _12247_;
wire _12248_;
wire _12249_;
wire _12250_;
wire _12251_;
wire _12252_;
wire _12253_;
wire _12254_;
wire _12255_;
wire _12256_;
wire _12257_;
wire _12258_;
wire _12259_;
wire _12260_;
wire _12261_;
wire _12262_;
wire _12263_;
wire _12264_;
wire _12265_;
wire _12266_;
wire _12267_;
wire _12268_;
wire _12269_;
wire _12270_;
wire _12271_;
wire _12272_;
wire _12273_;
wire _12274_;
wire _12275_;
wire _12276_;
wire _12277_;
wire _12278_;
wire _12279_;
wire _12280_;
wire _12281_;
wire _12282_;
wire _12283_;
wire _12284_;
wire _12285_;
wire _12286_;
wire _12287_;
wire _12288_;
wire _12289_;
wire _12290_;
wire _12291_;
wire _12292_;
wire _12293_;
wire _12294_;
wire _12295_;
wire _12296_;
wire _12297_;
wire _12298_;
wire _12299_;
wire _12300_;
wire _12301_;
wire _12302_;
wire _12303_;
wire _12304_;
wire _12305_;
wire _12306_;
wire _12307_;
wire _12308_;
wire _12309_;
wire _12310_;
wire _12311_;
wire _12312_;
wire _12313_;
wire _12314_;
wire _12315_;
wire _12316_;
wire _12317_;
wire _12318_;
wire _12319_;
wire _12320_;
wire _12321_;
wire _12322_;
wire _12323_;
wire _12324_;
wire _12325_;
wire _12326_;
wire _12327_;
wire _12328_;
wire _12329_;
wire _12330_;
wire _12331_;
wire _12332_;
wire _12333_;
wire _12334_;
wire _12335_;
wire _12336_;
wire _12337_;
wire _12338_;
wire _12339_;
wire _12340_;
wire _12341_;
wire _12342_;
wire _12343_;
wire _12344_;
wire _12345_;
wire _12346_;
wire _12347_;
wire _12348_;
wire _12349_;
wire _12350_;
wire _12351_;
wire _12352_;
wire _12353_;
wire _12354_;
wire _12355_;
wire _12356_;
wire _12357_;
wire _12358_;
wire _12359_;
wire _12360_;
wire _12361_;
wire _12362_;
wire _12363_;
wire _12364_;
wire _12365_;
wire _12366_;
wire _12367_;
wire _12368_;
wire _12369_;
wire _12370_;
wire _12371_;
wire _12372_;
wire _12373_;
wire _12374_;
wire _12375_;
wire _12376_;
wire _12377_;
wire _12378_;
wire _12379_;
wire _12380_;
wire _12381_;
wire _12382_;
wire _12383_;
wire _12384_;
wire _12385_;
wire _12386_;
wire _12387_;
wire _12388_;
wire _12389_;
wire _12390_;
wire _12391_;
wire _12392_;
wire _12393_;
wire _12394_;
wire _12395_;
wire _12396_;
wire _12397_;
wire _12398_;
wire _12399_;
wire _12400_;
wire _12401_;
wire _12402_;
wire _12403_;
wire _12404_;
wire _12405_;
wire _12406_;
wire _12407_;
wire _12408_;
wire _12409_;
wire _12410_;
wire _12411_;
wire _12412_;
wire _12413_;
wire _12414_;
wire _12415_;
wire _12416_;
wire _12417_;
wire _12418_;
wire _12419_;
wire _12420_;
wire _12421_;
wire _12422_;
wire _12423_;
wire _12424_;
wire _12425_;
wire _12426_;
wire _12427_;
wire _12428_;
wire _12429_;
wire _12430_;
wire _12431_;
wire _12432_;
wire _12433_;
wire _12434_;
wire _12435_;
wire _12436_;
wire _12437_;
wire _12438_;
wire _12439_;
wire _12440_;
wire _12441_;
wire _12442_;
wire _12443_;
wire _12444_;
wire _12445_;
wire _12446_;
wire _12447_;
wire _12448_;
wire _12449_;
wire _12450_;
wire _12451_;
wire _12452_;
wire _12453_;
wire _12454_;
wire _12455_;
wire _12456_;
wire _12457_;
wire _12458_;
wire _12459_;
wire _12460_;
wire _12461_;
wire _12462_;
wire _12463_;
wire _12464_;
wire _12465_;
wire _12466_;
wire _12467_;
wire _12468_;
wire _12469_;
wire _12470_;
wire _12471_;
wire _12472_;
wire _12473_;
wire _12474_;
wire _12475_;
wire _12476_;
wire _12477_;
wire _12478_;
wire _12479_;
wire _12480_;
wire _12481_;
wire _12482_;
wire _12483_;
wire _12484_;
wire _12485_;
wire _12486_;
wire _12487_;
wire _12488_;
wire _12489_;
wire _12490_;
wire _12491_;
wire _12492_;
wire _12493_;
wire _12494_;
wire _12495_;
wire _12496_;
wire _12497_;
wire _12498_;
wire _12499_;
wire _12500_;
wire _12501_;
wire _12502_;
wire _12503_;
wire _12504_;
wire _12505_;
wire _12506_;
wire _12507_;
wire _12508_;
wire _12509_;
wire _12510_;
wire _12511_;
wire _12512_;
wire _12513_;
wire _12514_;
wire _12515_;
wire _12516_;
wire _12517_;
wire _12518_;
wire _12519_;
wire _12520_;
wire _12521_;
wire _12522_;
wire _12523_;
wire _12524_;
wire _12525_;
wire _12526_;
wire _12527_;
wire _12528_;
wire _12529_;
wire _12530_;
wire _12531_;
wire _12532_;
wire _12533_;
wire _12534_;
wire _12535_;
wire _12536_;
wire _12537_;
wire _12538_;
wire _12539_;
wire _12540_;
wire _12541_;
wire _12542_;
wire _12543_;
wire _12544_;
wire _12545_;
wire _12546_;
wire _12547_;
wire _12548_;
wire _12549_;
wire _12550_;
wire _12551_;
wire _12552_;
wire _12553_;
wire _12554_;
wire _12555_;
wire _12556_;
wire _12557_;
wire _12558_;
wire _12559_;
wire _12560_;
wire _12561_;
wire _12562_;
wire _12563_;
wire _12564_;
wire _12565_;
wire _12566_;
wire _12567_;
wire _12568_;
wire _12569_;
wire _12570_;
wire _12571_;
wire _12572_;
wire _12573_;
wire _12574_;
wire _12575_;
wire _12576_;
wire _12577_;
wire _12578_;
wire _12579_;
wire _12580_;
wire _12581_;
wire _12582_;
wire _12583_;
wire _12584_;
wire _12585_;
wire _12586_;
wire _12587_;
wire _12588_;
wire _12589_;
wire _12590_;
wire _12591_;
wire _12592_;
wire _12593_;
wire _12594_;
wire _12595_;
wire _12596_;
wire _12597_;
wire _12598_;
wire _12599_;
wire _12600_;
wire _12601_;
wire _12602_;
wire _12603_;
wire _12604_;
wire _12605_;
wire _12606_;
wire _12607_;
wire _12608_;
wire _12609_;
wire _12610_;
wire _12611_;
wire _12612_;
wire _12613_;
wire _12614_;
wire _12615_;
wire _12616_;
wire _12617_;
wire _12618_;
wire _12619_;
wire _12620_;
wire _12621_;
wire _12622_;
wire _12623_;
wire _12624_;
wire _12625_;
wire _12626_;
wire _12627_;
wire _12628_;
wire _12629_;
wire _12630_;
wire _12631_;
wire _12632_;
wire _12633_;
wire _12634_;
wire _12635_;
wire _12636_;
wire _12637_;
wire _12638_;
wire _12639_;
wire _12640_;
wire _12641_;
wire _12642_;
wire _12643_;
wire _12644_;
wire _12645_;
wire _12646_;
wire _12647_;
wire _12648_;
wire _12649_;
wire _12650_;
wire _12651_;
wire _12652_;
wire _12653_;
wire _12654_;
wire _12655_;
wire _12656_;
wire _12657_;
wire _12658_;
wire _12659_;
wire _12660_;
wire _12661_;
wire _12662_;
wire _12663_;
wire _12664_;
wire _12665_;
wire _12666_;
wire _12667_;
wire _12668_;
wire _12669_;
wire _12670_;
wire _12671_;
wire _12672_;
wire _12673_;
wire _12674_;
wire _12675_;
wire _12676_;
wire _12677_;
wire _12678_;
wire _12679_;
wire _12680_;
wire _12681_;
wire _12682_;
wire _12683_;
wire _12684_;
wire _12685_;
wire _12686_;
wire _12687_;
wire _12688_;
wire _12689_;
wire _12690_;
wire _12691_;
wire _12692_;
wire _12693_;
wire _12694_;
wire _12695_;
wire _12696_;
wire _12697_;
wire _12698_;
wire _12699_;
wire _12700_;
wire _12701_;
wire _12702_;
wire _12703_;
wire _12704_;
wire _12705_;
wire _12706_;
wire _12707_;
wire _12708_;
wire _12709_;
wire _12710_;
wire _12711_;
wire _12712_;
wire _12713_;
wire _12714_;
wire _12715_;
wire _12716_;
wire _12717_;
wire _12718_;
wire _12719_;
wire _12720_;
wire _12721_;
wire _12722_;
wire _12723_;
wire _12724_;
wire _12725_;
wire _12726_;
wire _12727_;
wire _12728_;
wire _12729_;
wire _12730_;
wire _12731_;
wire _12732_;
wire _12733_;
wire _12734_;
wire _12735_;
wire _12736_;
wire _12737_;
wire _12738_;
wire _12739_;
wire _12740_;
wire _12741_;
wire _12742_;
wire _12743_;
wire _12744_;
wire _12745_;
wire _12746_;
wire _12747_;
wire _12748_;
wire _12749_;
wire _12750_;
wire _12751_;
wire _12752_;
wire _12753_;
wire _12754_;
wire _12755_;
wire _12756_;
wire _12757_;
wire _12758_;
wire _12759_;
wire _12760_;
wire _12761_;
wire _12762_;
wire _12763_;
wire _12764_;
wire _12765_;
wire _12766_;
wire _12767_;
wire _12768_;
wire _12769_;
wire _12770_;
wire _12771_;
wire _12772_;
wire _12773_;
wire _12774_;
wire _12775_;
wire _12776_;
wire _12777_;
wire _12778_;
wire _12779_;
wire _12780_;
wire _12781_;
wire _12782_;
wire _12783_;
wire _12784_;
wire _12785_;
wire _12786_;
wire _12787_;
wire _12788_;
wire _12789_;
wire _12790_;
wire _12791_;
wire _12792_;
wire _12793_;
wire _12794_;
wire _12795_;
wire _12796_;
wire _12797_;
wire _12798_;
wire _12799_;
wire _12800_;
wire _12801_;
wire _12802_;
wire _12803_;
wire _12804_;
wire _12805_;
wire _12806_;
wire _12807_;
wire _12808_;
wire _12809_;
wire _12810_;
wire _12811_;
wire _12812_;
wire _12813_;
wire _12814_;
wire _12815_;
wire _12816_;
wire _12817_;
wire _12818_;
wire _12819_;
wire _12820_;
wire _12821_;
wire _12822_;
wire _12823_;
wire _12824_;
wire _12825_;
wire _12826_;
wire _12827_;
wire _12828_;
wire _12829_;
wire _12830_;
wire _12831_;
wire _12832_;
wire _12833_;
wire _12834_;
wire _12835_;
wire _12836_;
wire _12837_;
wire _12838_;
wire _12839_;
wire _12840_;
wire _12841_;
wire _12842_;
wire _12843_;
wire _12844_;
wire _12845_;
wire _12846_;
wire _12847_;
wire _12848_;
wire _12849_;
wire _12850_;
wire _12851_;
wire _12852_;
wire _12853_;
wire _12854_;
wire _12855_;
wire _12856_;
wire _12857_;
wire _12858_;
wire _12859_;
wire _12860_;
wire _12861_;
wire _12862_;
wire _12863_;
wire _12864_;
wire _12865_;
wire _12866_;
wire _12867_;
wire _12868_;
wire _12869_;
wire _12870_;
wire _12871_;
wire _12872_;
wire _12873_;
wire _12874_;
wire _12875_;
wire _12876_;
wire _12877_;
wire _12878_;
wire _12879_;
wire _12880_;
wire _12881_;
wire _12882_;
wire _12883_;
wire _12884_;
wire _12885_;
wire _12886_;
wire _12887_;
wire _12888_;
wire _12889_;
wire _12890_;
wire _12891_;
wire _12892_;
wire _12893_;
wire _12894_;
wire _12895_;
wire _12896_;
wire _12897_;
wire _12898_;
wire _12899_;
wire _12900_;
wire _12901_;
wire _12902_;
wire _12903_;
wire _12904_;
wire _12905_;
wire _12906_;
wire _12907_;
wire _12908_;
wire _12909_;
wire _12910_;
wire _12911_;
wire _12912_;
wire _12913_;
wire _12914_;
wire _12915_;
wire _12916_;
wire _12917_;
wire _12918_;
wire _12919_;
wire _12920_;
wire _12921_;
wire _12922_;
wire _12923_;
wire _12924_;
wire _12925_;
wire _12926_;
wire _12927_;
wire _12928_;
wire _12929_;
wire _12930_;
wire _12931_;
wire _12932_;
wire _12933_;
wire _12934_;
wire _12935_;
wire _12936_;
wire _12937_;
wire _12938_;
wire _12939_;
wire _12940_;
wire _12941_;
wire _12942_;
wire _12943_;
wire _12944_;
wire _12945_;
wire _12946_;
wire _12947_;
wire _12948_;
wire _12949_;
wire _12950_;
wire _12951_;
wire _12952_;
wire _12953_;
wire _12954_;
wire _12955_;
wire _12956_;
wire _12957_;
wire _12958_;
wire _12959_;
wire _12960_;
wire _12961_;
wire _12962_;
wire _12963_;
wire _12964_;
wire _12965_;
wire _12966_;
wire _12967_;
wire _12968_;
wire _12969_;
wire _12970_;
wire _12971_;
wire _12972_;
wire _12973_;
wire _12974_;
wire _12975_;
wire _12976_;
wire _12977_;
wire _12978_;
wire _12979_;
wire _12980_;
wire _12981_;
wire _12982_;
wire _12983_;
wire _12984_;
wire _12985_;
wire _12986_;
wire _12987_;
wire _12988_;
wire _12989_;
wire _12990_;
wire _12991_;
wire _12992_;
wire _12993_;
wire _12994_;
wire _12995_;
wire _12996_;
wire _12997_;
wire _12998_;
wire _12999_;
wire _13000_;
wire _13001_;
wire _13002_;
wire _13003_;
wire _13004_;
wire _13005_;
wire _13006_;
wire _13007_;
wire _13008_;
wire _13009_;
wire _13010_;
wire _13011_;
wire _13012_;
wire _13013_;
wire _13014_;
wire _13015_;
wire _13016_;
wire _13017_;
wire _13018_;
wire _13019_;
wire _13020_;
wire _13021_;
wire _13022_;
wire _13023_;
wire _13024_;
wire _13025_;
wire _13026_;
wire _13027_;
wire _13028_;
wire _13029_;
wire _13030_;
wire _13031_;
wire _13032_;
wire _13033_;
wire _13034_;
wire _13035_;
wire _13036_;
wire _13037_;
wire _13038_;
wire _13039_;
wire _13040_;
wire _13041_;
wire _13042_;
wire _13043_;
wire _13044_;
wire _13045_;
wire _13046_;
wire _13047_;
wire _13048_;
wire _13049_;
wire _13050_;
wire _13051_;
wire _13052_;
wire _13053_;
wire _13054_;
wire _13055_;
wire _13056_;
wire _13057_;
wire _13058_;
wire _13059_;
wire _13060_;
wire _13061_;
wire _13062_;
wire _13063_;
wire _13064_;
wire _13065_;
wire _13066_;
wire _13067_;
wire _13068_;
wire _13069_;
wire _13070_;
wire _13071_;
wire _13072_;
wire _13073_;
wire _13074_;
wire _13075_;
wire _13076_;
wire _13077_;
wire _13078_;
wire _13079_;
wire _13080_;
wire _13081_;
wire _13082_;
wire _13083_;
wire _13084_;
wire _13085_;
wire _13086_;
wire _13087_;
wire _13088_;
wire _13089_;
wire _13090_;
wire _13091_;
wire _13092_;
wire _13093_;
wire _13094_;
wire _13095_;
wire _13096_;
wire _13097_;
wire _13098_;
wire _13099_;
wire _13100_;
wire _13101_;
wire _13102_;
wire _13103_;
wire _13104_;
wire _13105_;
wire _13106_;
wire _13107_;
wire _13108_;
wire _13109_;
wire _13110_;
wire _13111_;
wire _13112_;
wire _13113_;
wire _13114_;
wire _13115_;
wire _13116_;
wire _13117_;
wire _13118_;
wire _13119_;
wire _13120_;
wire _13121_;
wire _13122_;
wire _13123_;
wire _13124_;
wire _13125_;
wire _13126_;
wire _13127_;
wire _13128_;
wire _13129_;
wire _13130_;
wire _13131_;
wire _13132_;
wire _13133_;
wire _13134_;
wire _13135_;
wire _13136_;
wire _13137_;
wire _13138_;
wire _13139_;
wire _13140_;
wire _13141_;
wire _13142_;
wire _13143_;
wire _13144_;
wire _13145_;
wire _13146_;
wire _13147_;
wire _13148_;
wire _13149_;
wire _13150_;
wire _13151_;
wire _13152_;
wire _13153_;
wire _13154_;
wire _13155_;
wire _13156_;
wire _13157_;
wire _13158_;
wire _13159_;
wire _13160_;
wire _13161_;
wire _13162_;
wire _13163_;
wire _13164_;
wire _13165_;
wire _13166_;
wire _13167_;
wire _13168_;
wire _13169_;
wire _13170_;
wire _13171_;
wire _13172_;
wire _13173_;
wire _13174_;
wire _13175_;
wire _13176_;
wire _13177_;
wire _13178_;
wire _13179_;
wire _13180_;
wire _13181_;
wire _13182_;
wire _13183_;
wire _13184_;
wire _13185_;
wire _13186_;
wire _13187_;
wire _13188_;
wire _13189_;
wire _13190_;
wire _13191_;
wire _13192_;
wire _13193_;
wire _13194_;
wire _13195_;
wire _13196_;
wire _13197_;
wire _13198_;
wire _13199_;
wire _13200_;
wire _13201_;
wire _13202_;
wire _13203_;
wire _13204_;
wire _13205_;
wire _13206_;
wire _13207_;
wire _13208_;
wire _13209_;
wire _13210_;
wire _13211_;
wire _13212_;
wire _13213_;
wire _13214_;
wire _13215_;
wire _13216_;
wire _13217_;
wire _13218_;
wire _13219_;
wire _13220_;
wire _13221_;
wire _13222_;
wire _13223_;
wire _13224_;
wire _13225_;
wire _13226_;
wire _13227_;
wire _13228_;
wire _13229_;
wire _13230_;
wire _13231_;
wire _13232_;
wire _13233_;
wire _13234_;
wire _13235_;
wire _13236_;
wire _13237_;
wire _13238_;
wire _13239_;
wire _13240_;
wire _13241_;
wire _13242_;
wire _13243_;
wire _13244_;
wire _13245_;
wire _13246_;
wire _13247_;
wire _13248_;
wire _13249_;
wire _13250_;
wire _13251_;
wire _13252_;
wire _13253_;
wire _13254_;
wire _13255_;
wire _13256_;
wire _13257_;
wire _13258_;
wire _13259_;
wire _13260_;
wire _13261_;
wire _13262_;
wire _13263_;
wire _13264_;
wire _13265_;
wire _13266_;
wire _13267_;
wire _13268_;
wire _13269_;
wire _13270_;
wire _13271_;
wire _13272_;
wire _13273_;
wire _13274_;
wire _13275_;
wire _13276_;
wire _13277_;
wire _13278_;
wire _13279_;
wire _13280_;
wire _13281_;
wire _13282_;
wire _13283_;
wire _13284_;
wire _13285_;
wire _13286_;
wire _13287_;
wire _13288_;
wire _13289_;
wire _13290_;
wire _13291_;
wire _13292_;
wire _13293_;
wire _13294_;
wire _13295_;
wire _13296_;
wire _13297_;
wire _13298_;
wire _13299_;
wire _13300_;
wire _13301_;
wire _13302_;
wire _13303_;
wire _13304_;
wire _13305_;
wire _13306_;
wire _13307_;
wire _13308_;
wire _13309_;
wire _13310_;
wire _13311_;
wire _13312_;
wire _13313_;
wire _13314_;
wire _13315_;
wire _13316_;
wire _13317_;
wire _13318_;
wire _13319_;
wire _13320_;
wire _13321_;
wire _13322_;
wire _13323_;
wire _13324_;
wire _13325_;
wire _13326_;
wire _13327_;
wire _13328_;
wire _13329_;
wire _13330_;
wire _13331_;
wire _13332_;
wire _13333_;
wire _13334_;
wire _13335_;
wire _13336_;
wire _13337_;
wire _13338_;
wire _13339_;
wire _13340_;
wire _13341_;
wire _13342_;
wire _13343_;
wire _13344_;
wire _13345_;
wire _13346_;
wire _13347_;
wire _13348_;
wire _13349_;
wire _13350_;
wire _13351_;
wire _13352_;
wire _13353_;
wire _13354_;
wire _13355_;
wire _13356_;
wire _13357_;
wire _13358_;
wire _13359_;
wire _13360_;
wire _13361_;
wire _13362_;
wire _13363_;
wire _13364_;
wire _13365_;
wire _13366_;
wire _13367_;
wire _13368_;
wire _13369_;
wire _13370_;
wire _13371_;
wire _13372_;
wire _13373_;
wire _13374_;
wire _13375_;
wire _13376_;
wire _13377_;
wire _13378_;
wire _13379_;
wire _13380_;
wire _13381_;
wire _13382_;
wire _13383_;
wire _13384_;
wire _13385_;
wire _13386_;
wire _13387_;
wire _13388_;
wire _13389_;
wire _13390_;
wire _13391_;
wire _13392_;
wire _13393_;
wire _13394_;
wire _13395_;
wire _13396_;
wire _13397_;
wire _13398_;
wire _13399_;
wire _13400_;
wire _13401_;
wire _13402_;
wire _13403_;
wire _13404_;
wire _13405_;
wire _13406_;
wire _13407_;
wire _13408_;
wire _13409_;
wire _13410_;
wire _13411_;
wire _13412_;
wire _13413_;
wire _13414_;
wire _13415_;
wire _13416_;
wire _13417_;
wire _13418_;
wire _13419_;
wire _13420_;
wire _13421_;
wire _13422_;
wire _13423_;
wire _13424_;
wire _13425_;
wire _13426_;
wire _13427_;
wire _13428_;
wire _13429_;
wire _13430_;
wire _13431_;
wire _13432_;
wire _13433_;
wire _13434_;
wire _13435_;
wire _13436_;
wire _13437_;
wire _13438_;
wire _13439_;
wire _13440_;
wire _13441_;
wire _13442_;
wire _13443_;
wire _13444_;
wire _13445_;
wire _13446_;
wire _13447_;
wire _13448_;
wire _13449_;
wire _13450_;
wire _13451_;
wire _13452_;
wire _13453_;
wire _13454_;
wire _13455_;
wire _13456_;
wire _13457_;
wire _13458_;
wire _13459_;
wire _13460_;
wire _13461_;
wire _13462_;
wire _13463_;
wire _13464_;
wire _13465_;
wire _13466_;
wire _13467_;
wire _13468_;
wire _13469_;
wire _13470_;
wire _13471_;
wire _13472_;
wire _13473_;
wire _13474_;
wire _13475_;
wire _13476_;
wire _13477_;
wire _13478_;
wire _13479_;
wire _13480_;
wire _13481_;
wire _13482_;
wire _13483_;
wire _13484_;
wire _13485_;
wire _13486_;
wire _13487_;
wire _13488_;
wire _13489_;
wire _13490_;
wire _13491_;
wire _13492_;
wire _13493_;
wire _13494_;
wire _13495_;
wire _13496_;
wire _13497_;
wire _13498_;
wire _13499_;
wire _13500_;
wire _13501_;
wire _13502_;
wire _13503_;
wire _13504_;
wire _13505_;
wire _13506_;
wire _13507_;
wire _13508_;
wire _13509_;
wire _13510_;
wire _13511_;
wire _13512_;
wire _13513_;
wire _13514_;
wire _13515_;
wire _13516_;
wire _13517_;
wire _13518_;
wire _13519_;
wire _13520_;
wire _13521_;
wire _13522_;
wire _13523_;
wire _13524_;
wire _13525_;
wire _13526_;
wire _13527_;
wire _13528_;
wire _13529_;
wire _13530_;
wire _13531_;
wire _13532_;
wire _13533_;
wire _13534_;
wire _13535_;
wire _13536_;
wire _13537_;
wire _13538_;
wire _13539_;
wire _13540_;
wire _13541_;
wire _13542_;
wire _13543_;
wire _13544_;
wire _13545_;
wire _13546_;
wire _13547_;
wire _13548_;
wire _13549_;
wire _13550_;
wire _13551_;
wire _13552_;
wire _13553_;
wire _13554_;
wire _13555_;
wire _13556_;
wire _13557_;
wire _13558_;
wire _13559_;
wire _13560_;
wire _13561_;
wire _13562_;
wire _13563_;
wire _13564_;
wire _13565_;
wire _13566_;
wire _13567_;
wire _13568_;
wire _13569_;
wire _13570_;
wire _13571_;
wire _13572_;
wire _13573_;
wire _13574_;
wire _13575_;
wire _13576_;
wire _13577_;
wire _13578_;
wire _13579_;
wire _13580_;
wire _13581_;
wire _13582_;
wire _13583_;
wire _13584_;
wire _13585_;
wire _13586_;
wire _13587_;
wire _13588_;
wire _13589_;
wire _13590_;
wire _13591_;
wire _13592_;
wire _13593_;
wire _13594_;
wire _13595_;
wire _13596_;
wire _13597_;
wire _13598_;
wire _13599_;
wire _13600_;
wire _13601_;
wire _13602_;
wire _13603_;
wire _13604_;
wire _13605_;
wire _13606_;
wire _13607_;
wire _13608_;
wire _13609_;
wire _13610_;
wire _13611_;
wire _13612_;
wire _13613_;
wire _13614_;
wire _13615_;
wire _13616_;
wire _13617_;
wire _13618_;
wire _13619_;
wire _13620_;
wire _13621_;
wire _13622_;
wire _13623_;
wire _13624_;
wire _13625_;
wire _13626_;
wire _13627_;
wire _13628_;
wire _13629_;
wire _13630_;
wire _13631_;
wire _13632_;
wire _13633_;
wire _13634_;
wire _13635_;
wire _13636_;
wire _13637_;
wire _13638_;
wire _13639_;
wire _13640_;
wire _13641_;
wire _13642_;
wire _13643_;
wire _13644_;
wire _13645_;
wire _13646_;
wire _13647_;
wire _13648_;
wire _13649_;
wire _13650_;
wire _13651_;
wire _13652_;
wire _13653_;
wire _13654_;
wire _13655_;
wire _13656_;
wire _13657_;
wire _13658_;
wire _13659_;
wire _13660_;
wire _13661_;
wire _13662_;
wire _13663_;
wire _13664_;
wire _13665_;
wire _13666_;
wire _13667_;
wire _13668_;
wire _13669_;
wire _13670_;
wire _13671_;
wire _13672_;
wire _13673_;
wire _13674_;
wire _13675_;
wire _13676_;
wire _13677_;
wire _13678_;
wire _13679_;
wire _13680_;
wire _13681_;
wire _13682_;
wire _13683_;
wire _13684_;
wire _13685_;
wire _13686_;
wire _13687_;
wire _13688_;
wire _13689_;
wire _13690_;
wire _13691_;
wire _13692_;
wire _13693_;
wire _13694_;
wire _13695_;
wire _13696_;
wire _13697_;
wire _13698_;
wire _13699_;
wire _13700_;
wire _13701_;
wire _13702_;
wire _13703_;
wire _13704_;
wire _13705_;
wire _13706_;
wire _13707_;
wire _13708_;
wire _13709_;
wire _13710_;
wire _13711_;
wire _13712_;
wire _13713_;
wire _13714_;
wire _13715_;
wire _13716_;
wire _13717_;
wire _13718_;
wire _13719_;
wire _13720_;
wire _13721_;
wire _13722_;
wire _13723_;
wire _13724_;
wire _13725_;
wire _13726_;
wire _13727_;
wire _13728_;
wire _13729_;
wire _13730_;
wire _13731_;
wire _13732_;
wire _13733_;
wire _13734_;
wire _13735_;
wire _13736_;
wire _13737_;
wire _13738_;
wire _13739_;
wire _13740_;
wire _13741_;
wire _13742_;
wire _13743_;
wire _13744_;
wire _13745_;
wire _13746_;
wire _13747_;
wire _13748_;
wire _13749_;
wire _13750_;
wire _13751_;
wire _13752_;
wire _13753_;
wire _13754_;
wire _13755_;
wire _13756_;
wire _13757_;
wire _13758_;
wire _13759_;
wire _13760_;
wire _13761_;
wire _13762_;
wire _13763_;
wire _13764_;
wire _13765_;
wire _13766_;
wire _13767_;
wire _13768_;
wire _13769_;
wire _13770_;
wire _13771_;
wire _13772_;
wire _13773_;
wire _13774_;
wire _13775_;
wire _13776_;
wire _13777_;
wire _13778_;
wire _13779_;
wire _13780_;
wire _13781_;
wire _13782_;
wire _13783_;
wire _13784_;
wire _13785_;
wire _13786_;
wire _13787_;
wire _13788_;
wire _13789_;
wire _13790_;
wire _13791_;
wire _13792_;
wire _13793_;
wire _13794_;
wire _13795_;
wire _13796_;
wire _13797_;
wire _13798_;
wire _13799_;
wire _13800_;
wire _13801_;
wire _13802_;
wire _13803_;
wire _13804_;
wire _13805_;
wire _13806_;
wire _13807_;
wire _13808_;
wire _13809_;
wire _13810_;
wire _13811_;
wire _13812_;
wire _13813_;
wire _13814_;
wire _13815_;
wire _13816_;
wire _13817_;
wire _13818_;
wire _13819_;
wire _13820_;
wire _13821_;
wire _13822_;
wire _13823_;
wire _13824_;
wire _13825_;
wire _13826_;
wire _13827_;
wire _13828_;
wire _13829_;
wire _13830_;
wire _13831_;
wire _13832_;
wire _13833_;
wire _13834_;
wire _13835_;
wire _13836_;
wire _13837_;
wire _13838_;
wire _13839_;
wire _13840_;
wire _13841_;
wire _13842_;
wire _13843_;
wire _13844_;
wire _13845_;
wire _13846_;
wire _13847_;
wire _13848_;
wire _13849_;
wire _13850_;
wire _13851_;
wire _13852_;
wire _13853_;
wire _13854_;
wire _13855_;
wire _13856_;
wire _13857_;
wire _13858_;
wire _13859_;
wire _13860_;
wire _13861_;
wire _13862_;
wire _13863_;
wire _13864_;
wire _13865_;
wire _13866_;
wire _13867_;
wire _13868_;
wire _13869_;
wire _13870_;
wire _13871_;
wire _13872_;
wire _13873_;
wire _13874_;
wire _13875_;
wire _13876_;
wire _13877_;
wire _13878_;
wire _13879_;
wire _13880_;
wire _13881_;
wire _13882_;
wire _13883_;
wire _13884_;
wire _13885_;
wire _13886_;
wire _13887_;
wire _13888_;
wire _13889_;
wire _13890_;
wire _13891_;
wire _13892_;
wire _13893_;
wire _13894_;
wire _13895_;
wire _13896_;
wire _13897_;
wire _13898_;
wire _13899_;
wire _13900_;
wire _13901_;
wire _13902_;
wire _13903_;
wire _13904_;
wire _13905_;
wire _13906_;
wire _13907_;
wire _13908_;
wire _13909_;
wire _13910_;
wire _13911_;
wire _13912_;
wire _13913_;
wire _13914_;
wire _13915_;
wire _13916_;
wire _13917_;
wire _13918_;
wire _13919_;
wire _13920_;
wire _13921_;
wire _13922_;
wire _13923_;
wire _13924_;
wire _13925_;
wire _13926_;
wire _13927_;
wire _13928_;
wire _13929_;
wire _13930_;
wire _13931_;
wire _13932_;
wire _13933_;
wire _13934_;
wire _13935_;
wire _13936_;
wire _13937_;
wire _13938_;
wire _13939_;
wire _13940_;
wire _13941_;
wire _13942_;
wire _13943_;
wire _13944_;
wire _13945_;
wire _13946_;
wire _13947_;
wire _13948_;
wire _13949_;
wire _13950_;
wire _13951_;
wire _13952_;
wire _13953_;
wire _13954_;
wire _13955_;
wire _13956_;
wire _13957_;
wire _13958_;
wire _13959_;
wire _13960_;
wire _13961_;
wire _13962_;
wire _13963_;
wire _13964_;
wire _13965_;
wire _13966_;
wire _13967_;
wire _13968_;
wire _13969_;
wire _13970_;
wire _13971_;
wire _13972_;
wire _13973_;
wire _13974_;
wire _13975_;
wire _13976_;
wire _13977_;
wire _13978_;
wire _13979_;
wire _13980_;
wire _13981_;
wire _13982_;
wire _13983_;
wire _13984_;
wire _13985_;
wire _13986_;
wire _13987_;
wire _13988_;
wire _13989_;
wire _13990_;
wire _13991_;
wire _13992_;
wire _13993_;
wire _13994_;
wire _13995_;
wire _13996_;
wire _13997_;
wire _13998_;
wire _13999_;
wire _14000_;
wire _14001_;
wire _14002_;
wire _14003_;
wire _14004_;
wire _14005_;
wire _14006_;
wire _14007_;
wire _14008_;
wire _14009_;
wire _14010_;
wire _14011_;
wire _14012_;
wire _14013_;
wire _14014_;
wire _14015_;
wire _14016_;
wire _14017_;
wire _14018_;
wire _14019_;
wire _14020_;
wire _14021_;
wire _14022_;
wire _14023_;
wire _14024_;
wire _14025_;
wire _14026_;
wire _14027_;
wire _14028_;
wire _14029_;
wire _14030_;
wire _14031_;
wire _14032_;
wire _14033_;
wire _14034_;
wire _14035_;
wire _14036_;
wire _14037_;
wire _14038_;
wire _14039_;
wire _14040_;
wire _14041_;
wire _14042_;
wire _14043_;
wire _14044_;
wire _14045_;
wire _14046_;
wire _14047_;
wire _14048_;
wire _14049_;
wire _14050_;
wire _14051_;
wire _14052_;
wire _14053_;
wire _14054_;
wire _14055_;
wire _14056_;
wire _14057_;
wire _14058_;
wire _14059_;
wire _14060_;
wire _14061_;
wire _14062_;
wire _14063_;
wire _14064_;
wire _14065_;
wire _14066_;
wire _14067_;
wire _14068_;
wire _14069_;
wire _14070_;
wire _14071_;
wire _14072_;
wire _14073_;
wire _14074_;
wire _14075_;
wire _14076_;
wire _14077_;
wire _14078_;
wire _14079_;
wire _14080_;
wire _14081_;
wire _14082_;
wire _14083_;
wire _14084_;
wire _14085_;
wire _14086_;
wire _14087_;
wire _14088_;
wire _14089_;
wire _14090_;
wire _14091_;
wire _14092_;
wire _14093_;
wire _14094_;
wire _14095_;
wire _14096_;
wire _14097_;
wire _14098_;
wire _14099_;
wire _14100_;
wire _14101_;
wire _14102_;
wire _14103_;
wire _14104_;
wire _14105_;
wire _14106_;
wire _14107_;
wire _14108_;
wire _14109_;
wire _14110_;
wire _14111_;
wire _14112_;
wire _14113_;
wire _14114_;
wire _14115_;
wire _14116_;
wire _14117_;
wire _14118_;
wire _14119_;
wire _14120_;
wire _14121_;
wire _14122_;
wire _14123_;
wire _14124_;
wire _14125_;
wire _14126_;
wire _14127_;
wire _14128_;
wire _14129_;
wire _14130_;
wire _14131_;
wire _14132_;
wire _14133_;
wire _14134_;
wire _14135_;
wire _14136_;
wire _14137_;
wire _14138_;
wire _14139_;
wire _14140_;
wire _14141_;
wire _14142_;
wire _14143_;
wire _14144_;
wire _14145_;
wire _14146_;
wire _14147_;
wire _14148_;
wire _14149_;
wire _14150_;
wire _14151_;
wire _14152_;
wire _14153_;
wire _14154_;
wire _14155_;
wire _14156_;
wire _14157_;
wire _14158_;
wire _14159_;
wire _14160_;
wire _14161_;
wire _14162_;
wire _14163_;
wire _14164_;
wire _14165_;
wire _14166_;
wire _14167_;
wire _14168_;
wire _14169_;
wire _14170_;
wire _14171_;
wire _14172_;
wire _14173_;
wire _14174_;
wire _14175_;
wire _14176_;
wire _14177_;
wire _14178_;
wire _14179_;
wire _14180_;
wire _14181_;
wire _14182_;
wire _14183_;
wire _14184_;
wire _14185_;
wire _14186_;
wire _14187_;
wire _14188_;
wire _14189_;
wire _14190_;
wire _14191_;
wire _14192_;
wire _14193_;
wire _14194_;
wire _14195_;
wire _14196_;
wire _14197_;
wire _14198_;
wire _14199_;
wire _14200_;
wire _14201_;
wire _14202_;
wire _14203_;
wire _14204_;
wire _14205_;
wire _14206_;
wire _14207_;
wire _14208_;
wire _14209_;
wire _14210_;
wire _14211_;
wire _14212_;
wire _14213_;
wire _14214_;
wire _14215_;
wire _14216_;
wire _14217_;
wire _14218_;
wire _14219_;
wire _14220_;
wire _14221_;
wire _14222_;
wire _14223_;
wire _14224_;
wire _14225_;
wire _14226_;
wire _14227_;
wire _14228_;
wire _14229_;
wire _14230_;
wire _14231_;
wire _14232_;
wire _14233_;
wire _14234_;
wire _14235_;
wire _14236_;
wire _14237_;
wire _14238_;
wire _14239_;
wire _14240_;
wire _14241_;
wire _14242_;
wire _14243_;
wire _14244_;
wire _14245_;
wire _14246_;
wire _14247_;
wire _14248_;
wire _14249_;
wire _14250_;
wire _14251_;
wire _14252_;
wire _14253_;
wire _14254_;
wire _14255_;
wire _14256_;
wire _14257_;
wire _14258_;
wire _14259_;
wire _14260_;
wire _14261_;
wire _14262_;
wire _14263_;
wire _14264_;
wire _14265_;
wire _14266_;
wire _14267_;
wire _14268_;
wire _14269_;
wire _14270_;
wire _14271_;
wire _14272_;
wire _14273_;
wire _14274_;
wire _14275_;
wire _14276_;
wire _14277_;
wire _14278_;
wire _14279_;
wire _14280_;
wire _14281_;
wire _14282_;
wire _14283_;
wire _14284_;
wire _14285_;
wire _14286_;
wire _14287_;
wire _14288_;
wire _14289_;
wire _14290_;
wire _14291_;
wire _14292_;
wire _14293_;
wire _14294_;
wire _14295_;
wire _14296_;
wire _14297_;
wire _14298_;
wire _14299_;
wire _14300_;
wire _14301_;
wire _14302_;
wire _14303_;
wire _14304_;
wire _14305_;
wire _14306_;
wire _14307_;
wire _14308_;
wire _14309_;
wire _14310_;
wire _14311_;
wire _14312_;
wire _14313_;
wire _14314_;
wire _14315_;
wire _14316_;
wire _14317_;
wire _14318_;
wire _14319_;
wire _14320_;
wire _14321_;
wire _14322_;
wire _14323_;
wire _14324_;
wire _14325_;
wire _14326_;
wire _14327_;
wire _14328_;
wire _14329_;
wire _14330_;
wire _14331_;
wire _14332_;
wire _14333_;
wire _14334_;
wire _14335_;
wire _14336_;
wire _14337_;
wire _14338_;
wire _14339_;
wire _14340_;
wire _14341_;
wire _14342_;
wire _14343_;
wire _14344_;
wire _14345_;
wire _14346_;
wire _14347_;
wire _14348_;
wire _14349_;
wire _14350_;
wire _14351_;
wire _14352_;
wire _14353_;
wire _14354_;
wire _14355_;
wire _14356_;
wire _14357_;
wire _14358_;
wire _14359_;
wire _14360_;
wire _14361_;
wire _14362_;
wire _14363_;
wire _14364_;
wire _14365_;
wire _14366_;
wire _14367_;
wire _14368_;
wire _14369_;
wire _14370_;
wire _14371_;
wire _14372_;
wire _14373_;
wire _14374_;
wire _14375_;
wire _14376_;
wire _14377_;
wire _14378_;
wire _14379_;
wire _14380_;
wire _14381_;
wire _14382_;
wire _14383_;
wire _14384_;
wire _14385_;
wire _14386_;
wire _14387_;
wire _14388_;
wire _14389_;
wire _14390_;
wire _14391_;
wire _14392_;
wire _14393_;
wire _14394_;
wire _14395_;
wire _14396_;
wire _14397_;
wire _14398_;
wire _14399_;
wire _14400_;
wire _14401_;
wire _14402_;
wire _14403_;
wire _14404_;
wire _14405_;
wire _14406_;
wire _14407_;
wire _14408_;
wire _14409_;
wire _14410_;
wire _14411_;
wire _14412_;
wire _14413_;
wire _14414_;
wire _14415_;
wire _14416_;
wire _14417_;
wire _14418_;
wire _14419_;
wire _14420_;
wire _14421_;
wire _14422_;
wire _14423_;
wire _14424_;
wire _14425_;
wire _14426_;
wire _14427_;
wire _14428_;
wire _14429_;
wire _14430_;
wire _14431_;
wire _14432_;
wire _14433_;
wire _14434_;
wire _14435_;
wire _14436_;
wire _14437_;
wire _14438_;
wire _14439_;
wire _14440_;
wire _14441_;
wire _14442_;
wire _14443_;
wire _14444_;
wire _14445_;
wire _14446_;
wire _14447_;
wire _14448_;
wire _14449_;
wire _14450_;
wire _14451_;
wire _14452_;
wire _14453_;
wire _14454_;
wire _14455_;
wire _14456_;
wire _14457_;
wire _14458_;
wire _14459_;
wire _14460_;
wire _14461_;
wire _14462_;
wire _14463_;
wire _14464_;
wire _14465_;
wire _14466_;
wire _14467_;
wire _14468_;
wire _14469_;
wire _14470_;
wire _14471_;
wire _14472_;
wire _14473_;
wire _14474_;
wire _14475_;
wire _14476_;
wire _14477_;
wire _14478_;
wire _14479_;
wire _14480_;
wire _14481_;
wire _14482_;
wire _14483_;
wire _14484_;
wire _14485_;
wire _14486_;
wire _14487_;
wire _14488_;
wire _14489_;
wire _14490_;
wire _14491_;
wire _14492_;
wire _14493_;
wire _14494_;
wire _14495_;
wire _14496_;
wire _14497_;
wire _14498_;
wire _14499_;
wire _14500_;
wire _14501_;
wire _14502_;
wire _14503_;
wire _14504_;
wire _14505_;
wire _14506_;
wire _14507_;
wire _14508_;
wire _14509_;
wire _14510_;
wire _14511_;
wire _14512_;
wire _14513_;
wire _14514_;
wire _14515_;
wire _14516_;
wire _14517_;
wire _14518_;
wire _14519_;
wire _14520_;
wire _14521_;
wire _14522_;
wire _14523_;
wire _14524_;
wire _14525_;
wire _14526_;
wire _14527_;
wire _14528_;
wire _14529_;
wire _14530_;
wire _14531_;
wire _14532_;
wire _14533_;
wire _14534_;
wire _14535_;
wire _14536_;
wire _14537_;
wire _14538_;
wire _14539_;
wire _14540_;
wire _14541_;
wire _14542_;
wire _14543_;
wire _14544_;
wire _14545_;
wire _14546_;
wire _14547_;
wire _14548_;
wire _14549_;
wire _14550_;
wire _14551_;
wire _14552_;
wire _14553_;
wire _14554_;
wire _14555_;
wire _14556_;
wire _14557_;
wire _14558_;
wire _14559_;
wire _14560_;
wire _14561_;
wire _14562_;
wire _14563_;
wire _14564_;
wire _14565_;
wire _14566_;
wire _14567_;
wire _14568_;
wire _14569_;
wire _14570_;
wire _14571_;
wire _14572_;
wire _14573_;
wire _14574_;
wire _14575_;
wire _14576_;
wire _14577_;
wire _14578_;
wire _14579_;
wire _14580_;
wire _14581_;
wire _14582_;
wire _14583_;
wire _14584_;
wire _14585_;
wire _14586_;
wire _14587_;
wire _14588_;
wire _14589_;
wire _14590_;
wire _14591_;
wire _14592_;
wire _14593_;
wire _14594_;
wire _14595_;
wire _14596_;
wire _14597_;
wire _14598_;
wire _14599_;
wire _14600_;
wire _14601_;
wire _14602_;
wire _14603_;
wire _14604_;
wire _14605_;
wire _14606_;
wire _14607_;
wire _14608_;
wire _14609_;
wire _14610_;
wire _14611_;
wire _14612_;
wire _14613_;
wire _14614_;
wire _14615_;
wire _14616_;
wire _14617_;
wire _14618_;
wire _14619_;
wire _14620_;
wire _14621_;
wire _14622_;
wire _14623_;
wire _14624_;
wire _14625_;
wire _14626_;
wire _14627_;
wire _14628_;
wire _14629_;
wire _14630_;
wire _14631_;
wire _14632_;
wire _14633_;
wire _14634_;
wire _14635_;
wire _14636_;
wire _14637_;
wire _14638_;
wire _14639_;
wire _14640_;
wire _14641_;
wire _14642_;
wire _14643_;
wire _14644_;
wire _14645_;
wire _14646_;
wire _14647_;
wire _14648_;
wire _14649_;
wire _14650_;
wire _14651_;
wire _14652_;
wire _14653_;
wire _14654_;
wire _14655_;
wire _14656_;
wire _14657_;
wire _14658_;
wire _14659_;
wire _14660_;
wire _14661_;
wire _14662_;
wire _14663_;
wire _14664_;
wire _14665_;
wire _14666_;
wire _14667_;
wire _14668_;
wire _14669_;
wire _14670_;
wire _14671_;
wire _14672_;
wire _14673_;
wire _14674_;
wire _14675_;
wire _14676_;
wire _14677_;
wire _14678_;
wire _14679_;
wire _14680_;
wire _14681_;
wire _14682_;
wire _14683_;
wire _14684_;
wire _14685_;
wire _14686_;
wire _14687_;
wire _14688_;
wire _14689_;
wire _14690_;
wire _14691_;
wire _14692_;
wire _14693_;
wire _14694_;
wire _14695_;
wire _14696_;
wire _14697_;
wire _14698_;
wire _14699_;
wire _14700_;
wire _14701_;
wire _14702_;
wire _14703_;
wire _14704_;
wire _14705_;
wire _14706_;
wire _14707_;
wire _14708_;
wire _14709_;
wire _14710_;
wire _14711_;
wire _14712_;
wire _14713_;
wire _14714_;
wire _14715_;
wire _14716_;
wire _14717_;
wire _14718_;
wire _14719_;
wire _14720_;
wire _14721_;
wire _14722_;
wire _14723_;
wire _14724_;
wire _14725_;
wire _14726_;
wire _14727_;
wire _14728_;
wire _14729_;
wire _14730_;
wire _14731_;
wire _14732_;
wire _14733_;
wire _14734_;
wire _14735_;
wire _14736_;
wire _14737_;
wire _14738_;
wire _14739_;
wire _14740_;
wire _14741_;
wire _14742_;
wire _14743_;
wire _14744_;
wire _14745_;
wire _14746_;
wire _14747_;
wire _14748_;
wire _14749_;
wire _14750_;
wire _14751_;
wire _14752_;
wire _14753_;
wire _14754_;
wire _14755_;
wire _14756_;
wire _14757_;
wire _14758_;
wire _14759_;
wire _14760_;
wire _14761_;
wire _14762_;
wire _14763_;
wire _14764_;
wire _14765_;
wire _14766_;
wire _14767_;
wire _14768_;
wire _14769_;
wire _14770_;
wire _14771_;
wire _14772_;
wire _14773_;
wire _14774_;
wire _14775_;
wire _14776_;
wire _14777_;
wire _14778_;
wire _14779_;
wire _14780_;
wire _14781_;
wire _14782_;
wire _14783_;
wire _14784_;
wire _14785_;
wire _14786_;
wire _14787_;
wire _14788_;
wire _14789_;
wire _14790_;
wire _14791_;
wire _14792_;
wire _14793_;
wire _14794_;
wire _14795_;
wire _14796_;
wire _14797_;
wire _14798_;
wire _14799_;
wire _14800_;
wire _14801_;
wire _14802_;
wire _14803_;
wire _14804_;
wire _14805_;
wire _14806_;
wire _14807_;
wire _14808_;
wire _14809_;
wire _14810_;
wire _14811_;
wire _14812_;
wire _14813_;
wire _14814_;
wire _14815_;
wire _14816_;
wire _14817_;
wire _14818_;
wire _14819_;
wire _14820_;
wire _14821_;
wire _14822_;
wire _14823_;
wire _14824_;
wire _14825_;
wire _14826_;
wire _14827_;
wire _14828_;
wire _14829_;
wire _14830_;
wire _14831_;
wire _14832_;
wire _14833_;
wire _14834_;
wire _14835_;
wire _14836_;
wire _14837_;
wire _14838_;
wire _14839_;
wire _14840_;
wire _14841_;
wire _14842_;
wire _14843_;
wire _14844_;
wire _14845_;
wire _14846_;
wire _14847_;
wire _14848_;
wire _14849_;
wire _14850_;
wire _14851_;
wire _14852_;
wire _14853_;
wire _14854_;
wire _14855_;
wire _14856_;
wire _14857_;
wire _14858_;
wire _14859_;
wire _14860_;
wire _14861_;
wire _14862_;
wire _14863_;
wire _14864_;
wire _14865_;
wire _14866_;
wire _14867_;
wire _14868_;
wire _14869_;
wire _14870_;
wire _14871_;
wire _14872_;
wire _14873_;
wire _14874_;
wire _14875_;
wire _14876_;
wire _14877_;
wire _14878_;
wire _14879_;
wire _14880_;
wire _14881_;
wire _14882_;
wire _14883_;
wire _14884_;
wire _14885_;
wire _14886_;
wire _14887_;
wire _14888_;
wire _14889_;
wire _14890_;
wire _14891_;
wire _14892_;
wire _14893_;
wire _14894_;
wire _14895_;
wire _14896_;
wire _14897_;
wire _14898_;
wire _14899_;
wire _14900_;
wire _14901_;
wire _14902_;
wire _14903_;
wire _14904_;
wire _14905_;
wire _14906_;
wire _14907_;
wire _14908_;
wire _14909_;
wire _14910_;
wire _14911_;
wire _14912_;
wire _14913_;
wire _14914_;
wire _14915_;
wire _14916_;
wire _14917_;
wire _14918_;
wire _14919_;
wire _14920_;
wire _14921_;
wire _14922_;
wire _14923_;
wire _14924_;
wire _14925_;
wire _14926_;
wire _14927_;
wire _14928_;
wire _14929_;
wire _14930_;
wire _14931_;
wire _14932_;
wire _14933_;
wire _14934_;
wire _14935_;
wire _14936_;
wire _14937_;
wire _14938_;
wire _14939_;
wire _14940_;
wire _14941_;
wire _14942_;
wire _14943_;
wire _14944_;
wire _14945_;
wire _14946_;
wire _14947_;
wire _14948_;
wire _14949_;
wire _14950_;
wire _14951_;
wire _14952_;
wire _14953_;
wire _14954_;
wire _14955_;
wire _14956_;
wire _14957_;
wire _14958_;
wire _14959_;
wire _14960_;
wire _14961_;
wire _14962_;
wire _14963_;
wire _14964_;
wire _14965_;
wire _14966_;
wire _14967_;
wire _14968_;
wire _14969_;
wire _14970_;
wire _14971_;
wire _14972_;
wire _14973_;
wire _14974_;
wire _14975_;
wire _14976_;
wire _14977_;
wire _14978_;
wire _14979_;
wire _14980_;
wire _14981_;
wire _14982_;
wire _14983_;
wire _14984_;
wire _14985_;
wire _14986_;
wire _14987_;
wire _14988_;
wire _14989_;
wire _14990_;
wire _14991_;
wire _14992_;
wire _14993_;
wire _14994_;
wire _14995_;
wire _14996_;
wire _14997_;
wire _14998_;
wire _14999_;
wire _15000_;
wire _15001_;
wire _15002_;
wire _15003_;
wire _15004_;
wire _15005_;
wire _15006_;
wire _15007_;
wire _15008_;
wire _15009_;
wire _15010_;
wire _15011_;
wire _15012_;
wire _15013_;
wire _15014_;
wire _15015_;
wire _15016_;
wire _15017_;
wire _15018_;
wire _15019_;
wire _15020_;
wire _15021_;
wire _15022_;
wire _15023_;
wire _15024_;
wire _15025_;
wire _15026_;
wire _15027_;
wire _15028_;
wire _15029_;
wire _15030_;
wire _15031_;
wire _15032_;
wire _15033_;
wire _15034_;
wire _15035_;
wire _15036_;
wire _15037_;
wire _15038_;
wire _15039_;
wire _15040_;
wire _15041_;
wire _15042_;
wire _15043_;
wire _15044_;
wire _15045_;
wire _15046_;
wire _15047_;
wire _15048_;
wire _15049_;
wire _15050_;
wire _15051_;
wire _15052_;
wire _15053_;
wire _15054_;
wire _15055_;
wire _15056_;
wire _15057_;
wire _15058_;
wire _15059_;
wire _15060_;
wire _15061_;
wire _15062_;
wire _15063_;
wire _15064_;
wire _15065_;
wire _15066_;
wire _15067_;
wire _15068_;
wire _15069_;
wire _15070_;
wire _15071_;
wire _15072_;
wire _15073_;
wire _15074_;
wire _15075_;
wire _15076_;
wire _15077_;
wire _15078_;
wire _15079_;
wire _15080_;
wire _15081_;
wire _15082_;
wire _15083_;
wire _15084_;
wire _15085_;
wire _15086_;
wire _15087_;
wire _15088_;
wire _15089_;
wire _15090_;
wire _15091_;
wire _15092_;
wire _15093_;
wire _15094_;
wire _15095_;
wire _15096_;
wire _15097_;
wire _15098_;
wire _15099_;
wire _15100_;
wire _15101_;
wire _15102_;
wire _15103_;
wire _15104_;
wire _15105_;
wire _15106_;
wire _15107_;
wire _15108_;
wire _15109_;
wire _15110_;
wire _15111_;
wire _15112_;
wire _15113_;
wire _15114_;
wire _15115_;
wire _15116_;
wire _15117_;
wire _15118_;
wire _15119_;
wire _15120_;
wire _15121_;
wire _15122_;
wire _15123_;
wire _15124_;
wire _15125_;
wire _15126_;
wire _15127_;
wire _15128_;
wire _15129_;
wire _15130_;
wire _15131_;
wire _15132_;
wire _15133_;
wire _15134_;
wire _15135_;
wire _15136_;
wire _15137_;
wire _15138_;
wire _15139_;
wire _15140_;
wire _15141_;
wire _15142_;
wire _15143_;
wire _15144_;
wire _15145_;
wire _15146_;
wire _15147_;
wire _15148_;
wire _15149_;
wire _15150_;
wire _15151_;
wire _15152_;
wire _15153_;
wire _15154_;
wire _15155_;
wire _15156_;
wire _15157_;
wire _15158_;
wire _15159_;
wire _15160_;
wire _15161_;
wire _15162_;
wire _15163_;
wire _15164_;
wire _15165_;
wire _15166_;
wire _15167_;
wire _15168_;
wire _15169_;
wire _15170_;
wire _15171_;
wire _15172_;
wire _15173_;
wire _15174_;
wire _15175_;
wire _15176_;
wire _15177_;
wire _15178_;
wire _15179_;
wire _15180_;
wire _15181_;
wire _15182_;
wire _15183_;
wire _15184_;
wire _15185_;
wire _15186_;
wire _15187_;
wire _15188_;
wire _15189_;
wire _15190_;
wire _15191_;
wire _15192_;
wire _15193_;
wire _15194_;
wire _15195_;
wire _15196_;
wire _15197_;
wire _15198_;
wire _15199_;
wire _15200_;
wire _15201_;
wire _15202_;
wire _15203_;
wire _15204_;
wire _15205_;
wire _15206_;
wire _15207_;
wire _15208_;
wire _15209_;
wire _15210_;
wire _15211_;
wire _15212_;
wire _15213_;
wire _15214_;
wire _15215_;
wire _15216_;
wire _15217_;
wire _15218_;
wire _15219_;
wire _15220_;
wire _15221_;
wire _15222_;
wire _15223_;
wire _15224_;
wire _15225_;
wire _15226_;
wire _15227_;
wire _15228_;
wire _15229_;
wire _15230_;
wire _15231_;
wire _15232_;
wire _15233_;
wire _15234_;
wire _15235_;
wire _15236_;
wire _15237_;
wire _15238_;
wire _15239_;
wire _15240_;
wire _15241_;
wire _15242_;
wire _15243_;
wire _15244_;
wire _15245_;
wire _15246_;
wire _15247_;
wire _15248_;
wire _15249_;
wire _15250_;
wire _15251_;
wire _15252_;
wire _15253_;
wire _15254_;
wire _15255_;
wire _15256_;
wire _15257_;
wire _15258_;
wire _15259_;
wire _15260_;
wire _15261_;
wire _15262_;
wire _15263_;
wire _15264_;
wire _15265_;
wire _15266_;
wire _15267_;
wire _15268_;
wire _15269_;
wire _15270_;
wire _15271_;
wire _15272_;
wire _15273_;
wire _15274_;
wire _15275_;
wire _15276_;
wire _15277_;
wire _15278_;
wire _15279_;
wire _15280_;
wire _15281_;
wire _15282_;
wire _15283_;
wire _15284_;
wire _15285_;
wire _15286_;
wire _15287_;
wire _15288_;
wire _15289_;
wire _15290_;
wire _15291_;
wire _15292_;
wire _15293_;
wire _15294_;
wire _15295_;
wire _15296_;
wire _15297_;
wire _15298_;
wire _15299_;
wire _15300_;
wire _15301_;
wire _15302_;
wire _15303_;
wire _15304_;
wire _15305_;
wire _15306_;
wire _15307_;
wire _15308_;
wire _15309_;
wire _15310_;
wire _15311_;
wire _15312_;
wire _15313_;
wire _15314_;
wire _15315_;
wire _15316_;
wire _15317_;
wire _15318_;
wire _15319_;
wire _15320_;
wire _15321_;
wire _15322_;
wire _15323_;
wire _15324_;
wire _15325_;
wire _15326_;
wire _15327_;
wire _15328_;
wire _15329_;
wire _15330_;
wire _15331_;
wire _15332_;
wire _15333_;
wire _15334_;
wire _15335_;
wire _15336_;
wire _15337_;
wire _15338_;
wire _15339_;
wire _15340_;
wire _15341_;
wire _15342_;
wire _15343_;
wire _15344_;
wire _15345_;
wire _15346_;
wire _15347_;
wire _15348_;
wire _15349_;
wire _15350_;
wire _15351_;
wire _15352_;
wire _15353_;
wire _15354_;
wire _15355_;
wire _15356_;
wire _15357_;
wire _15358_;
wire _15359_;
wire _15360_;
wire _15361_;
wire _15362_;
wire _15363_;
wire _15364_;
wire _15365_;
wire _15366_;
wire _15367_;
wire _15368_;
wire _15369_;
wire _15370_;
wire _15371_;
wire _15372_;
wire _15373_;
wire _15374_;
wire _15375_;
wire _15376_;
wire _15377_;
wire _15378_;
wire _15379_;
wire _15380_;
wire _15381_;
wire _15382_;
wire _15383_;
wire _15384_;
wire _15385_;
wire _15386_;
wire _15387_;
wire _15388_;
wire _15389_;
wire _15390_;
wire _15391_;
wire _15392_;
wire _15393_;
wire _15394_;
wire _15395_;
wire _15396_;
wire _15397_;
wire _15398_;
wire _15399_;
wire _15400_;
wire _15401_;
wire _15402_;
wire _15403_;
wire _15404_;
wire _15405_;
wire _15406_;
wire _15407_;
wire _15408_;
wire _15409_;
wire _15410_;
wire _15411_;
wire _15412_;
wire _15413_;
wire _15414_;
wire _15415_;
wire _15416_;
wire _15417_;
wire _15418_;
wire _15419_;
wire _15420_;
wire _15421_;
wire _15422_;
wire _15423_;
wire _15424_;
wire _15425_;
wire _15426_;
wire _15427_;
wire _15428_;
wire _15429_;
wire _15430_;
wire _15431_;
wire _15432_;
wire _15433_;
wire _15434_;
wire _15435_;
wire _15436_;
wire _15437_;
wire _15438_;
wire _15439_;
wire _15440_;
wire _15441_;
wire _15442_;
wire _15443_;
wire _15444_;
wire _15445_;
wire _15446_;
wire _15447_;
wire _15448_;
wire _15449_;
wire _15450_;
wire _15451_;
wire _15452_;
wire _15453_;
wire _15454_;
wire _15455_;
wire _15456_;
wire _15457_;
wire _15458_;
wire _15459_;
wire _15460_;
wire _15461_;
wire _15462_;
wire _15463_;
wire _15464_;
wire _15465_;
wire _15466_;
wire _15467_;
wire _15468_;
wire _15469_;
wire _15470_;
wire _15471_;
wire _15472_;
wire _15473_;
wire _15474_;
wire _15475_;
wire _15476_;
wire _15477_;
wire _15478_;
wire _15479_;
wire _15480_;
wire _15481_;
wire _15482_;
wire _15483_;
wire _15484_;
wire _15485_;
wire _15486_;
wire _15487_;
wire _15488_;
wire _15489_;
wire _15490_;
wire _15491_;
wire _15492_;
wire _15493_;
wire _15494_;
wire _15495_;
wire _15496_;
wire _15497_;
wire _15498_;
wire _15499_;
wire _15500_;
wire _15501_;
wire _15502_;
wire _15503_;
wire _15504_;
wire _15505_;
wire _15506_;
wire _15507_;
wire _15508_;
wire _15509_;
wire _15510_;
wire _15511_;
wire _15512_;
wire _15513_;
wire _15514_;
wire _15515_;
wire _15516_;
wire _15517_;
wire _15518_;
wire _15519_;
wire _15520_;
wire _15521_;
wire _15522_;
wire _15523_;
wire _15524_;
wire _15525_;
wire _15526_;
wire _15527_;
wire _15528_;
wire _15529_;
wire _15530_;
wire _15531_;
wire _15532_;
wire _15533_;
wire _15534_;
wire _15535_;
wire _15536_;
wire _15537_;
wire _15538_;
wire _15539_;
wire _15540_;
wire _15541_;
wire _15542_;
wire _15543_;
wire _15544_;
wire _15545_;
wire _15546_;
wire _15547_;
wire _15548_;
wire _15549_;
wire _15550_;
wire _15551_;
wire _15552_;
wire _15553_;
wire _15554_;
wire _15555_;
wire _15556_;
wire _15557_;
wire _15558_;
wire _15559_;
wire _15560_;
wire _15561_;
wire _15562_;
wire _15563_;
wire _15564_;
wire _15565_;
wire _15566_;
wire _15567_;
wire _15568_;
wire _15569_;
wire _15570_;
wire _15571_;
wire _15572_;
wire _15573_;
wire _15574_;
wire _15575_;
wire _15576_;
wire _15577_;
wire _15578_;
wire _15579_;
wire _15580_;
wire _15581_;
wire _15582_;
wire _15583_;
wire _15584_;
wire _15585_;
wire _15586_;
wire _15587_;
wire _15588_;
wire _15589_;
wire _15590_;
wire _15591_;
wire _15592_;
wire _15593_;
wire _15594_;
wire _15595_;
wire _15596_;
wire _15597_;
wire _15598_;
wire _15599_;
wire _15600_;
wire _15601_;
wire _15602_;
wire _15603_;
wire _15604_;
wire _15605_;
wire _15606_;
wire _15607_;
wire _15608_;
wire _15609_;
wire _15610_;
wire _15611_;
wire _15612_;
wire _15613_;
wire _15614_;
wire _15615_;
wire _15616_;
wire _15617_;
wire _15618_;
wire _15619_;
wire _15620_;
wire _15621_;
wire _15622_;
wire _15623_;
wire _15624_;
wire _15625_;
wire _15626_;
wire _15627_;
wire _15628_;
wire _15629_;
wire _15630_;
wire _15631_;
wire _15632_;
wire _15633_;
wire _15634_;
wire _15635_;
wire _15636_;
wire _15637_;
wire _15638_;
wire _15639_;
wire _15640_;
wire _15641_;
wire _15642_;
wire _15643_;
wire _15644_;
wire _15645_;
wire _15646_;
wire _15647_;
wire _15648_;
wire _15649_;
wire _15650_;
wire _15651_;
wire _15652_;
wire _15653_;
wire _15654_;
wire _15655_;
wire _15656_;
wire _15657_;
wire _15658_;
wire _15659_;
wire _15660_;
wire _15661_;
wire _15662_;
wire _15663_;
wire _15664_;
wire _15665_;
wire _15666_;
wire _15667_;
wire _15668_;
wire _15669_;
wire _15670_;
wire _15671_;
wire _15672_;
wire _15673_;
wire _15674_;
wire _15675_;
wire _15676_;
wire _15677_;
wire _15678_;
wire _15679_;
wire _15680_;
wire _15681_;
wire _15682_;
wire _15683_;
wire _15684_;
wire _15685_;
wire _15686_;
wire _15687_;
wire _15688_;
wire _15689_;
wire _15690_;
wire _15691_;
wire _15692_;
wire _15693_;
wire _15694_;
wire _15695_;
wire _15696_;
wire _15697_;
wire _15698_;
wire _15699_;
wire _15700_;
wire _15701_;
wire _15702_;
wire _15703_;
wire _15704_;
wire _15705_;
wire _15706_;
wire _15707_;
wire _15708_;
wire _15709_;
wire _15710_;
wire _15711_;
wire _15712_;
wire _15713_;
wire _15714_;
wire _15715_;
wire _15716_;
wire _15717_;
wire _15718_;
wire _15719_;
wire _15720_;
wire _15721_;
wire _15722_;
wire _15723_;
wire _15724_;
wire _15725_;
wire _15726_;
wire _15727_;
wire _15728_;
wire _15729_;
wire _15730_;
wire _15731_;
wire _15732_;
wire _15733_;
wire _15734_;
wire _15735_;
wire _15736_;
wire _15737_;
wire _15738_;
wire _15739_;
wire _15740_;
wire _15741_;
wire _15742_;
wire _15743_;
wire _15744_;
wire _15745_;
wire _15746_;
wire _15747_;
wire _15748_;
wire _15749_;
wire _15750_;
wire _15751_;
wire _15752_;
wire _15753_;
wire _15754_;
wire _15755_;
wire _15756_;
wire _15757_;
wire _15758_;
wire _15759_;
wire _15760_;
wire _15761_;
wire _15762_;
wire _15763_;
wire _15764_;
wire _15765_;
wire _15766_;
wire _15767_;
wire _15768_;
wire _15769_;
wire _15770_;
wire _15771_;
wire _15772_;
wire _15773_;
wire _15774_;
wire _15775_;
wire _15776_;
wire _15777_;
wire _15778_;
wire _15779_;
wire _15780_;
wire _15781_;
wire _15782_;
wire _15783_;
wire _15784_;
wire _15785_;
wire _15786_;
wire _15787_;
wire _15788_;
wire _15789_;
wire _15790_;
wire _15791_;
wire _15792_;
wire _15793_;
wire _15794_;
wire _15795_;
wire _15796_;
wire _15797_;
wire _15798_;
wire _15799_;
wire _15800_;
wire _15801_;
wire _15802_;
wire _15803_;
wire _15804_;
wire _15805_;
wire _15806_;
wire _15807_;
wire _15808_;
wire _15809_;
wire _15810_;
wire _15811_;
wire _15812_;
wire _15813_;
wire _15814_;
wire _15815_;
wire _15816_;
wire _15817_;
wire _15818_;
wire _15819_;
wire _15820_;
wire _15821_;
wire _15822_;
wire _15823_;
wire _15824_;
wire _15825_;
wire _15826_;
wire _15827_;
wire _15828_;
wire _15829_;
wire _15830_;
wire _15831_;
wire _15832_;
wire _15833_;
wire _15834_;
wire _15835_;
wire _15836_;
wire _15837_;
wire _15838_;
wire _15839_;
wire _15840_;
wire _15841_;
wire _15842_;
wire _15843_;
wire _15844_;
wire _15845_;
wire _15846_;
wire _15847_;
wire _15848_;
wire _15849_;
wire _15850_;
wire _15851_;
wire _15852_;
wire _15853_;
wire _15854_;
wire _15855_;
wire _15856_;
wire _15857_;
wire _15858_;
wire _15859_;
wire _15860_;
wire _15861_;
wire _15862_;
wire _15863_;
wire _15864_;
wire _15865_;
wire _15866_;
wire _15867_;
wire _15868_;
wire _15869_;
wire _15870_;
wire _15871_;
wire _15872_;
wire _15873_;
wire _15874_;
wire _15875_;
wire _15876_;
wire _15877_;
wire _15878_;
wire _15879_;
wire _15880_;
wire _15881_;
wire _15882_;
wire _15883_;
wire _15884_;
wire _15885_;
wire _15886_;
wire _15887_;
wire _15888_;
wire _15889_;
wire _15890_;
wire _15891_;
wire _15892_;
wire _15893_;
wire _15894_;
wire _15895_;
wire _15896_;
wire _15897_;
wire _15898_;
wire _15899_;
wire _15900_;
wire _15901_;
wire _15902_;
wire _15903_;
wire _15904_;
wire _15905_;
wire _15906_;
wire _15907_;
wire _15908_;
wire _15909_;
wire _15910_;
wire _15911_;
wire _15912_;
wire _15913_;
wire _15914_;
wire _15915_;
wire _15916_;
wire _15917_;
wire _15918_;
wire _15919_;
wire _15920_;
wire _15921_;
wire _15922_;
wire _15923_;
wire _15924_;
wire _15925_;
wire _15926_;
wire _15927_;
wire _15928_;
wire _15929_;
wire _15930_;
wire _15931_;
wire _15932_;
wire _15933_;
wire _15934_;
wire _15935_;
wire _15936_;
wire _15937_;
wire _15938_;
wire _15939_;
wire _15940_;
wire _15941_;
wire _15942_;
wire _15943_;
wire _15944_;
wire _15945_;
wire _15946_;
wire _15947_;
wire _15948_;
wire _15949_;
wire _15950_;
wire _15951_;
wire _15952_;
wire _15953_;
wire _15954_;
wire _15955_;
wire _15956_;
wire _15957_;
wire _15958_;
wire _15959_;
wire _15960_;
wire _15961_;
wire _15962_;
wire _15963_;
wire _15964_;
wire _15965_;
wire _15966_;
wire _15967_;
wire _15968_;
wire _15969_;
wire _15970_;
wire _15971_;
wire _15972_;
wire _15973_;
wire _15974_;
wire _15975_;
wire _15976_;
wire _15977_;
wire _15978_;
wire _15979_;
wire _15980_;
wire _15981_;
wire _15982_;
wire _15983_;
wire _15984_;
wire _15985_;
wire _15986_;
wire _15987_;
wire _15988_;
wire _15989_;
wire _15990_;
wire _15991_;
wire _15992_;
wire _15993_;
wire _15994_;
wire _15995_;
wire _15996_;
wire _15997_;
wire _15998_;
wire _15999_;
wire _16000_;
wire _16001_;
wire _16002_;
wire _16003_;
wire _16004_;
wire _16005_;
wire _16006_;
wire _16007_;
wire _16008_;
wire _16009_;
wire _16010_;
wire _16011_;
wire _16012_;
wire _16013_;
wire _16014_;
wire _16015_;
wire _16016_;
wire _16017_;
wire _16018_;
wire _16019_;
wire _16020_;
wire _16021_;
wire _16022_;
wire _16023_;
wire _16024_;
wire _16025_;
wire _16026_;
wire _16027_;
wire _16028_;
wire _16029_;
wire _16030_;
wire _16031_;
wire _16032_;
wire _16033_;
wire _16034_;
wire _16035_;
wire _16036_;
wire _16037_;
wire _16038_;
wire _16039_;
wire _16040_;
wire _16041_;
wire _16042_;
wire _16043_;
wire _16044_;
wire _16045_;
wire _16046_;
wire _16047_;
wire _16048_;
wire _16049_;
wire _16050_;
wire _16051_;
wire _16052_;
wire _16053_;
wire _16054_;
wire _16055_;
wire _16056_;
wire _16057_;
wire _16058_;
wire _16059_;
wire _16060_;
wire _16061_;
wire _16062_;
wire _16063_;
wire _16064_;
wire _16065_;
wire _16066_;
wire _16067_;
wire _16068_;
wire _16069_;
wire _16070_;
wire _16071_;
wire _16072_;
wire _16073_;
wire _16074_;
wire _16075_;
wire _16076_;
wire _16077_;
wire _16078_;
wire _16079_;
wire _16080_;
wire _16081_;
wire _16082_;
wire _16083_;
wire _16084_;
wire _16085_;
wire _16086_;
wire _16087_;
wire _16088_;
wire _16089_;
wire _16090_;
wire _16091_;
wire _16092_;
wire _16093_;
wire _16094_;
wire _16095_;
wire _16096_;
wire _16097_;
wire _16098_;
wire _16099_;
wire _16100_;
wire _16101_;
wire _16102_;
wire _16103_;
wire _16104_;
wire _16105_;
wire _16106_;
wire _16107_;
wire _16108_;
wire _16109_;
wire _16110_;
wire _16111_;
wire _16112_;
wire _16113_;
wire _16114_;
wire _16115_;
wire _16116_;
wire _16117_;
wire _16118_;
wire _16119_;
wire _16120_;
wire _16121_;
wire _16122_;
wire _16123_;
wire _16124_;
wire _16125_;
wire _16126_;
wire _16127_;
wire _16128_;
wire _16129_;
wire _16130_;
wire _16131_;
wire _16132_;
wire _16133_;
wire _16134_;
wire _16135_;
wire _16136_;
wire _16137_;
wire _16138_;
wire _16139_;
wire _16140_;
wire _16141_;
wire _16142_;
wire _16143_;
wire _16144_;
wire _16145_;
wire _16146_;
wire _16147_;
wire _16148_;
wire _16149_;
wire _16150_;
wire _16151_;
wire _16152_;
wire _16153_;
wire _16154_;
wire _16155_;
wire _16156_;
wire _16157_;
wire _16158_;
wire _16159_;
wire _16160_;
wire _16161_;
wire _16162_;
wire _16163_;
wire _16164_;
wire _16165_;
wire _16166_;
wire _16167_;
wire _16168_;
wire _16169_;
wire _16170_;
wire _16171_;
wire _16172_;
wire _16173_;
wire _16174_;
wire _16175_;
wire _16176_;
wire _16177_;
wire _16178_;
wire _16179_;
wire _16180_;
wire _16181_;
wire _16182_;
wire _16183_;
wire _16184_;
wire _16185_;
wire _16186_;
wire _16187_;
wire _16188_;
wire _16189_;
wire _16190_;
wire _16191_;
wire _16192_;
wire _16193_;
wire _16194_;
wire _16195_;
wire _16196_;
wire _16197_;
wire _16198_;
wire _16199_;
wire _16200_;
wire _16201_;
wire _16202_;
wire _16203_;
wire _16204_;
wire _16205_;
wire _16206_;
wire _16207_;
wire _16208_;
wire _16209_;
wire _16210_;
wire _16211_;
wire _16212_;
wire _16213_;
wire _16214_;
wire _16215_;
wire _16216_;
wire _16217_;
wire _16218_;
wire _16219_;
wire _16220_;
wire _16221_;
wire _16222_;
wire _16223_;
wire _16224_;
wire _16225_;
wire _16226_;
wire _16227_;
wire _16228_;
wire _16229_;
wire _16230_;
wire _16231_;
wire _16232_;
wire _16233_;
wire _16234_;
wire _16235_;
wire _16236_;
wire _16237_;
wire _16238_;
wire _16239_;
wire _16240_;
wire _16241_;
wire _16242_;
wire _16243_;
wire _16244_;
wire _16245_;
wire _16246_;
wire _16247_;
wire _16248_;
wire _16249_;
wire _16250_;
wire _16251_;
wire _16252_;
wire _16253_;
wire _16254_;
wire _16255_;
wire _16256_;
wire _16257_;
wire _16258_;
wire _16259_;
wire _16260_;
wire _16261_;
wire _16262_;
wire _16263_;
wire _16264_;
wire _16265_;
wire _16266_;
wire _16267_;
wire _16268_;
wire _16269_;
wire _16270_;
wire _16271_;
wire _16272_;
wire _16273_;
wire _16274_;
wire _16275_;
wire _16276_;
wire _16277_;
wire _16278_;
wire _16279_;
wire _16280_;
wire _16281_;
wire _16282_;
wire _16283_;
wire _16284_;
wire _16285_;
wire _16286_;
wire _16287_;
wire _16288_;
wire _16289_;
wire _16290_;
wire _16291_;
wire _16292_;
wire _16293_;
wire _16294_;
wire _16295_;
wire _16296_;
wire _16297_;
wire _16298_;
wire _16299_;
wire _16300_;
wire _16301_;
wire _16302_;
wire _16303_;
wire _16304_;
wire _16305_;
wire _16306_;
wire _16307_;
wire _16308_;
wire _16309_;
wire _16310_;
wire _16311_;
wire _16312_;
wire _16313_;
wire _16314_;
wire _16315_;
wire _16316_;
wire _16317_;
wire _16318_;
wire _16319_;
wire _16320_;
wire _16321_;
wire _16322_;
wire _16323_;
wire _16324_;
wire _16325_;
wire _16326_;
wire _16327_;
wire _16328_;
wire _16329_;
wire _16330_;
wire _16331_;
wire _16332_;
wire _16333_;
wire _16334_;
wire _16335_;
wire _16336_;
wire _16337_;
wire _16338_;
wire _16339_;
wire _16340_;
wire _16341_;
wire _16342_;
wire _16343_;
wire _16344_;
wire _16345_;
wire _16346_;
wire _16347_;
wire _16348_;
wire _16349_;
wire _16350_;
wire _16351_;
wire _16352_;
wire _16353_;
wire _16354_;
wire _16355_;
wire _16356_;
wire _16357_;
wire _16358_;
wire _16359_;
wire _16360_;
wire _16361_;
wire _16362_;
wire _16363_;
wire _16364_;
wire _16365_;
wire _16366_;
wire _16367_;
wire _16368_;
wire _16369_;
wire _16370_;
wire _16371_;
wire _16372_;
wire _16373_;
wire _16374_;
wire _16375_;
wire _16376_;
wire _16377_;
wire _16378_;
wire _16379_;
wire _16380_;
wire _16381_;
wire _16382_;
wire _16383_;
wire _16384_;
wire _16385_;
wire _16386_;
wire _16387_;
wire _16388_;
wire _16389_;
wire _16390_;
wire _16391_;
wire _16392_;
wire _16393_;
wire _16394_;
wire _16395_;
wire _16396_;
wire _16397_;
wire _16398_;
wire _16399_;
wire _16400_;
wire _16401_;
wire _16402_;
wire _16403_;
wire _16404_;
wire _16405_;
wire _16406_;
wire _16407_;
wire _16408_;
wire _16409_;
wire _16410_;
wire _16411_;
wire _16412_;
wire _16413_;
wire _16414_;
wire _16415_;
wire _16416_;
wire _16417_;
wire _16418_;
wire _16419_;
wire _16420_;
wire _16421_;
wire _16422_;
wire _16423_;
wire _16424_;
wire _16425_;
wire _16426_;
wire _16427_;
wire _16428_;
wire _16429_;
wire _16430_;
wire _16431_;
wire _16432_;
wire _16433_;
wire _16434_;
wire _16435_;
wire _16436_;
wire _16437_;
wire _16438_;
wire _16439_;
wire _16440_;
wire _16441_;
wire _16442_;
wire _16443_;
wire _16444_;
wire _16445_;
wire _16446_;
wire _16447_;
wire _16448_;
wire _16449_;
wire _16450_;
wire _16451_;
wire _16452_;
wire _16453_;
wire _16454_;
wire _16455_;
wire _16456_;
wire _16457_;
wire _16458_;
wire _16459_;
wire [31:0] alu_out;
wire [31:0] alu_out_q;
wire [63:0] cached_ascii_instr;
wire [31:0] cached_insn_imm;
wire [4:0] cached_insn_rd;
wire [4:0] cached_insn_rs1;
wire [4:0] cached_insn_rs2;
input clk;
wire clk;
wire [63:0] count_cycle;
wire [63:0] count_instr;
wire [7:0] cpu_state;
wire [31:0] cpuregs_0;
wire [31:0] cpuregs_10;
wire [31:0] cpuregs_11;
wire [31:0] cpuregs_12;
wire [31:0] cpuregs_13;
wire [31:0] cpuregs_14;
wire [31:0] cpuregs_15;
wire [31:0] cpuregs_16;
wire [31:0] cpuregs_17;
wire [31:0] cpuregs_18;
wire [31:0] cpuregs_19;
wire [31:0] cpuregs_1;
wire [31:0] cpuregs_20;
wire [31:0] cpuregs_21;
wire [31:0] cpuregs_22;
wire [31:0] cpuregs_23;
wire [31:0] cpuregs_24;
wire [31:0] cpuregs_25;
wire [31:0] cpuregs_26;
wire [31:0] cpuregs_27;
wire [31:0] cpuregs_28;
wire [31:0] cpuregs_29;
wire [31:0] cpuregs_2;
wire [31:0] cpuregs_30;
wire [31:0] cpuregs_31;
wire [31:0] cpuregs_3;
wire [31:0] cpuregs_4;
wire [31:0] cpuregs_5;
wire [31:0] cpuregs_6;
wire [31:0] cpuregs_7;
wire [31:0] cpuregs_8;
wire [31:0] cpuregs_9;
wire [63:0] dbg_ascii_instr;
wire [127:0] dbg_ascii_state;
wire [31:0] dbg_insn_imm;
wire [4:0] dbg_insn_rd;
wire [4:0] dbg_insn_rs1;
wire [4:0] dbg_insn_rs2;
wire dbg_next;
wire [31:0] dbg_rs1val;
wire dbg_rs1val_valid;
wire [31:0] dbg_rs2val;
wire dbg_rs2val_valid;
wire [31:0] decoded_imm;
wire [31:0] decoded_imm_j;
wire [4:0] decoded_rd;
wire decoder_pseudo_trigger;
wire decoder_pseudo_trigger_q;
wire decoder_trigger;
wire decoder_trigger_q;
output [31:0] eoi;
wire [31:0] eoi;
wire instr_add;
wire instr_addi;
wire instr_and;
wire instr_andi;
wire instr_auipc;
wire instr_beq;
wire instr_bge;
wire instr_bgeu;
wire instr_blt;
wire instr_bltu;
wire instr_bne;
wire instr_jal;
wire instr_jalr;
wire instr_lb;
wire instr_lbu;
wire instr_lh;
wire instr_lhu;
wire instr_lui;
wire instr_lw;
wire instr_or;
wire instr_ori;
wire instr_rdcycle;
wire instr_rdcycleh;
wire instr_rdinstr;
wire instr_rdinstrh;
wire instr_sb;
wire instr_sh;
wire instr_sll;
wire instr_slli;
wire instr_slt;
wire instr_slti;
wire instr_sltiu;
wire instr_sltu;
wire instr_sra;
wire instr_srai;
wire instr_srl;
wire instr_srli;
wire instr_sub;
wire instr_sw;
wire instr_xor;
wire instr_xori;
input [31:0] irq;
wire [31:0] irq;
wire is_alu_reg_imm;
wire is_alu_reg_reg;
wire is_beq_bne_blt_bge_bltu_bgeu;
wire is_compare;
wire is_jalr_addi_slti_sltiu_xori_ori_andi;
wire is_lb_lh_lw_lbu_lhu;
wire is_lbu_lhu_lw;
wire is_lui_auipc_jal;
wire is_lui_auipc_jal_jalr_addi_add_sub;
wire is_sb_sh_sw;
wire is_sll_srl_sra;
wire is_slli_srli_srai;
wire is_slti_blt_slt;
wire is_sltiu_bltu_sltu;
wire latched_branch;
wire latched_is_lb;
wire latched_is_lh;
wire latched_is_lu;
wire [4:0] latched_rd;
wire latched_stalu;
wire latched_store;
wire launch_next_insn;
output [31:0] mem_addr;
wire [31:0] mem_addr;
wire mem_do_prefetch;
wire mem_do_rdata;
wire mem_do_rinst;
wire mem_do_wdata;
output mem_instr;
wire mem_instr;
output [31:0] mem_la_addr;
wire [31:0] mem_la_addr;
output mem_la_read;
wire mem_la_read;
output [31:0] mem_la_wdata;
wire [31:0] mem_la_wdata;
output mem_la_write;
wire mem_la_write;
output [3:0] mem_la_wstrb;
wire [3:0] mem_la_wstrb;
input [31:0] mem_rdata;
wire [31:0] mem_rdata;
wire [31:0] mem_rdata_q;
input mem_ready;
wire mem_ready;
wire [1:0] mem_state;
output mem_valid;
wire mem_valid;
output [31:0] mem_wdata;
wire [31:0] mem_wdata;
wire [1:0] mem_wordsize;
output [3:0] mem_wstrb;
wire [3:0] mem_wstrb;
output [31:0] pcpi_insn;
wire [31:0] pcpi_insn;
input [31:0] pcpi_rd;
wire [31:0] pcpi_rd;
input pcpi_ready;
wire pcpi_ready;
output [31:0] pcpi_rs1;
wire [31:0] pcpi_rs1;
output [31:0] pcpi_rs2;
wire [31:0] pcpi_rs2;
output pcpi_valid;
wire pcpi_valid;
input pcpi_wait;
wire pcpi_wait;
input pcpi_wr;
wire pcpi_wr;
wire [63:0] q_ascii_instr;
wire [31:0] q_insn_imm;
wire [4:0] q_insn_rd;
wire [4:0] q_insn_rs1;
wire [4:0] q_insn_rs2;
wire [31:0] reg_next_pc;
wire [31:0] reg_out;
wire [31:0] reg_pc;
wire [4:0] reg_sh;
input resetn;
wire resetn;
output [35:0] trace_data;
wire [35:0] trace_data;
output trace_valid;
wire trace_valid;
output trap;
wire trap;
NOT_g _16460_ (.A(count_instr[62]), .Y(_10854_));
NOT_g _16461_ (.A(count_instr[60]), .Y(_10855_));
NOT_g _16462_ (.A(count_instr[58]), .Y(_10856_));
NOT_g _16463_ (.A(count_instr[56]), .Y(_10857_));
NOT_g _16464_ (.A(count_instr[54]), .Y(_10858_));
NOT_g _16465_ (.A(count_instr[53]), .Y(_10859_));
NOT_g _16466_ (.A(count_instr[51]), .Y(_10860_));
NOT_g _16467_ (.A(count_instr[50]), .Y(_10861_));
NOT_g _16468_ (.A(count_instr[46]), .Y(_10862_));
NOT_g _16469_ (.A(count_instr[45]), .Y(_10863_));
NOT_g _16470_ (.A(count_instr[44]), .Y(_10864_));
NOT_g _16471_ (.A(count_instr[43]), .Y(_10865_));
NOT_g _16472_ (.A(count_instr[41]), .Y(_10866_));
NOT_g _16473_ (.A(count_instr[38]), .Y(_10867_));
NOT_g _16474_ (.A(count_instr[37]), .Y(_10868_));
NOT_g _16475_ (.A(count_instr[35]), .Y(_10869_));
NOT_g _16476_ (.A(count_instr[34]), .Y(_10870_));
NOT_g _16477_ (.A(count_instr[33]), .Y(_10871_));
NOT_g _16478_ (.A(count_instr[31]), .Y(_10872_));
NOT_g _16479_ (.A(count_instr[30]), .Y(_10873_));
NOT_g _16480_ (.A(count_instr[29]), .Y(_10874_));
NOT_g _16481_ (.A(count_instr[27]), .Y(_10875_));
NOT_g _16482_ (.A(count_instr[26]), .Y(_10876_));
NOT_g _16483_ (.A(count_instr[24]), .Y(_10877_));
NOT_g _16484_ (.A(count_instr[23]), .Y(_10878_));
NOT_g _16485_ (.A(count_instr[22]), .Y(_10879_));
NOT_g _16486_ (.A(count_instr[21]), .Y(_10880_));
NOT_g _16487_ (.A(count_instr[20]), .Y(_10881_));
NOT_g _16488_ (.A(count_instr[18]), .Y(_10882_));
NOT_g _16489_ (.A(count_instr[16]), .Y(_10883_));
NOT_g _16490_ (.A(count_instr[15]), .Y(_10884_));
NOT_g _16491_ (.A(count_instr[12]), .Y(_10885_));
NOT_g _16492_ (.A(count_instr[11]), .Y(_10886_));
NOT_g _16493_ (.A(count_instr[9]), .Y(_10887_));
NOT_g _16494_ (.A(count_instr[7]), .Y(_10888_));
NOT_g _16495_ (.A(count_instr[6]), .Y(_10889_));
NOT_g _16496_ (.A(count_instr[5]), .Y(_10890_));
NOT_g _16497_ (.A(count_instr[3]), .Y(_10891_));
NOT_g _16498_ (.A(count_instr[1]), .Y(_10892_));
NOT_g _16499_ (.A(mem_do_wdata), .Y(_10893_));
NOT_g _16500_ (.A(latched_is_lh), .Y(_10894_));
NOT_g _16501_ (.A(latched_is_lu), .Y(_10895_));
NOT_g _16502_ (.A(latched_branch), .Y(_10896_));
NOT_g _16503_ (.A(latched_stalu), .Y(_10897_));
NOT_g _16504_ (.A(mem_do_rinst), .Y(_10898_));
NOT_g _16505_ (.A(reg_pc[31]), .Y(_10899_));
NOT_g _16506_ (.A(reg_pc[2]), .Y(_10900_));
NOT_g _16507_ (.A(mem_do_prefetch), .Y(_10901_));
NOT_g _16508_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .Y(_10902_));
NOT_g _16509_ (.A(instr_and), .Y(_10903_));
NOT_g _16510_ (.A(instr_or), .Y(_10904_));
NOT_g _16511_ (.A(instr_sra), .Y(_10905_));
NOT_g _16512_ (.A(instr_srl), .Y(_10906_));
NOT_g _16513_ (.A(instr_xor), .Y(_10907_));
NOT_g _16514_ (.A(instr_sltu), .Y(_10908_));
NOT_g _16515_ (.A(instr_sll), .Y(_10909_));
NOT_g _16516_ (.A(instr_sub), .Y(_10910_));
NOT_g _16517_ (.A(instr_add), .Y(_10911_));
NOT_g _16518_ (.A(instr_andi), .Y(_10912_));
NOT_g _16519_ (.A(instr_ori), .Y(_10913_));
NOT_g _16520_ (.A(instr_xori), .Y(_10914_));
NOT_g _16521_ (.A(instr_sltiu), .Y(_10915_));
NOT_g _16522_ (.A(instr_slti), .Y(_10916_));
NOT_g _16523_ (.A(instr_addi), .Y(_10917_));
NOT_g _16524_ (.A(instr_bgeu), .Y(_10918_));
NOT_g _16525_ (.A(instr_bltu), .Y(_10919_));
NOT_g _16526_ (.A(instr_bge), .Y(_10920_));
NOT_g _16527_ (.A(instr_blt), .Y(_10921_));
NOT_g _16528_ (.A(cpuregs_29[0]), .Y(_10922_));
NOT_g _16529_ (.A(cpuregs_29[4]), .Y(_10923_));
NOT_g _16530_ (.A(cpuregs_29[5]), .Y(_10924_));
NOT_g _16531_ (.A(cpuregs_29[6]), .Y(_10925_));
NOT_g _16532_ (.A(cpuregs_29[8]), .Y(_10926_));
NOT_g _16533_ (.A(cpuregs_29[12]), .Y(_10927_));
NOT_g _16534_ (.A(cpuregs_29[13]), .Y(_10928_));
NOT_g _16535_ (.A(cpuregs_29[15]), .Y(_10929_));
NOT_g _16536_ (.A(cpuregs_29[17]), .Y(_10930_));
NOT_g _16537_ (.A(cpuregs_29[18]), .Y(_10931_));
NOT_g _16538_ (.A(cpuregs_29[20]), .Y(_10932_));
NOT_g _16539_ (.A(cpuregs_29[29]), .Y(_10933_));
NOT_g _16540_ (.A(cpuregs_9[19]), .Y(_10934_));
NOT_g _16541_ (.A(cpuregs_9[25]), .Y(_10935_));
NOT_g _16542_ (.A(cpuregs_9[27]), .Y(_10936_));
NOT_g _16543_ (.A(cpuregs_6[2]), .Y(_10937_));
NOT_g _16544_ (.A(cpuregs_6[3]), .Y(_10938_));
NOT_g _16545_ (.A(cpuregs_6[6]), .Y(_10939_));
NOT_g _16546_ (.A(cpuregs_6[7]), .Y(_10940_));
NOT_g _16547_ (.A(cpuregs_6[10]), .Y(_10941_));
NOT_g _16548_ (.A(cpuregs_6[11]), .Y(_10942_));
NOT_g _16549_ (.A(cpuregs_6[14]), .Y(_10943_));
NOT_g _16550_ (.A(cpuregs_6[18]), .Y(_10944_));
NOT_g _16551_ (.A(cpuregs_6[20]), .Y(_10945_));
NOT_g _16552_ (.A(cpuregs_6[22]), .Y(_10946_));
NOT_g _16553_ (.A(cpuregs_6[23]), .Y(_10947_));
NOT_g _16554_ (.A(cpuregs_6[30]), .Y(_10948_));
NOT_g _16555_ (.A(cpuregs_4[2]), .Y(_10949_));
NOT_g _16556_ (.A(cpuregs_4[3]), .Y(_10950_));
NOT_g _16557_ (.A(cpuregs_4[6]), .Y(_10951_));
NOT_g _16558_ (.A(cpuregs_4[7]), .Y(_10952_));
NOT_g _16559_ (.A(cpuregs_4[10]), .Y(_10953_));
NOT_g _16560_ (.A(cpuregs_4[11]), .Y(_10954_));
NOT_g _16561_ (.A(cpuregs_4[14]), .Y(_10955_));
NOT_g _16562_ (.A(cpuregs_4[18]), .Y(_10956_));
NOT_g _16563_ (.A(cpuregs_4[20]), .Y(_10957_));
NOT_g _16564_ (.A(cpuregs_4[22]), .Y(_10958_));
NOT_g _16565_ (.A(cpuregs_4[23]), .Y(_10959_));
NOT_g _16566_ (.A(cpuregs_4[30]), .Y(_10960_));
NOT_g _16567_ (.A(instr_auipc), .Y(_10961_));
NOT_g _16568_ (.A(instr_jal), .Y(_10962_));
NOT_g _16569_ (.A(resetn), .Y(_10963_));
NOT_g _16570_ (.A(is_sll_srl_sra), .Y(_10964_));
NOT_g _16571_ (.A(instr_lw), .Y(_10965_));
NOT_g _16572_ (.A(instr_sb), .Y(_10966_));
NOT_g _16573_ (.A(instr_sh), .Y(_10967_));
NOT_g _16574_ (.A(instr_sw), .Y(_10968_));
NOT_g _16575_ (.A(instr_slli), .Y(_10969_));
NOT_g _16576_ (.A(instr_srli), .Y(_10970_));
NOT_g _16577_ (.A(instr_srai), .Y(_10971_));
NOT_g _16578_ (.A(instr_rdcycle), .Y(_10972_));
NOT_g _16579_ (.A(instr_rdcycleh), .Y(_10973_));
NOT_g _16580_ (.A(instr_rdinstr), .Y(_10974_));
NOT_g _16581_ (.A(instr_rdinstrh), .Y(_10975_));
NOT_g _16582_ (.A(decoded_imm_j[3]), .Y(_10976_));
NOT_g _16583_ (.A(is_slli_srli_srai), .Y(_10977_));
NOT_g _16584_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi), .Y(_10978_));
NOT_g _16585_ (.A(instr_lui), .Y(_10979_));
NOT_g _16586_ (.A(is_sb_sh_sw), .Y(_10980_));
NOT_g _16587_ (.A(is_alu_reg_imm), .Y(_10981_));
NOT_g _16588_ (.A(pcpi_rs2[1]), .Y(_10982_));
NOT_g _16589_ (.A(pcpi_rs2[2]), .Y(_10983_));
NOT_g _16590_ (.A(pcpi_rs2[4]), .Y(_10984_));
NOT_g _16591_ (.A(pcpi_rs2[5]), .Y(_10985_));
NOT_g _16592_ (.A(pcpi_rs2[6]), .Y(_10986_));
NOT_g _16593_ (.A(pcpi_rs2[7]), .Y(_10987_));
NOT_g _16594_ (.A(pcpi_rs2[8]), .Y(_10988_));
NOT_g _16595_ (.A(pcpi_rs2[9]), .Y(_10989_));
NOT_g _16596_ (.A(pcpi_rs2[10]), .Y(_10990_));
NOT_g _16597_ (.A(pcpi_rs2[11]), .Y(_10991_));
NOT_g _16598_ (.A(pcpi_rs2[12]), .Y(_10992_));
NOT_g _16599_ (.A(pcpi_rs2[13]), .Y(_10993_));
NOT_g _16600_ (.A(pcpi_rs2[14]), .Y(_10994_));
NOT_g _16601_ (.A(pcpi_rs2[15]), .Y(_10995_));
NOT_g _16602_ (.A(pcpi_rs2[16]), .Y(_10996_));
NOT_g _16603_ (.A(pcpi_rs2[17]), .Y(_10997_));
NOT_g _16604_ (.A(pcpi_rs2[18]), .Y(_10998_));
NOT_g _16605_ (.A(pcpi_rs2[19]), .Y(_10999_));
NOT_g _16606_ (.A(pcpi_rs2[20]), .Y(_11000_));
NOT_g _16607_ (.A(pcpi_rs2[21]), .Y(_11001_));
NOT_g _16608_ (.A(pcpi_rs2[22]), .Y(_11002_));
NOT_g _16609_ (.A(pcpi_rs2[23]), .Y(_11003_));
NOT_g _16610_ (.A(pcpi_rs2[24]), .Y(_11004_));
NOT_g _16611_ (.A(pcpi_rs2[25]), .Y(_11005_));
NOT_g _16612_ (.A(pcpi_rs2[26]), .Y(_11006_));
NOT_g _16613_ (.A(pcpi_rs2[27]), .Y(_11007_));
NOT_g _16614_ (.A(pcpi_rs2[28]), .Y(_11008_));
NOT_g _16615_ (.A(pcpi_rs2[29]), .Y(_11009_));
NOT_g _16616_ (.A(pcpi_rs2[30]), .Y(_11010_));
NOT_g _16617_ (.A(pcpi_rs2[31]), .Y(_11011_));
NOT_g _16618_ (.A(mem_wordsize[0]), .Y(_11012_));
NOT_g _16619_ (.A(mem_wordsize[1]), .Y(_11013_));
NOT_g _16620_ (.A(cpuregs_22[1]), .Y(_11014_));
NOT_g _16621_ (.A(cpuregs_22[10]), .Y(_11015_));
NOT_g _16622_ (.A(cpuregs_22[11]), .Y(_11016_));
NOT_g _16623_ (.A(cpuregs_22[17]), .Y(_11017_));
NOT_g _16624_ (.A(cpuregs_22[18]), .Y(_11018_));
NOT_g _16625_ (.A(cpuregs_22[21]), .Y(_11019_));
NOT_g _16626_ (.A(cpuregs_22[26]), .Y(_11020_));
NOT_g _16627_ (.A(cpuregs_22[29]), .Y(_11021_));
NOT_g _16628_ (.A(cpuregs_21[1]), .Y(_11022_));
NOT_g _16629_ (.A(cpuregs_21[2]), .Y(_11023_));
NOT_g _16630_ (.A(cpuregs_21[5]), .Y(_11024_));
NOT_g _16631_ (.A(cpuregs_21[6]), .Y(_11025_));
NOT_g _16632_ (.A(cpuregs_21[10]), .Y(_11026_));
NOT_g _16633_ (.A(cpuregs_21[11]), .Y(_11027_));
NOT_g _16634_ (.A(cpuregs_21[12]), .Y(_11028_));
NOT_g _16635_ (.A(cpuregs_21[14]), .Y(_11029_));
NOT_g _16636_ (.A(cpuregs_21[15]), .Y(_11030_));
NOT_g _16637_ (.A(cpuregs_21[17]), .Y(_11031_));
NOT_g _16638_ (.A(cpuregs_21[18]), .Y(_11032_));
NOT_g _16639_ (.A(cpuregs_21[21]), .Y(_11033_));
NOT_g _16640_ (.A(cpuregs_21[22]), .Y(_11034_));
NOT_g _16641_ (.A(cpuregs_21[25]), .Y(_11035_));
NOT_g _16642_ (.A(cpuregs_21[26]), .Y(_11036_));
NOT_g _16643_ (.A(cpuregs_21[29]), .Y(_11037_));
NOT_g _16644_ (.A(cpuregs_21[30]), .Y(_11038_));
NOT_g _16645_ (.A(cpuregs_21[31]), .Y(_11039_));
NOT_g _16646_ (.A(dbg_next), .Y(_11040_));
NOT_g _16647_ (.A(latched_rd[0]), .Y(_11041_));
NOT_g _16648_ (.A(latched_rd[2]), .Y(_11042_));
NOT_g _16649_ (.A(latched_rd[3]), .Y(_11043_));
NOT_g _16650_ (.A(latched_rd[4]), .Y(_11044_));
NOT_g _16651_ (.A(decoder_trigger_q), .Y(_11045_));
NOT_g _16652_ (.A(decoded_imm_j[15]), .Y(_11046_));
NOT_g _16653_ (.A(decoded_imm_j[17]), .Y(_11047_));
NOT_g _16654_ (.A(decoded_imm_j[19]), .Y(_11048_));
NOT_g _16655_ (.A(decoded_imm_j[4]), .Y(_11049_));
NOT_g _16656_ (.A(cached_ascii_instr[0]), .Y(_11050_));
NOT_g _16657_ (.A(cached_ascii_instr[1]), .Y(_11051_));
NOT_g _16658_ (.A(cached_ascii_instr[2]), .Y(_11052_));
NOT_g _16659_ (.A(cached_ascii_instr[3]), .Y(_11053_));
NOT_g _16660_ (.A(cached_ascii_instr[4]), .Y(_11054_));
NOT_g _16661_ (.A(cached_ascii_instr[8]), .Y(_11055_));
NOT_g _16662_ (.A(cached_ascii_instr[9]), .Y(_11056_));
NOT_g _16663_ (.A(cached_ascii_instr[10]), .Y(_11057_));
NOT_g _16664_ (.A(cached_ascii_instr[11]), .Y(_11058_));
NOT_g _16665_ (.A(cached_ascii_instr[12]), .Y(_11059_));
NOT_g _16666_ (.A(cached_ascii_instr[16]), .Y(_11060_));
NOT_g _16667_ (.A(cached_ascii_instr[17]), .Y(_11061_));
NOT_g _16668_ (.A(cached_ascii_instr[18]), .Y(_11062_));
NOT_g _16669_ (.A(cached_ascii_instr[19]), .Y(_11063_));
NOT_g _16670_ (.A(cached_ascii_instr[20]), .Y(_11064_));
NOT_g _16671_ (.A(cached_ascii_instr[22]), .Y(_11065_));
NOT_g _16672_ (.A(cached_ascii_instr[24]), .Y(_11066_));
NOT_g _16673_ (.A(cached_ascii_instr[25]), .Y(_11067_));
NOT_g _16674_ (.A(cached_ascii_instr[26]), .Y(_11068_));
NOT_g _16675_ (.A(cached_ascii_instr[27]), .Y(_11069_));
NOT_g _16676_ (.A(cached_ascii_instr[28]), .Y(_11070_));
NOT_g _16677_ (.A(cached_ascii_instr[30]), .Y(_11071_));
NOT_g _16678_ (.A(cached_ascii_instr[32]), .Y(_11072_));
NOT_g _16679_ (.A(cached_ascii_instr[33]), .Y(_11073_));
NOT_g _16680_ (.A(cached_ascii_instr[35]), .Y(_11074_));
NOT_g _16681_ (.A(cached_ascii_instr[36]), .Y(_11075_));
NOT_g _16682_ (.A(cached_ascii_instr[38]), .Y(_11076_));
NOT_g _16683_ (.A(mem_rdata_q[12]), .Y(_11077_));
NOT_g _16684_ (.A(mem_rdata_q[13]), .Y(_11078_));
NOT_g _16685_ (.A(mem_rdata_q[14]), .Y(_11079_));
NOT_g _16686_ (.A(mem_rdata_q[20]), .Y(_11080_));
NOT_g _16687_ (.A(mem_rdata_q[27]), .Y(_11081_));
NOT_g _16688_ (.A(mem_rdata_q[29]), .Y(_11082_));
NOT_g _16689_ (.A(mem_rdata_q[31]), .Y(_11083_));
NOT_g _16690_ (.A(mem_state[1]), .Y(_11084_));
NOT_g _16691_ (.A(mem_rdata_q[2]), .Y(_11085_));
NOT_g _16692_ (.A(mem_rdata_q[3]), .Y(_11086_));
NOT_g _16693_ (.A(cpuregs_31[0]), .Y(_11087_));
NOT_g _16694_ (.A(cpuregs_31[4]), .Y(_11088_));
NOT_g _16695_ (.A(cpuregs_31[8]), .Y(_11089_));
NOT_g _16696_ (.A(cpuregs_31[13]), .Y(_11090_));
NOT_g _16697_ (.A(cpuregs_31[18]), .Y(_11091_));
NOT_g _16698_ (.A(cpuregs_31[20]), .Y(_11092_));
NOT_g _16699_ (.A(cpuregs_28[0]), .Y(_11093_));
NOT_g _16700_ (.A(cpuregs_28[4]), .Y(_11094_));
NOT_g _16701_ (.A(cpuregs_28[6]), .Y(_11095_));
NOT_g _16702_ (.A(cpuregs_28[8]), .Y(_11096_));
NOT_g _16703_ (.A(cpuregs_28[13]), .Y(_11097_));
NOT_g _16704_ (.A(cpuregs_28[17]), .Y(_11098_));
NOT_g _16705_ (.A(cpuregs_28[18]), .Y(_11099_));
NOT_g _16706_ (.A(cpuregs_28[20]), .Y(_11100_));
NOT_g _16707_ (.A(cpuregs_28[29]), .Y(_11101_));
NOT_g _16708_ (.A(cpuregs_14[8]), .Y(_11102_));
NOT_g _16709_ (.A(cpuregs_14[16]), .Y(_11103_));
NOT_g _16710_ (.A(cpuregs_14[18]), .Y(_11104_));
NOT_g _16711_ (.A(cpuregs_14[19]), .Y(_11105_));
NOT_g _16712_ (.A(cpuregs_14[27]), .Y(_11106_));
NOT_g _16713_ (.A(cpuregs_5[2]), .Y(_11107_));
NOT_g _16714_ (.A(cpuregs_5[3]), .Y(_11108_));
NOT_g _16715_ (.A(cpuregs_5[6]), .Y(_11109_));
NOT_g _16716_ (.A(cpuregs_5[7]), .Y(_11110_));
NOT_g _16717_ (.A(cpuregs_5[10]), .Y(_11111_));
NOT_g _16718_ (.A(cpuregs_5[11]), .Y(_11112_));
NOT_g _16719_ (.A(cpuregs_5[14]), .Y(_11113_));
NOT_g _16720_ (.A(cpuregs_5[18]), .Y(_11114_));
NOT_g _16721_ (.A(cpuregs_5[20]), .Y(_11115_));
NOT_g _16722_ (.A(cpuregs_5[22]), .Y(_11116_));
NOT_g _16723_ (.A(cpuregs_5[23]), .Y(_11117_));
NOT_g _16724_ (.A(cpuregs_5[30]), .Y(_11118_));
NOT_g _16725_ (.A(cpuregs_12[15]), .Y(_11119_));
NOT_g _16726_ (.A(cpuregs_12[18]), .Y(_11120_));
NOT_g _16727_ (.A(cpuregs_12[19]), .Y(_11121_));
NOT_g _16728_ (.A(cpuregs_12[27]), .Y(_11122_));
NOT_g _16729_ (.A(cpuregs_7[2]), .Y(_11123_));
NOT_g _16730_ (.A(cpuregs_7[3]), .Y(_11124_));
NOT_g _16731_ (.A(cpuregs_7[6]), .Y(_11125_));
NOT_g _16732_ (.A(cpuregs_7[7]), .Y(_11126_));
NOT_g _16733_ (.A(cpuregs_7[10]), .Y(_11127_));
NOT_g _16734_ (.A(cpuregs_7[11]), .Y(_11128_));
NOT_g _16735_ (.A(cpuregs_7[14]), .Y(_11129_));
NOT_g _16736_ (.A(cpuregs_7[18]), .Y(_11130_));
NOT_g _16737_ (.A(cpuregs_7[20]), .Y(_11131_));
NOT_g _16738_ (.A(cpuregs_7[22]), .Y(_11132_));
NOT_g _16739_ (.A(cpuregs_7[23]), .Y(_11133_));
NOT_g _16740_ (.A(cpuregs_7[30]), .Y(_11134_));
NOT_g _16741_ (.A(pcpi_rs1[0]), .Y(_11135_));
NOT_g _16742_ (.A(pcpi_rs1[1]), .Y(_11136_));
NOT_g _16743_ (.A(decoded_imm_j[7]), .Y(_11137_));
NOT_g _16744_ (.A(decoded_imm_j[31]), .Y(_11138_));
NOT_g _16745_ (.A(cpuregs_13[0]), .Y(_11139_));
NOT_g _16746_ (.A(cpuregs_13[1]), .Y(_11140_));
NOT_g _16747_ (.A(cpuregs_13[4]), .Y(_11141_));
NOT_g _16748_ (.A(cpuregs_13[5]), .Y(_11142_));
NOT_g _16749_ (.A(cpuregs_13[6]), .Y(_11143_));
NOT_g _16750_ (.A(cpuregs_13[8]), .Y(_11144_));
NOT_g _16751_ (.A(cpuregs_13[9]), .Y(_11145_));
NOT_g _16752_ (.A(cpuregs_13[12]), .Y(_11146_));
NOT_g _16753_ (.A(cpuregs_13[13]), .Y(_11147_));
NOT_g _16754_ (.A(cpuregs_13[15]), .Y(_11148_));
NOT_g _16755_ (.A(cpuregs_13[17]), .Y(_11149_));
NOT_g _16756_ (.A(cpuregs_13[18]), .Y(_11150_));
NOT_g _16757_ (.A(cpuregs_13[19]), .Y(_11151_));
NOT_g _16758_ (.A(cpuregs_13[20]), .Y(_11152_));
NOT_g _16759_ (.A(cpuregs_13[25]), .Y(_11153_));
NOT_g _16760_ (.A(cpuregs_13[27]), .Y(_11154_));
NOT_g _16761_ (.A(decoded_imm_j[13]), .Y(_11155_));
NOT_g _16762_ (.A(cpuregs_15[0]), .Y(_11156_));
NOT_g _16763_ (.A(cpuregs_15[1]), .Y(_11157_));
NOT_g _16764_ (.A(cpuregs_15[4]), .Y(_11158_));
NOT_g _16765_ (.A(cpuregs_15[8]), .Y(_11159_));
NOT_g _16766_ (.A(cpuregs_15[9]), .Y(_11160_));
NOT_g _16767_ (.A(cpuregs_15[12]), .Y(_11161_));
NOT_g _16768_ (.A(cpuregs_15[13]), .Y(_11162_));
NOT_g _16769_ (.A(cpuregs_15[15]), .Y(_11163_));
NOT_g _16770_ (.A(cpuregs_15[16]), .Y(_11164_));
NOT_g _16771_ (.A(cpuregs_15[17]), .Y(_11165_));
NOT_g _16772_ (.A(cpuregs_15[18]), .Y(_11166_));
NOT_g _16773_ (.A(cpuregs_15[19]), .Y(_11167_));
NOT_g _16774_ (.A(cpuregs_15[20]), .Y(_11168_));
NOT_g _16775_ (.A(cpuregs_15[25]), .Y(_11169_));
NOT_g _16776_ (.A(cpuregs_15[27]), .Y(_11170_));
NOT_g _16777_ (.A(cpuregs_30[0]), .Y(_11171_));
NOT_g _16778_ (.A(cpuregs_30[4]), .Y(_11172_));
NOT_g _16779_ (.A(cpuregs_30[8]), .Y(_11173_));
NOT_g _16780_ (.A(cpuregs_30[13]), .Y(_11174_));
NOT_g _16781_ (.A(cpuregs_30[18]), .Y(_11175_));
NOT_g _16782_ (.A(cpuregs_30[20]), .Y(_11176_));
NOT_g _16783_ (.A(cpuregs_23[1]), .Y(_11177_));
NOT_g _16784_ (.A(cpuregs_23[2]), .Y(_11178_));
NOT_g _16785_ (.A(cpuregs_23[6]), .Y(_11179_));
NOT_g _16786_ (.A(cpuregs_23[10]), .Y(_11180_));
NOT_g _16787_ (.A(cpuregs_23[11]), .Y(_11181_));
NOT_g _16788_ (.A(cpuregs_23[12]), .Y(_11182_));
NOT_g _16789_ (.A(cpuregs_23[14]), .Y(_11183_));
NOT_g _16790_ (.A(cpuregs_23[17]), .Y(_11184_));
NOT_g _16791_ (.A(cpuregs_23[18]), .Y(_11185_));
NOT_g _16792_ (.A(cpuregs_23[21]), .Y(_11186_));
NOT_g _16793_ (.A(cpuregs_23[22]), .Y(_11187_));
NOT_g _16794_ (.A(cpuregs_23[25]), .Y(_11188_));
NOT_g _16795_ (.A(cpuregs_23[26]), .Y(_11189_));
NOT_g _16796_ (.A(cpuregs_23[29]), .Y(_11190_));
NOT_g _16797_ (.A(cpuregs_23[30]), .Y(_11191_));
NOT_g _16798_ (.A(cpuregs_23[31]), .Y(_11192_));
NOT_g _16799_ (.A(cpuregs_20[1]), .Y(_11193_));
NOT_g _16800_ (.A(cpuregs_20[6]), .Y(_11194_));
NOT_g _16801_ (.A(cpuregs_20[10]), .Y(_11195_));
NOT_g _16802_ (.A(cpuregs_20[11]), .Y(_11196_));
NOT_g _16803_ (.A(cpuregs_20[12]), .Y(_11197_));
NOT_g _16804_ (.A(cpuregs_20[17]), .Y(_11198_));
NOT_g _16805_ (.A(cpuregs_20[18]), .Y(_11199_));
NOT_g _16806_ (.A(cpuregs_20[21]), .Y(_11200_));
NOT_g _16807_ (.A(cpuregs_20[26]), .Y(_11201_));
NOT_g _16808_ (.A(cpuregs_20[29]), .Y(_11202_));
NOT_g _16809_ (.A(cpu_state[7]), .Y(_11203_));
NOT_g _16810_ (.A(cpu_state[4]), .Y(_11204_));
NOT_g _16811_ (.A(cpu_state[3]), .Y(_11205_));
NOT_g _16812_ (.A(cpu_state[0]), .Y(_11206_));
NOT_g _16813_ (.A(reg_sh[0]), .Y(_11207_));
NOT_g _16814_ (.A(reg_sh[4]), .Y(_11208_));
NOT_g _16815_ (.A(is_lui_auipc_jal), .Y(_11209_));
NOT_g _16816_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(_11210_));
NOT_g _16817_ (.A(decoder_pseudo_trigger), .Y(_11211_));
NOT_g _16818_ (.A(_00012_[0]), .Y(_11212_));
NOT_g _16819_ (.A(_00012_[1]), .Y(_11213_));
NOT_g _16820_ (.A(_00012_[2]), .Y(_11214_));
NOT_g _16821_ (.A(_00012_[3]), .Y(_11215_));
NOT_g _16822_ (.A(_00012_[4]), .Y(_11216_));
NOT_g _16823_ (.A(_00011_[0]), .Y(_11217_));
NOT_g _16824_ (.A(_00011_[1]), .Y(_11218_));
NOT_g _16825_ (.A(_00011_[2]), .Y(_11219_));
NOT_g _16826_ (.A(_00011_[3]), .Y(_11220_));
NOT_g _16827_ (.A(_00011_[4]), .Y(_11221_));
NOT_g _16828_ (.A(alu_out_q[0]), .Y(_11222_));
NOT_g _16829_ (.A(decoder_pseudo_trigger_q), .Y(_11223_));
NOT_g _16830_ (.A(count_cycle[2]), .Y(_11224_));
NOT_g _16831_ (.A(count_cycle[4]), .Y(_11225_));
NOT_g _16832_ (.A(count_cycle[6]), .Y(_11226_));
NOT_g _16833_ (.A(count_cycle[8]), .Y(_11227_));
NOT_g _16834_ (.A(count_cycle[10]), .Y(_11228_));
NOT_g _16835_ (.A(count_cycle[12]), .Y(_11229_));
NOT_g _16836_ (.A(count_cycle[14]), .Y(_11230_));
NOT_g _16837_ (.A(count_cycle[16]), .Y(_11231_));
NOT_g _16838_ (.A(count_cycle[18]), .Y(_11232_));
NOT_g _16839_ (.A(count_cycle[20]), .Y(_11233_));
NOT_g _16840_ (.A(count_cycle[22]), .Y(_11234_));
NOT_g _16841_ (.A(count_cycle[24]), .Y(_11235_));
NOT_g _16842_ (.A(count_cycle[26]), .Y(_11236_));
NOT_g _16843_ (.A(count_cycle[28]), .Y(_11237_));
NOT_g _16844_ (.A(count_cycle[30]), .Y(_11238_));
NOT_g _16845_ (.A(count_cycle[32]), .Y(_11239_));
NOT_g _16846_ (.A(count_cycle[34]), .Y(_11240_));
NOT_g _16847_ (.A(count_cycle[36]), .Y(_11241_));
NOT_g _16848_ (.A(count_cycle[38]), .Y(_11242_));
NOT_g _16849_ (.A(count_cycle[40]), .Y(_11243_));
NOT_g _16850_ (.A(count_cycle[42]), .Y(_11244_));
NOT_g _16851_ (.A(count_cycle[44]), .Y(_11245_));
NOT_g _16852_ (.A(count_cycle[46]), .Y(_11246_));
NOT_g _16853_ (.A(count_cycle[48]), .Y(_11247_));
NOT_g _16854_ (.A(count_cycle[50]), .Y(_11248_));
NOT_g _16855_ (.A(count_cycle[52]), .Y(_11249_));
NOT_g _16856_ (.A(count_cycle[54]), .Y(_11250_));
NOT_g _16857_ (.A(count_cycle[56]), .Y(_11251_));
NOT_g _16858_ (.A(count_cycle[58]), .Y(_11252_));
NOT_g _16859_ (.A(count_cycle[60]), .Y(_11253_));
NOT_g _16860_ (.A(count_cycle[62]), .Y(_11254_));
NOR_g _16861_ (.A(cpu_state[0]), .B(cpu_state[1]), .Y(_11255_));
NOR_g _16862_ (.A(cpu_state[3]), .B(cpu_state[2]), .Y(_11256_));
AND_g _16863_ (.A(_11205_), .B(_11255_), .Y(_11257_));
AND_g _16864_ (.A(_11255_), .B(_11256_), .Y(_11258_));
NOR_g _16865_ (.A(cpu_state[4]), .B(cpu_state[5]), .Y(_11259_));
AND_g _16866_ (.A(_11203_), .B(_11259_), .Y(_11260_));
AND_g _16867_ (.A(cpu_state[6]), .B(_11260_), .Y(_11261_));
AND_g _16868_ (.A(_11258_), .B(_11261_), .Y(_11262_));
NAND_g _16869_ (.A(_11258_), .B(_11261_), .Y(_11263_));
NAND_g _16870_ (.A(decoder_trigger), .B(_11262_), .Y(_11264_));
NOT_g _16871_ (.A(_11264_), .Y(launch_next_insn));
NOR_g _16872_ (.A(latched_branch), .B(latched_store), .Y(_11265_));
NOT_g _16873_ (.A(_11265_), .Y(_11266_));
NOR_g _16874_ (.A(cpu_state[7]), .B(cpu_state[6]), .Y(_11267_));
AND_g _16875_ (.A(_11259_), .B(_11267_), .Y(_11268_));
NAND_g _16876_ (.A(cpu_state[3]), .B(_11255_), .Y(_11269_));
NOR_g _16877_ (.A(cpu_state[2]), .B(_11269_), .Y(_11270_));
AND_g _16878_ (.A(_11268_), .B(_11270_), .Y(_11271_));
NAND_g _16879_ (.A(_11268_), .B(_11270_), .Y(_11272_));
AND_g _16880_ (.A(_10902_), .B(_11271_), .Y(_11273_));
NOT_g _16881_ (.A(_11273_), .Y(_11274_));
AND_g _16882_ (.A(resetn), .B(_11262_), .Y(_11275_));
NAND_g _16883_ (.A(_11266_), .B(_11275_), .Y(_11276_));
NOR_g _16884_ (.A(latched_rd[2]), .B(latched_rd[4]), .Y(_11277_));
NOR_g _16885_ (.A(latched_rd[0]), .B(latched_rd[1]), .Y(_11278_));
NOT_g _16886_ (.A(_11278_), .Y(_11279_));
AND_g _16887_ (.A(_11277_), .B(_11278_), .Y(_11280_));
AND_g _16888_ (.A(_11043_), .B(_11280_), .Y(_11281_));
NOR_g _16889_ (.A(_11276_), .B(_11281_), .Y(_11282_));
NOR_g _16890_ (.A(_11043_), .B(_11276_), .Y(_11283_));
NOR_g _16891_ (.A(_11042_), .B(_11276_), .Y(_11284_));
NAND_g _16892_ (.A(latched_rd[2]), .B(_11282_), .Y(_11285_));
AND_g _16893_ (.A(latched_rd[2]), .B(_11283_), .Y(_11286_));
AND_g _16894_ (.A(latched_rd[4]), .B(_11286_), .Y(_11287_));
NAND_g _16895_ (.A(latched_rd[0]), .B(_11282_), .Y(_11288_));
NOR_g _16896_ (.A(latched_rd[1]), .B(_11288_), .Y(_11289_));
AND_g _16897_ (.A(_11287_), .B(_11289_), .Y(_11290_));
NAND_g _16898_ (.A(_11287_), .B(_11289_), .Y(_11291_));
NAND_g _16899_ (.A(cpuregs_29[0]), .B(_11291_), .Y(_11292_));
NAND_g _16900_ (.A(reg_next_pc[0]), .B(latched_branch), .Y(_11293_));
NAND_g _16901_ (.A(latched_stalu), .B(_11222_), .Y(_11294_));
NOR_g _16902_ (.A(latched_stalu), .B(reg_out[0]), .Y(_11295_));
NOT_g _16903_ (.A(_11295_), .Y(_11296_));
AND_g _16904_ (.A(_10896_), .B(latched_store), .Y(_11297_));
AND_g _16905_ (.A(_11296_), .B(_11297_), .Y(_11298_));
NAND_g _16906_ (.A(_11294_), .B(_11298_), .Y(_11299_));
NAND_g _16907_ (.A(_11293_), .B(_11299_), .Y(_11300_));
AND_g _16908_ (.A(_11282_), .B(_11300_), .Y(_11301_));
NAND_g _16909_ (.A(_11290_), .B(_11301_), .Y(_11302_));
NAND_g _16910_ (.A(_11292_), .B(_11302_), .Y(_00023_));
NAND_g _16911_ (.A(cpuregs_29[1]), .B(_11291_), .Y(_11303_));
NAND_g _16912_ (.A(latched_stalu), .B(alu_out_q[1]), .Y(_11304_));
NAND_g _16913_ (.A(_10897_), .B(reg_out[1]), .Y(_11305_));
NAND_g _16914_ (.A(_11304_), .B(_11305_), .Y(_11306_));
NAND_g _16915_ (.A(_11297_), .B(_11306_), .Y(_11307_));
NAND_g _16916_ (.A(latched_branch), .B(reg_pc[1]), .Y(_11308_));
NAND_g _16917_ (.A(_11307_), .B(_11308_), .Y(_11309_));
AND_g _16918_ (.A(_11282_), .B(_11309_), .Y(_11310_));
NAND_g _16919_ (.A(_11290_), .B(_11310_), .Y(_11311_));
NAND_g _16920_ (.A(_11303_), .B(_11311_), .Y(_00024_));
NAND_g _16921_ (.A(cpuregs_29[2]), .B(_11291_), .Y(_11312_));
NAND_g _16922_ (.A(latched_stalu), .B(alu_out_q[2]), .Y(_11313_));
NAND_g _16923_ (.A(_10897_), .B(reg_out[2]), .Y(_11314_));
NAND_g _16924_ (.A(_11313_), .B(_11314_), .Y(_11315_));
NAND_g _16925_ (.A(_11297_), .B(_11315_), .Y(_11316_));
NAND_g _16926_ (.A(latched_branch), .B(_10900_), .Y(_11317_));
NAND_g _16927_ (.A(_11316_), .B(_11317_), .Y(_11318_));
AND_g _16928_ (.A(_11282_), .B(_11318_), .Y(_11319_));
NAND_g _16929_ (.A(_11290_), .B(_11319_), .Y(_11320_));
NAND_g _16930_ (.A(_11312_), .B(_11320_), .Y(_00025_));
NAND_g _16931_ (.A(cpuregs_29[3]), .B(_11291_), .Y(_11321_));
NAND_g _16932_ (.A(latched_stalu), .B(alu_out_q[3]), .Y(_11322_));
NAND_g _16933_ (.A(_10897_), .B(reg_out[3]), .Y(_11323_));
NAND_g _16934_ (.A(_11322_), .B(_11323_), .Y(_11324_));
NAND_g _16935_ (.A(_11297_), .B(_11324_), .Y(_11325_));
NOR_g _16936_ (.A(reg_pc[3]), .B(reg_pc[2]), .Y(_11326_));
AND_g _16937_ (.A(reg_pc[3]), .B(reg_pc[2]), .Y(_11327_));
NAND_g _16938_ (.A(reg_pc[3]), .B(reg_pc[2]), .Y(_11328_));
NOR_g _16939_ (.A(_10896_), .B(_11326_), .Y(_11329_));
NAND_g _16940_ (.A(_11328_), .B(_11329_), .Y(_11330_));
NAND_g _16941_ (.A(_11325_), .B(_11330_), .Y(_11331_));
AND_g _16942_ (.A(_11282_), .B(_11331_), .Y(_11332_));
NAND_g _16943_ (.A(_11290_), .B(_11332_), .Y(_11333_));
NAND_g _16944_ (.A(_11321_), .B(_11333_), .Y(_00026_));
NAND_g _16945_ (.A(cpuregs_29[4]), .B(_11291_), .Y(_11334_));
NAND_g _16946_ (.A(latched_stalu), .B(alu_out_q[4]), .Y(_11335_));
NAND_g _16947_ (.A(_10897_), .B(reg_out[4]), .Y(_11336_));
NAND_g _16948_ (.A(_11335_), .B(_11336_), .Y(_11337_));
NAND_g _16949_ (.A(_11297_), .B(_11337_), .Y(_11338_));
NOR_g _16950_ (.A(reg_pc[4]), .B(_11327_), .Y(_11339_));
AND_g _16951_ (.A(reg_pc[4]), .B(_11327_), .Y(_11340_));
NAND_g _16952_ (.A(reg_pc[4]), .B(_11327_), .Y(_11341_));
NOR_g _16953_ (.A(_10896_), .B(_11339_), .Y(_11342_));
NAND_g _16954_ (.A(_11341_), .B(_11342_), .Y(_11343_));
NAND_g _16955_ (.A(_11338_), .B(_11343_), .Y(_11344_));
AND_g _16956_ (.A(_11282_), .B(_11344_), .Y(_11345_));
NAND_g _16957_ (.A(_11290_), .B(_11345_), .Y(_11346_));
NAND_g _16958_ (.A(_11334_), .B(_11346_), .Y(_00027_));
NAND_g _16959_ (.A(cpuregs_29[5]), .B(_11291_), .Y(_11347_));
NAND_g _16960_ (.A(latched_stalu), .B(alu_out_q[5]), .Y(_11348_));
NAND_g _16961_ (.A(_10897_), .B(reg_out[5]), .Y(_11349_));
NAND_g _16962_ (.A(_11348_), .B(_11349_), .Y(_11350_));
NAND_g _16963_ (.A(_11297_), .B(_11350_), .Y(_11351_));
NOR_g _16964_ (.A(reg_pc[5]), .B(_11340_), .Y(_11352_));
AND_g _16965_ (.A(reg_pc[5]), .B(_11340_), .Y(_11353_));
NAND_g _16966_ (.A(reg_pc[5]), .B(_11340_), .Y(_11354_));
NOR_g _16967_ (.A(_10896_), .B(_11352_), .Y(_11355_));
NAND_g _16968_ (.A(_11354_), .B(_11355_), .Y(_11356_));
NAND_g _16969_ (.A(_11351_), .B(_11356_), .Y(_11357_));
AND_g _16970_ (.A(_11282_), .B(_11357_), .Y(_11358_));
NAND_g _16971_ (.A(_11290_), .B(_11358_), .Y(_11359_));
NAND_g _16972_ (.A(_11347_), .B(_11359_), .Y(_00028_));
NAND_g _16973_ (.A(cpuregs_29[6]), .B(_11291_), .Y(_11360_));
NAND_g _16974_ (.A(latched_stalu), .B(alu_out_q[6]), .Y(_11361_));
NAND_g _16975_ (.A(_10897_), .B(reg_out[6]), .Y(_11362_));
NAND_g _16976_ (.A(_11361_), .B(_11362_), .Y(_11363_));
NAND_g _16977_ (.A(_11297_), .B(_11363_), .Y(_11364_));
NOR_g _16978_ (.A(reg_pc[6]), .B(_11353_), .Y(_11365_));
AND_g _16979_ (.A(reg_pc[6]), .B(_11353_), .Y(_11366_));
NAND_g _16980_ (.A(reg_pc[6]), .B(_11353_), .Y(_11367_));
NOR_g _16981_ (.A(_10896_), .B(_11365_), .Y(_11368_));
NAND_g _16982_ (.A(_11367_), .B(_11368_), .Y(_11369_));
NAND_g _16983_ (.A(_11364_), .B(_11369_), .Y(_11370_));
AND_g _16984_ (.A(_11282_), .B(_11370_), .Y(_11371_));
NAND_g _16985_ (.A(_11290_), .B(_11371_), .Y(_11372_));
NAND_g _16986_ (.A(_11360_), .B(_11372_), .Y(_00029_));
NAND_g _16987_ (.A(cpuregs_29[7]), .B(_11291_), .Y(_11373_));
NAND_g _16988_ (.A(latched_stalu), .B(alu_out_q[7]), .Y(_11374_));
NAND_g _16989_ (.A(_10897_), .B(reg_out[7]), .Y(_11375_));
NAND_g _16990_ (.A(_11374_), .B(_11375_), .Y(_11376_));
NAND_g _16991_ (.A(_11297_), .B(_11376_), .Y(_11377_));
NOR_g _16992_ (.A(reg_pc[7]), .B(_11366_), .Y(_11378_));
AND_g _16993_ (.A(reg_pc[7]), .B(_11366_), .Y(_11379_));
NAND_g _16994_ (.A(reg_pc[7]), .B(_11366_), .Y(_11380_));
NOR_g _16995_ (.A(_10896_), .B(_11378_), .Y(_11381_));
NAND_g _16996_ (.A(_11380_), .B(_11381_), .Y(_11382_));
NAND_g _16997_ (.A(_11377_), .B(_11382_), .Y(_11383_));
AND_g _16998_ (.A(_11282_), .B(_11383_), .Y(_11384_));
NAND_g _16999_ (.A(_11290_), .B(_11384_), .Y(_11385_));
NAND_g _17000_ (.A(_11373_), .B(_11385_), .Y(_00030_));
NAND_g _17001_ (.A(cpuregs_29[8]), .B(_11291_), .Y(_11386_));
NAND_g _17002_ (.A(latched_stalu), .B(alu_out_q[8]), .Y(_11387_));
NAND_g _17003_ (.A(_10897_), .B(reg_out[8]), .Y(_11388_));
NAND_g _17004_ (.A(_11387_), .B(_11388_), .Y(_11389_));
NAND_g _17005_ (.A(_11297_), .B(_11389_), .Y(_11390_));
NOR_g _17006_ (.A(reg_pc[8]), .B(_11379_), .Y(_11391_));
AND_g _17007_ (.A(reg_pc[8]), .B(_11379_), .Y(_11392_));
NAND_g _17008_ (.A(reg_pc[8]), .B(_11379_), .Y(_11393_));
NOR_g _17009_ (.A(_10896_), .B(_11391_), .Y(_11394_));
NAND_g _17010_ (.A(_11393_), .B(_11394_), .Y(_11395_));
NAND_g _17011_ (.A(_11390_), .B(_11395_), .Y(_11396_));
AND_g _17012_ (.A(_11282_), .B(_11396_), .Y(_11397_));
NAND_g _17013_ (.A(_11290_), .B(_11397_), .Y(_11398_));
NAND_g _17014_ (.A(_11386_), .B(_11398_), .Y(_00031_));
NAND_g _17015_ (.A(cpuregs_29[9]), .B(_11291_), .Y(_11399_));
NAND_g _17016_ (.A(latched_stalu), .B(alu_out_q[9]), .Y(_11400_));
NAND_g _17017_ (.A(_10897_), .B(reg_out[9]), .Y(_11401_));
NAND_g _17018_ (.A(_11400_), .B(_11401_), .Y(_11402_));
NAND_g _17019_ (.A(_11297_), .B(_11402_), .Y(_11403_));
NOR_g _17020_ (.A(reg_pc[9]), .B(_11392_), .Y(_11404_));
AND_g _17021_ (.A(reg_pc[9]), .B(_11392_), .Y(_11405_));
NAND_g _17022_ (.A(reg_pc[9]), .B(_11392_), .Y(_11406_));
NOR_g _17023_ (.A(_10896_), .B(_11404_), .Y(_11407_));
NAND_g _17024_ (.A(_11406_), .B(_11407_), .Y(_11408_));
NAND_g _17025_ (.A(_11403_), .B(_11408_), .Y(_11409_));
AND_g _17026_ (.A(_11282_), .B(_11409_), .Y(_11410_));
NAND_g _17027_ (.A(_11290_), .B(_11410_), .Y(_11411_));
NAND_g _17028_ (.A(_11399_), .B(_11411_), .Y(_00032_));
NAND_g _17029_ (.A(cpuregs_29[10]), .B(_11291_), .Y(_11412_));
NAND_g _17030_ (.A(latched_stalu), .B(alu_out_q[10]), .Y(_11413_));
NAND_g _17031_ (.A(_10897_), .B(reg_out[10]), .Y(_11414_));
NAND_g _17032_ (.A(_11413_), .B(_11414_), .Y(_11415_));
NAND_g _17033_ (.A(_11297_), .B(_11415_), .Y(_11416_));
NOR_g _17034_ (.A(reg_pc[10]), .B(_11405_), .Y(_11417_));
AND_g _17035_ (.A(reg_pc[10]), .B(_11405_), .Y(_11418_));
NAND_g _17036_ (.A(reg_pc[10]), .B(_11405_), .Y(_11419_));
NOR_g _17037_ (.A(_10896_), .B(_11417_), .Y(_11420_));
NAND_g _17038_ (.A(_11419_), .B(_11420_), .Y(_11421_));
NAND_g _17039_ (.A(_11416_), .B(_11421_), .Y(_11422_));
AND_g _17040_ (.A(_11282_), .B(_11422_), .Y(_11423_));
NAND_g _17041_ (.A(_11290_), .B(_11423_), .Y(_11424_));
NAND_g _17042_ (.A(_11412_), .B(_11424_), .Y(_00033_));
NAND_g _17043_ (.A(cpuregs_29[11]), .B(_11291_), .Y(_11425_));
NAND_g _17044_ (.A(latched_stalu), .B(alu_out_q[11]), .Y(_11426_));
NAND_g _17045_ (.A(_10897_), .B(reg_out[11]), .Y(_11427_));
NAND_g _17046_ (.A(_11426_), .B(_11427_), .Y(_11428_));
NAND_g _17047_ (.A(_11297_), .B(_11428_), .Y(_11429_));
NOR_g _17048_ (.A(reg_pc[11]), .B(_11418_), .Y(_11430_));
AND_g _17049_ (.A(reg_pc[11]), .B(_11418_), .Y(_11431_));
NAND_g _17050_ (.A(reg_pc[11]), .B(_11418_), .Y(_11432_));
NOR_g _17051_ (.A(_10896_), .B(_11430_), .Y(_11433_));
NAND_g _17052_ (.A(_11432_), .B(_11433_), .Y(_11434_));
NAND_g _17053_ (.A(_11429_), .B(_11434_), .Y(_11435_));
AND_g _17054_ (.A(_11282_), .B(_11435_), .Y(_11436_));
NAND_g _17055_ (.A(_11290_), .B(_11436_), .Y(_11437_));
NAND_g _17056_ (.A(_11425_), .B(_11437_), .Y(_00034_));
NAND_g _17057_ (.A(cpuregs_29[12]), .B(_11291_), .Y(_11438_));
NAND_g _17058_ (.A(latched_stalu), .B(alu_out_q[12]), .Y(_11439_));
NAND_g _17059_ (.A(_10897_), .B(reg_out[12]), .Y(_11440_));
NAND_g _17060_ (.A(_11439_), .B(_11440_), .Y(_11441_));
NAND_g _17061_ (.A(_11297_), .B(_11441_), .Y(_11442_));
NOR_g _17062_ (.A(reg_pc[12]), .B(_11431_), .Y(_11443_));
AND_g _17063_ (.A(reg_pc[12]), .B(_11431_), .Y(_11444_));
NAND_g _17064_ (.A(reg_pc[12]), .B(_11431_), .Y(_11445_));
NOR_g _17065_ (.A(_10896_), .B(_11443_), .Y(_11446_));
NAND_g _17066_ (.A(_11445_), .B(_11446_), .Y(_11447_));
NAND_g _17067_ (.A(_11442_), .B(_11447_), .Y(_11448_));
AND_g _17068_ (.A(_11282_), .B(_11448_), .Y(_11449_));
NAND_g _17069_ (.A(_11290_), .B(_11449_), .Y(_11450_));
NAND_g _17070_ (.A(_11438_), .B(_11450_), .Y(_00035_));
NAND_g _17071_ (.A(cpuregs_29[13]), .B(_11291_), .Y(_11451_));
NAND_g _17072_ (.A(latched_stalu), .B(alu_out_q[13]), .Y(_11452_));
NAND_g _17073_ (.A(_10897_), .B(reg_out[13]), .Y(_11453_));
NAND_g _17074_ (.A(_11452_), .B(_11453_), .Y(_11454_));
NAND_g _17075_ (.A(_11297_), .B(_11454_), .Y(_11455_));
NOR_g _17076_ (.A(reg_pc[13]), .B(_11444_), .Y(_11456_));
AND_g _17077_ (.A(reg_pc[13]), .B(_11444_), .Y(_11457_));
NAND_g _17078_ (.A(reg_pc[13]), .B(_11444_), .Y(_11458_));
NOR_g _17079_ (.A(_10896_), .B(_11456_), .Y(_11459_));
NAND_g _17080_ (.A(_11458_), .B(_11459_), .Y(_11460_));
NAND_g _17081_ (.A(_11455_), .B(_11460_), .Y(_11461_));
AND_g _17082_ (.A(_11282_), .B(_11461_), .Y(_11462_));
NAND_g _17083_ (.A(_11290_), .B(_11462_), .Y(_11463_));
NAND_g _17084_ (.A(_11451_), .B(_11463_), .Y(_00036_));
NAND_g _17085_ (.A(cpuregs_29[14]), .B(_11291_), .Y(_11464_));
NAND_g _17086_ (.A(latched_stalu), .B(alu_out_q[14]), .Y(_11465_));
NAND_g _17087_ (.A(_10897_), .B(reg_out[14]), .Y(_11466_));
NAND_g _17088_ (.A(_11465_), .B(_11466_), .Y(_11467_));
NAND_g _17089_ (.A(_11297_), .B(_11467_), .Y(_11468_));
NOR_g _17090_ (.A(reg_pc[14]), .B(_11457_), .Y(_11469_));
AND_g _17091_ (.A(reg_pc[14]), .B(_11457_), .Y(_11470_));
NAND_g _17092_ (.A(reg_pc[14]), .B(_11457_), .Y(_11471_));
NOR_g _17093_ (.A(_10896_), .B(_11469_), .Y(_11472_));
NAND_g _17094_ (.A(_11471_), .B(_11472_), .Y(_11473_));
NAND_g _17095_ (.A(_11468_), .B(_11473_), .Y(_11474_));
AND_g _17096_ (.A(_11282_), .B(_11474_), .Y(_11475_));
NAND_g _17097_ (.A(_11290_), .B(_11475_), .Y(_11476_));
NAND_g _17098_ (.A(_11464_), .B(_11476_), .Y(_00037_));
NAND_g _17099_ (.A(cpuregs_29[15]), .B(_11291_), .Y(_11477_));
NAND_g _17100_ (.A(latched_stalu), .B(alu_out_q[15]), .Y(_11478_));
NAND_g _17101_ (.A(_10897_), .B(reg_out[15]), .Y(_11479_));
NAND_g _17102_ (.A(_11478_), .B(_11479_), .Y(_11480_));
NAND_g _17103_ (.A(_11297_), .B(_11480_), .Y(_11481_));
NOR_g _17104_ (.A(reg_pc[15]), .B(_11470_), .Y(_11482_));
AND_g _17105_ (.A(reg_pc[15]), .B(_11470_), .Y(_11483_));
NAND_g _17106_ (.A(reg_pc[15]), .B(_11470_), .Y(_11484_));
NOR_g _17107_ (.A(_10896_), .B(_11482_), .Y(_11485_));
NAND_g _17108_ (.A(_11484_), .B(_11485_), .Y(_11486_));
NAND_g _17109_ (.A(_11481_), .B(_11486_), .Y(_11487_));
AND_g _17110_ (.A(_11282_), .B(_11487_), .Y(_11488_));
NAND_g _17111_ (.A(_11290_), .B(_11488_), .Y(_11489_));
NAND_g _17112_ (.A(_11477_), .B(_11489_), .Y(_00038_));
NAND_g _17113_ (.A(cpuregs_29[16]), .B(_11291_), .Y(_11490_));
NAND_g _17114_ (.A(latched_stalu), .B(alu_out_q[16]), .Y(_11491_));
NAND_g _17115_ (.A(_10897_), .B(reg_out[16]), .Y(_11492_));
NAND_g _17116_ (.A(_11491_), .B(_11492_), .Y(_11493_));
NAND_g _17117_ (.A(_11297_), .B(_11493_), .Y(_11494_));
NOR_g _17118_ (.A(reg_pc[16]), .B(_11483_), .Y(_11495_));
AND_g _17119_ (.A(reg_pc[16]), .B(_11483_), .Y(_11496_));
NAND_g _17120_ (.A(reg_pc[16]), .B(_11483_), .Y(_11497_));
NOR_g _17121_ (.A(_10896_), .B(_11495_), .Y(_11498_));
NAND_g _17122_ (.A(_11497_), .B(_11498_), .Y(_11499_));
NAND_g _17123_ (.A(_11494_), .B(_11499_), .Y(_11500_));
AND_g _17124_ (.A(_11282_), .B(_11500_), .Y(_11501_));
NAND_g _17125_ (.A(_11290_), .B(_11501_), .Y(_11502_));
NAND_g _17126_ (.A(_11490_), .B(_11502_), .Y(_00039_));
NAND_g _17127_ (.A(cpuregs_29[17]), .B(_11291_), .Y(_11503_));
NAND_g _17128_ (.A(latched_stalu), .B(alu_out_q[17]), .Y(_11504_));
NAND_g _17129_ (.A(_10897_), .B(reg_out[17]), .Y(_11505_));
NAND_g _17130_ (.A(_11504_), .B(_11505_), .Y(_11506_));
NAND_g _17131_ (.A(_11297_), .B(_11506_), .Y(_11507_));
NOR_g _17132_ (.A(reg_pc[17]), .B(_11496_), .Y(_11508_));
AND_g _17133_ (.A(reg_pc[17]), .B(_11496_), .Y(_11509_));
NAND_g _17134_ (.A(reg_pc[17]), .B(_11496_), .Y(_11510_));
NOR_g _17135_ (.A(_10896_), .B(_11508_), .Y(_11511_));
NAND_g _17136_ (.A(_11510_), .B(_11511_), .Y(_11512_));
NAND_g _17137_ (.A(_11507_), .B(_11512_), .Y(_11513_));
AND_g _17138_ (.A(_11282_), .B(_11513_), .Y(_11514_));
NAND_g _17139_ (.A(_11290_), .B(_11514_), .Y(_11515_));
NAND_g _17140_ (.A(_11503_), .B(_11515_), .Y(_00040_));
NAND_g _17141_ (.A(cpuregs_29[18]), .B(_11291_), .Y(_11516_));
NAND_g _17142_ (.A(latched_stalu), .B(alu_out_q[18]), .Y(_11517_));
NAND_g _17143_ (.A(_10897_), .B(reg_out[18]), .Y(_11518_));
NAND_g _17144_ (.A(_11517_), .B(_11518_), .Y(_11519_));
NAND_g _17145_ (.A(_11297_), .B(_11519_), .Y(_11520_));
NOR_g _17146_ (.A(reg_pc[18]), .B(_11509_), .Y(_11521_));
AND_g _17147_ (.A(reg_pc[18]), .B(_11509_), .Y(_11522_));
NAND_g _17148_ (.A(reg_pc[18]), .B(_11509_), .Y(_11523_));
NOR_g _17149_ (.A(_10896_), .B(_11521_), .Y(_11524_));
NAND_g _17150_ (.A(_11523_), .B(_11524_), .Y(_11525_));
NAND_g _17151_ (.A(_11520_), .B(_11525_), .Y(_11526_));
AND_g _17152_ (.A(_11282_), .B(_11526_), .Y(_11527_));
NAND_g _17153_ (.A(_11290_), .B(_11527_), .Y(_11528_));
NAND_g _17154_ (.A(_11516_), .B(_11528_), .Y(_00041_));
NAND_g _17155_ (.A(cpuregs_29[19]), .B(_11291_), .Y(_11529_));
NAND_g _17156_ (.A(latched_stalu), .B(alu_out_q[19]), .Y(_11530_));
NAND_g _17157_ (.A(_10897_), .B(reg_out[19]), .Y(_11531_));
NAND_g _17158_ (.A(_11530_), .B(_11531_), .Y(_11532_));
NAND_g _17159_ (.A(_11297_), .B(_11532_), .Y(_11533_));
NOR_g _17160_ (.A(reg_pc[19]), .B(_11522_), .Y(_11534_));
AND_g _17161_ (.A(reg_pc[19]), .B(_11522_), .Y(_11535_));
NAND_g _17162_ (.A(reg_pc[19]), .B(_11522_), .Y(_11536_));
NOR_g _17163_ (.A(_10896_), .B(_11534_), .Y(_11537_));
NAND_g _17164_ (.A(_11536_), .B(_11537_), .Y(_11538_));
NAND_g _17165_ (.A(_11533_), .B(_11538_), .Y(_11539_));
AND_g _17166_ (.A(_11282_), .B(_11539_), .Y(_11540_));
NAND_g _17167_ (.A(_11290_), .B(_11540_), .Y(_11541_));
NAND_g _17168_ (.A(_11529_), .B(_11541_), .Y(_00042_));
NAND_g _17169_ (.A(cpuregs_29[20]), .B(_11291_), .Y(_11542_));
NAND_g _17170_ (.A(latched_stalu), .B(alu_out_q[20]), .Y(_11543_));
NAND_g _17171_ (.A(_10897_), .B(reg_out[20]), .Y(_11544_));
NAND_g _17172_ (.A(_11543_), .B(_11544_), .Y(_11545_));
NAND_g _17173_ (.A(_11297_), .B(_11545_), .Y(_11546_));
NOR_g _17174_ (.A(reg_pc[20]), .B(_11535_), .Y(_11547_));
AND_g _17175_ (.A(reg_pc[20]), .B(_11535_), .Y(_11548_));
NAND_g _17176_ (.A(reg_pc[20]), .B(_11535_), .Y(_11549_));
NOR_g _17177_ (.A(_10896_), .B(_11547_), .Y(_11550_));
NAND_g _17178_ (.A(_11549_), .B(_11550_), .Y(_11551_));
NAND_g _17179_ (.A(_11546_), .B(_11551_), .Y(_11552_));
AND_g _17180_ (.A(_11282_), .B(_11552_), .Y(_11553_));
NAND_g _17181_ (.A(_11290_), .B(_11553_), .Y(_11554_));
NAND_g _17182_ (.A(_11542_), .B(_11554_), .Y(_00043_));
NAND_g _17183_ (.A(cpuregs_29[21]), .B(_11291_), .Y(_11555_));
NAND_g _17184_ (.A(latched_stalu), .B(alu_out_q[21]), .Y(_11556_));
NAND_g _17185_ (.A(_10897_), .B(reg_out[21]), .Y(_11557_));
NAND_g _17186_ (.A(_11556_), .B(_11557_), .Y(_11558_));
NAND_g _17187_ (.A(_11297_), .B(_11558_), .Y(_11559_));
NOR_g _17188_ (.A(reg_pc[21]), .B(_11548_), .Y(_11560_));
AND_g _17189_ (.A(reg_pc[21]), .B(_11548_), .Y(_11561_));
NAND_g _17190_ (.A(reg_pc[21]), .B(_11548_), .Y(_11562_));
NOR_g _17191_ (.A(_10896_), .B(_11560_), .Y(_11563_));
NAND_g _17192_ (.A(_11562_), .B(_11563_), .Y(_11564_));
NAND_g _17193_ (.A(_11559_), .B(_11564_), .Y(_11565_));
AND_g _17194_ (.A(_11282_), .B(_11565_), .Y(_11566_));
NAND_g _17195_ (.A(_11290_), .B(_11566_), .Y(_11567_));
NAND_g _17196_ (.A(_11555_), .B(_11567_), .Y(_00044_));
NAND_g _17197_ (.A(cpuregs_29[22]), .B(_11291_), .Y(_11568_));
NAND_g _17198_ (.A(latched_stalu), .B(alu_out_q[22]), .Y(_11569_));
NAND_g _17199_ (.A(_10897_), .B(reg_out[22]), .Y(_11570_));
NAND_g _17200_ (.A(_11569_), .B(_11570_), .Y(_11571_));
NAND_g _17201_ (.A(_11297_), .B(_11571_), .Y(_11572_));
NOR_g _17202_ (.A(reg_pc[22]), .B(_11561_), .Y(_11573_));
AND_g _17203_ (.A(reg_pc[22]), .B(_11561_), .Y(_11574_));
NAND_g _17204_ (.A(reg_pc[22]), .B(_11561_), .Y(_11575_));
NOR_g _17205_ (.A(_10896_), .B(_11573_), .Y(_11576_));
NAND_g _17206_ (.A(_11575_), .B(_11576_), .Y(_11577_));
NAND_g _17207_ (.A(_11572_), .B(_11577_), .Y(_11578_));
AND_g _17208_ (.A(_11282_), .B(_11578_), .Y(_11579_));
NAND_g _17209_ (.A(_11290_), .B(_11579_), .Y(_11580_));
NAND_g _17210_ (.A(_11568_), .B(_11580_), .Y(_00045_));
NAND_g _17211_ (.A(cpuregs_29[23]), .B(_11291_), .Y(_11581_));
NAND_g _17212_ (.A(latched_stalu), .B(alu_out_q[23]), .Y(_11582_));
NAND_g _17213_ (.A(_10897_), .B(reg_out[23]), .Y(_11583_));
NAND_g _17214_ (.A(_11582_), .B(_11583_), .Y(_11584_));
NAND_g _17215_ (.A(_11297_), .B(_11584_), .Y(_11585_));
NOR_g _17216_ (.A(reg_pc[23]), .B(_11574_), .Y(_11586_));
AND_g _17217_ (.A(reg_pc[23]), .B(_11574_), .Y(_11587_));
NAND_g _17218_ (.A(reg_pc[23]), .B(_11574_), .Y(_11588_));
NOR_g _17219_ (.A(_10896_), .B(_11586_), .Y(_11589_));
NAND_g _17220_ (.A(_11588_), .B(_11589_), .Y(_11590_));
NAND_g _17221_ (.A(_11585_), .B(_11590_), .Y(_11591_));
AND_g _17222_ (.A(_11282_), .B(_11591_), .Y(_11592_));
NAND_g _17223_ (.A(_11290_), .B(_11592_), .Y(_11593_));
NAND_g _17224_ (.A(_11581_), .B(_11593_), .Y(_00046_));
NAND_g _17225_ (.A(cpuregs_29[24]), .B(_11291_), .Y(_11594_));
NAND_g _17226_ (.A(latched_stalu), .B(alu_out_q[24]), .Y(_11595_));
NAND_g _17227_ (.A(_10897_), .B(reg_out[24]), .Y(_11596_));
NAND_g _17228_ (.A(_11595_), .B(_11596_), .Y(_11597_));
NAND_g _17229_ (.A(_11297_), .B(_11597_), .Y(_11598_));
NOR_g _17230_ (.A(reg_pc[24]), .B(_11587_), .Y(_11599_));
AND_g _17231_ (.A(reg_pc[24]), .B(_11587_), .Y(_11600_));
NAND_g _17232_ (.A(reg_pc[24]), .B(_11587_), .Y(_11601_));
NOR_g _17233_ (.A(_10896_), .B(_11599_), .Y(_11602_));
NAND_g _17234_ (.A(_11601_), .B(_11602_), .Y(_11603_));
NAND_g _17235_ (.A(_11598_), .B(_11603_), .Y(_11604_));
AND_g _17236_ (.A(_11282_), .B(_11604_), .Y(_11605_));
NAND_g _17237_ (.A(_11290_), .B(_11605_), .Y(_11606_));
NAND_g _17238_ (.A(_11594_), .B(_11606_), .Y(_00047_));
NAND_g _17239_ (.A(cpuregs_29[25]), .B(_11291_), .Y(_11607_));
NAND_g _17240_ (.A(latched_stalu), .B(alu_out_q[25]), .Y(_11608_));
NAND_g _17241_ (.A(_10897_), .B(reg_out[25]), .Y(_11609_));
NAND_g _17242_ (.A(_11608_), .B(_11609_), .Y(_11610_));
NAND_g _17243_ (.A(_11297_), .B(_11610_), .Y(_11611_));
NOR_g _17244_ (.A(reg_pc[25]), .B(_11600_), .Y(_11612_));
AND_g _17245_ (.A(reg_pc[25]), .B(_11600_), .Y(_11613_));
NAND_g _17246_ (.A(reg_pc[25]), .B(_11600_), .Y(_11614_));
NOR_g _17247_ (.A(_10896_), .B(_11612_), .Y(_11615_));
NAND_g _17248_ (.A(_11614_), .B(_11615_), .Y(_11616_));
NAND_g _17249_ (.A(_11611_), .B(_11616_), .Y(_11617_));
AND_g _17250_ (.A(_11282_), .B(_11617_), .Y(_11618_));
NAND_g _17251_ (.A(_11290_), .B(_11618_), .Y(_11619_));
NAND_g _17252_ (.A(_11607_), .B(_11619_), .Y(_00048_));
NAND_g _17253_ (.A(cpuregs_29[26]), .B(_11291_), .Y(_11620_));
NAND_g _17254_ (.A(latched_stalu), .B(alu_out_q[26]), .Y(_11621_));
NAND_g _17255_ (.A(_10897_), .B(reg_out[26]), .Y(_11622_));
NAND_g _17256_ (.A(_11621_), .B(_11622_), .Y(_11623_));
NAND_g _17257_ (.A(_11297_), .B(_11623_), .Y(_11624_));
NOR_g _17258_ (.A(reg_pc[26]), .B(_11613_), .Y(_11625_));
AND_g _17259_ (.A(reg_pc[26]), .B(_11613_), .Y(_11626_));
NAND_g _17260_ (.A(reg_pc[26]), .B(_11613_), .Y(_11627_));
NOR_g _17261_ (.A(_10896_), .B(_11625_), .Y(_11628_));
NAND_g _17262_ (.A(_11627_), .B(_11628_), .Y(_11629_));
NAND_g _17263_ (.A(_11624_), .B(_11629_), .Y(_11630_));
AND_g _17264_ (.A(_11282_), .B(_11630_), .Y(_11631_));
NAND_g _17265_ (.A(_11290_), .B(_11631_), .Y(_11632_));
NAND_g _17266_ (.A(_11620_), .B(_11632_), .Y(_00049_));
NAND_g _17267_ (.A(cpuregs_29[27]), .B(_11291_), .Y(_11633_));
NAND_g _17268_ (.A(latched_stalu), .B(alu_out_q[27]), .Y(_11634_));
NAND_g _17269_ (.A(_10897_), .B(reg_out[27]), .Y(_11635_));
NAND_g _17270_ (.A(_11634_), .B(_11635_), .Y(_11636_));
NAND_g _17271_ (.A(_11297_), .B(_11636_), .Y(_11637_));
NOR_g _17272_ (.A(reg_pc[27]), .B(_11626_), .Y(_11638_));
AND_g _17273_ (.A(reg_pc[27]), .B(_11626_), .Y(_11639_));
NAND_g _17274_ (.A(reg_pc[27]), .B(_11626_), .Y(_11640_));
NOR_g _17275_ (.A(_10896_), .B(_11638_), .Y(_11641_));
NAND_g _17276_ (.A(_11640_), .B(_11641_), .Y(_11642_));
NAND_g _17277_ (.A(_11637_), .B(_11642_), .Y(_11643_));
AND_g _17278_ (.A(_11282_), .B(_11643_), .Y(_11644_));
NAND_g _17279_ (.A(_11290_), .B(_11644_), .Y(_11645_));
NAND_g _17280_ (.A(_11633_), .B(_11645_), .Y(_00050_));
NAND_g _17281_ (.A(cpuregs_29[28]), .B(_11291_), .Y(_11646_));
NAND_g _17282_ (.A(latched_stalu), .B(alu_out_q[28]), .Y(_11647_));
NAND_g _17283_ (.A(_10897_), .B(reg_out[28]), .Y(_11648_));
NAND_g _17284_ (.A(_11647_), .B(_11648_), .Y(_11649_));
NAND_g _17285_ (.A(_11297_), .B(_11649_), .Y(_11650_));
NOR_g _17286_ (.A(reg_pc[28]), .B(_11639_), .Y(_11651_));
AND_g _17287_ (.A(reg_pc[28]), .B(_11639_), .Y(_11652_));
NAND_g _17288_ (.A(reg_pc[28]), .B(_11639_), .Y(_11653_));
NOR_g _17289_ (.A(_10896_), .B(_11651_), .Y(_11654_));
NAND_g _17290_ (.A(_11653_), .B(_11654_), .Y(_11655_));
NAND_g _17291_ (.A(_11650_), .B(_11655_), .Y(_11656_));
AND_g _17292_ (.A(_11282_), .B(_11656_), .Y(_11657_));
NAND_g _17293_ (.A(_11290_), .B(_11657_), .Y(_11658_));
NAND_g _17294_ (.A(_11646_), .B(_11658_), .Y(_00051_));
NAND_g _17295_ (.A(cpuregs_29[29]), .B(_11291_), .Y(_11659_));
NAND_g _17296_ (.A(latched_stalu), .B(alu_out_q[29]), .Y(_11660_));
NAND_g _17297_ (.A(_10897_), .B(reg_out[29]), .Y(_11661_));
NAND_g _17298_ (.A(_11660_), .B(_11661_), .Y(_11662_));
NAND_g _17299_ (.A(_11297_), .B(_11662_), .Y(_11663_));
NOR_g _17300_ (.A(reg_pc[29]), .B(_11652_), .Y(_11664_));
AND_g _17301_ (.A(reg_pc[29]), .B(_11652_), .Y(_11665_));
NAND_g _17302_ (.A(reg_pc[29]), .B(_11652_), .Y(_11666_));
NOR_g _17303_ (.A(_10896_), .B(_11664_), .Y(_11667_));
NAND_g _17304_ (.A(_11666_), .B(_11667_), .Y(_11668_));
NAND_g _17305_ (.A(_11663_), .B(_11668_), .Y(_11669_));
AND_g _17306_ (.A(_11282_), .B(_11669_), .Y(_11670_));
NAND_g _17307_ (.A(_11290_), .B(_11670_), .Y(_11671_));
NAND_g _17308_ (.A(_11659_), .B(_11671_), .Y(_00052_));
NAND_g _17309_ (.A(cpuregs_29[30]), .B(_11291_), .Y(_11672_));
NAND_g _17310_ (.A(latched_stalu), .B(alu_out_q[30]), .Y(_11673_));
NAND_g _17311_ (.A(_10897_), .B(reg_out[30]), .Y(_11674_));
NAND_g _17312_ (.A(_11673_), .B(_11674_), .Y(_11675_));
NAND_g _17313_ (.A(_11297_), .B(_11675_), .Y(_11676_));
NOR_g _17314_ (.A(reg_pc[30]), .B(_11665_), .Y(_11677_));
NAND_g _17315_ (.A(reg_pc[30]), .B(_11665_), .Y(_11678_));
NOT_g _17316_ (.A(_11678_), .Y(_11679_));
NOR_g _17317_ (.A(_10896_), .B(_11677_), .Y(_11680_));
NAND_g _17318_ (.A(_11678_), .B(_11680_), .Y(_11681_));
NAND_g _17319_ (.A(_11676_), .B(_11681_), .Y(_11682_));
AND_g _17320_ (.A(_11282_), .B(_11682_), .Y(_11683_));
NAND_g _17321_ (.A(_11290_), .B(_11683_), .Y(_11684_));
NAND_g _17322_ (.A(_11672_), .B(_11684_), .Y(_00053_));
NAND_g _17323_ (.A(cpuregs_29[31]), .B(_11291_), .Y(_11685_));
NAND_g _17324_ (.A(latched_stalu), .B(alu_out_q[31]), .Y(_11686_));
NAND_g _17325_ (.A(_10897_), .B(reg_out[31]), .Y(_11687_));
NAND_g _17326_ (.A(_11686_), .B(_11687_), .Y(_11688_));
NAND_g _17327_ (.A(_11297_), .B(_11688_), .Y(_11689_));
NAND_g _17328_ (.A(reg_pc[31]), .B(_11679_), .Y(_11690_));
NAND_g _17329_ (.A(_10899_), .B(_11678_), .Y(_11691_));
AND_g _17330_ (.A(latched_branch), .B(_11691_), .Y(_11692_));
NAND_g _17331_ (.A(_11690_), .B(_11692_), .Y(_11693_));
NAND_g _17332_ (.A(_11689_), .B(_11693_), .Y(_11694_));
AND_g _17333_ (.A(_11282_), .B(_11694_), .Y(_11695_));
NAND_g _17334_ (.A(_11290_), .B(_11695_), .Y(_11696_));
NAND_g _17335_ (.A(_11685_), .B(_11696_), .Y(_00054_));
AND_g _17336_ (.A(_11277_), .B(_11283_), .Y(_11697_));
AND_g _17337_ (.A(_11289_), .B(_11697_), .Y(_11698_));
NAND_g _17338_ (.A(_11289_), .B(_11697_), .Y(_11699_));
NAND_g _17339_ (.A(cpuregs_9[0]), .B(_11699_), .Y(_11700_));
NAND_g _17340_ (.A(_11301_), .B(_11698_), .Y(_11701_));
NAND_g _17341_ (.A(_11700_), .B(_11701_), .Y(_00055_));
NAND_g _17342_ (.A(cpuregs_9[1]), .B(_11699_), .Y(_11702_));
NAND_g _17343_ (.A(_11310_), .B(_11698_), .Y(_11703_));
NAND_g _17344_ (.A(_11702_), .B(_11703_), .Y(_00056_));
NAND_g _17345_ (.A(cpuregs_9[2]), .B(_11699_), .Y(_11704_));
NAND_g _17346_ (.A(_11319_), .B(_11698_), .Y(_11705_));
NAND_g _17347_ (.A(_11704_), .B(_11705_), .Y(_00057_));
NAND_g _17348_ (.A(cpuregs_9[3]), .B(_11699_), .Y(_11706_));
NAND_g _17349_ (.A(_11332_), .B(_11698_), .Y(_11707_));
NAND_g _17350_ (.A(_11706_), .B(_11707_), .Y(_00058_));
NAND_g _17351_ (.A(cpuregs_9[4]), .B(_11699_), .Y(_11708_));
NAND_g _17352_ (.A(_11345_), .B(_11698_), .Y(_11709_));
NAND_g _17353_ (.A(_11708_), .B(_11709_), .Y(_00059_));
NAND_g _17354_ (.A(cpuregs_9[5]), .B(_11699_), .Y(_11710_));
NAND_g _17355_ (.A(_11358_), .B(_11698_), .Y(_11711_));
NAND_g _17356_ (.A(_11710_), .B(_11711_), .Y(_00060_));
NAND_g _17357_ (.A(cpuregs_9[6]), .B(_11699_), .Y(_11712_));
NAND_g _17358_ (.A(_11371_), .B(_11698_), .Y(_11713_));
NAND_g _17359_ (.A(_11712_), .B(_11713_), .Y(_00061_));
NAND_g _17360_ (.A(cpuregs_9[7]), .B(_11699_), .Y(_11714_));
NAND_g _17361_ (.A(_11384_), .B(_11698_), .Y(_11715_));
NAND_g _17362_ (.A(_11714_), .B(_11715_), .Y(_00062_));
NAND_g _17363_ (.A(cpuregs_9[8]), .B(_11699_), .Y(_11716_));
NAND_g _17364_ (.A(_11397_), .B(_11698_), .Y(_11717_));
NAND_g _17365_ (.A(_11716_), .B(_11717_), .Y(_00063_));
NAND_g _17366_ (.A(cpuregs_9[9]), .B(_11699_), .Y(_11718_));
NAND_g _17367_ (.A(_11410_), .B(_11698_), .Y(_11719_));
NAND_g _17368_ (.A(_11718_), .B(_11719_), .Y(_00064_));
NAND_g _17369_ (.A(cpuregs_9[10]), .B(_11699_), .Y(_11720_));
NAND_g _17370_ (.A(_11423_), .B(_11698_), .Y(_11721_));
NAND_g _17371_ (.A(_11720_), .B(_11721_), .Y(_00065_));
NAND_g _17372_ (.A(cpuregs_9[11]), .B(_11699_), .Y(_11722_));
NAND_g _17373_ (.A(_11436_), .B(_11698_), .Y(_11723_));
NAND_g _17374_ (.A(_11722_), .B(_11723_), .Y(_00066_));
NAND_g _17375_ (.A(cpuregs_9[12]), .B(_11699_), .Y(_11724_));
NAND_g _17376_ (.A(_11449_), .B(_11698_), .Y(_11725_));
NAND_g _17377_ (.A(_11724_), .B(_11725_), .Y(_00067_));
NAND_g _17378_ (.A(cpuregs_9[13]), .B(_11699_), .Y(_11726_));
NAND_g _17379_ (.A(_11462_), .B(_11698_), .Y(_11727_));
NAND_g _17380_ (.A(_11726_), .B(_11727_), .Y(_00068_));
NAND_g _17381_ (.A(cpuregs_9[14]), .B(_11699_), .Y(_11728_));
NAND_g _17382_ (.A(_11475_), .B(_11698_), .Y(_11729_));
NAND_g _17383_ (.A(_11728_), .B(_11729_), .Y(_00069_));
NAND_g _17384_ (.A(cpuregs_9[15]), .B(_11699_), .Y(_11730_));
NAND_g _17385_ (.A(_11488_), .B(_11698_), .Y(_11731_));
NAND_g _17386_ (.A(_11730_), .B(_11731_), .Y(_00070_));
NAND_g _17387_ (.A(cpuregs_9[16]), .B(_11699_), .Y(_11732_));
NAND_g _17388_ (.A(_11501_), .B(_11698_), .Y(_11733_));
NAND_g _17389_ (.A(_11732_), .B(_11733_), .Y(_00071_));
NAND_g _17390_ (.A(cpuregs_9[17]), .B(_11699_), .Y(_11734_));
NAND_g _17391_ (.A(_11514_), .B(_11698_), .Y(_11735_));
NAND_g _17392_ (.A(_11734_), .B(_11735_), .Y(_00072_));
NAND_g _17393_ (.A(cpuregs_9[18]), .B(_11699_), .Y(_11736_));
NAND_g _17394_ (.A(_11527_), .B(_11698_), .Y(_11737_));
NAND_g _17395_ (.A(_11736_), .B(_11737_), .Y(_00073_));
NAND_g _17396_ (.A(cpuregs_9[19]), .B(_11699_), .Y(_11738_));
NAND_g _17397_ (.A(_11540_), .B(_11698_), .Y(_11739_));
NAND_g _17398_ (.A(_11738_), .B(_11739_), .Y(_00074_));
NAND_g _17399_ (.A(cpuregs_9[20]), .B(_11699_), .Y(_11740_));
NAND_g _17400_ (.A(_11553_), .B(_11698_), .Y(_11741_));
NAND_g _17401_ (.A(_11740_), .B(_11741_), .Y(_00075_));
NAND_g _17402_ (.A(cpuregs_9[21]), .B(_11699_), .Y(_11742_));
NAND_g _17403_ (.A(_11566_), .B(_11698_), .Y(_11743_));
NAND_g _17404_ (.A(_11742_), .B(_11743_), .Y(_00076_));
NAND_g _17405_ (.A(cpuregs_9[22]), .B(_11699_), .Y(_11744_));
NAND_g _17406_ (.A(_11579_), .B(_11698_), .Y(_11745_));
NAND_g _17407_ (.A(_11744_), .B(_11745_), .Y(_00077_));
NAND_g _17408_ (.A(cpuregs_9[23]), .B(_11699_), .Y(_11746_));
NAND_g _17409_ (.A(_11592_), .B(_11698_), .Y(_11747_));
NAND_g _17410_ (.A(_11746_), .B(_11747_), .Y(_00078_));
NAND_g _17411_ (.A(cpuregs_9[24]), .B(_11699_), .Y(_11748_));
NAND_g _17412_ (.A(_11605_), .B(_11698_), .Y(_11749_));
NAND_g _17413_ (.A(_11748_), .B(_11749_), .Y(_00079_));
NAND_g _17414_ (.A(cpuregs_9[25]), .B(_11699_), .Y(_11750_));
NAND_g _17415_ (.A(_11618_), .B(_11698_), .Y(_11751_));
NAND_g _17416_ (.A(_11750_), .B(_11751_), .Y(_00080_));
NAND_g _17417_ (.A(cpuregs_9[26]), .B(_11699_), .Y(_11752_));
NAND_g _17418_ (.A(_11631_), .B(_11698_), .Y(_11753_));
NAND_g _17419_ (.A(_11752_), .B(_11753_), .Y(_00081_));
NAND_g _17420_ (.A(cpuregs_9[27]), .B(_11699_), .Y(_11754_));
NAND_g _17421_ (.A(_11644_), .B(_11698_), .Y(_11755_));
NAND_g _17422_ (.A(_11754_), .B(_11755_), .Y(_00082_));
NAND_g _17423_ (.A(cpuregs_9[28]), .B(_11699_), .Y(_11756_));
NAND_g _17424_ (.A(_11657_), .B(_11698_), .Y(_11757_));
NAND_g _17425_ (.A(_11756_), .B(_11757_), .Y(_00083_));
NAND_g _17426_ (.A(cpuregs_9[29]), .B(_11699_), .Y(_11758_));
NAND_g _17427_ (.A(_11670_), .B(_11698_), .Y(_11759_));
NAND_g _17428_ (.A(_11758_), .B(_11759_), .Y(_00084_));
NAND_g _17429_ (.A(cpuregs_9[30]), .B(_11699_), .Y(_11760_));
NAND_g _17430_ (.A(_11683_), .B(_11698_), .Y(_11761_));
NAND_g _17431_ (.A(_11760_), .B(_11761_), .Y(_00085_));
NAND_g _17432_ (.A(cpuregs_9[31]), .B(_11699_), .Y(_11762_));
NAND_g _17433_ (.A(_11695_), .B(_11698_), .Y(_11763_));
NAND_g _17434_ (.A(_11762_), .B(_11763_), .Y(_00086_));
NAND_g _17435_ (.A(latched_rd[1]), .B(_11282_), .Y(_11764_));
NOR_g _17436_ (.A(latched_rd[0]), .B(_11764_), .Y(_11765_));
NOR_g _17437_ (.A(_11044_), .B(_11276_), .Y(_11766_));
NOR_g _17438_ (.A(_11283_), .B(_11766_), .Y(_11767_));
AND_g _17439_ (.A(_11284_), .B(_11767_), .Y(_11768_));
AND_g _17440_ (.A(_11765_), .B(_11768_), .Y(_11769_));
NAND_g _17441_ (.A(_11765_), .B(_11768_), .Y(_11770_));
NAND_g _17442_ (.A(_11301_), .B(_11769_), .Y(_11771_));
NAND_g _17443_ (.A(cpuregs_6[0]), .B(_11770_), .Y(_11772_));
NAND_g _17444_ (.A(_11771_), .B(_11772_), .Y(_00087_));
NAND_g _17445_ (.A(_11310_), .B(_11769_), .Y(_11773_));
NAND_g _17446_ (.A(cpuregs_6[1]), .B(_11770_), .Y(_11774_));
NAND_g _17447_ (.A(_11773_), .B(_11774_), .Y(_00088_));
NAND_g _17448_ (.A(_11319_), .B(_11769_), .Y(_11775_));
NAND_g _17449_ (.A(cpuregs_6[2]), .B(_11770_), .Y(_11776_));
NAND_g _17450_ (.A(_11775_), .B(_11776_), .Y(_00089_));
NAND_g _17451_ (.A(_11332_), .B(_11769_), .Y(_11777_));
NAND_g _17452_ (.A(cpuregs_6[3]), .B(_11770_), .Y(_11778_));
NAND_g _17453_ (.A(_11777_), .B(_11778_), .Y(_00090_));
NAND_g _17454_ (.A(_11345_), .B(_11769_), .Y(_11779_));
NAND_g _17455_ (.A(cpuregs_6[4]), .B(_11770_), .Y(_11780_));
NAND_g _17456_ (.A(_11779_), .B(_11780_), .Y(_00091_));
NAND_g _17457_ (.A(_11358_), .B(_11769_), .Y(_11781_));
NAND_g _17458_ (.A(cpuregs_6[5]), .B(_11770_), .Y(_11782_));
NAND_g _17459_ (.A(_11781_), .B(_11782_), .Y(_00092_));
NAND_g _17460_ (.A(_11371_), .B(_11769_), .Y(_11783_));
NAND_g _17461_ (.A(cpuregs_6[6]), .B(_11770_), .Y(_11784_));
NAND_g _17462_ (.A(_11783_), .B(_11784_), .Y(_00093_));
NAND_g _17463_ (.A(_11384_), .B(_11769_), .Y(_11785_));
NAND_g _17464_ (.A(cpuregs_6[7]), .B(_11770_), .Y(_11786_));
NAND_g _17465_ (.A(_11785_), .B(_11786_), .Y(_00094_));
NAND_g _17466_ (.A(_11397_), .B(_11769_), .Y(_11787_));
NAND_g _17467_ (.A(cpuregs_6[8]), .B(_11770_), .Y(_11788_));
NAND_g _17468_ (.A(_11787_), .B(_11788_), .Y(_00095_));
NAND_g _17469_ (.A(_11410_), .B(_11769_), .Y(_11789_));
NAND_g _17470_ (.A(cpuregs_6[9]), .B(_11770_), .Y(_11790_));
NAND_g _17471_ (.A(_11789_), .B(_11790_), .Y(_00096_));
NAND_g _17472_ (.A(_11423_), .B(_11769_), .Y(_11791_));
NAND_g _17473_ (.A(cpuregs_6[10]), .B(_11770_), .Y(_11792_));
NAND_g _17474_ (.A(_11791_), .B(_11792_), .Y(_00097_));
NAND_g _17475_ (.A(_11436_), .B(_11769_), .Y(_11793_));
NAND_g _17476_ (.A(cpuregs_6[11]), .B(_11770_), .Y(_11794_));
NAND_g _17477_ (.A(_11793_), .B(_11794_), .Y(_00098_));
NAND_g _17478_ (.A(_11449_), .B(_11769_), .Y(_11795_));
NAND_g _17479_ (.A(cpuregs_6[12]), .B(_11770_), .Y(_11796_));
NAND_g _17480_ (.A(_11795_), .B(_11796_), .Y(_00099_));
NAND_g _17481_ (.A(_11462_), .B(_11769_), .Y(_11797_));
NAND_g _17482_ (.A(cpuregs_6[13]), .B(_11770_), .Y(_11798_));
NAND_g _17483_ (.A(_11797_), .B(_11798_), .Y(_00100_));
NAND_g _17484_ (.A(_11475_), .B(_11769_), .Y(_11799_));
NAND_g _17485_ (.A(cpuregs_6[14]), .B(_11770_), .Y(_11800_));
NAND_g _17486_ (.A(_11799_), .B(_11800_), .Y(_00101_));
NAND_g _17487_ (.A(_11488_), .B(_11769_), .Y(_11801_));
NAND_g _17488_ (.A(cpuregs_6[15]), .B(_11770_), .Y(_11802_));
NAND_g _17489_ (.A(_11801_), .B(_11802_), .Y(_00102_));
NAND_g _17490_ (.A(_11501_), .B(_11769_), .Y(_11803_));
NAND_g _17491_ (.A(cpuregs_6[16]), .B(_11770_), .Y(_11804_));
NAND_g _17492_ (.A(_11803_), .B(_11804_), .Y(_00103_));
NOR_g _17493_ (.A(cpuregs_6[17]), .B(_11769_), .Y(_11805_));
NOR_g _17494_ (.A(_11514_), .B(_11770_), .Y(_11806_));
NOR_g _17495_ (.A(_11805_), .B(_11806_), .Y(_00104_));
NAND_g _17496_ (.A(_11527_), .B(_11769_), .Y(_11807_));
NAND_g _17497_ (.A(cpuregs_6[18]), .B(_11770_), .Y(_11808_));
NAND_g _17498_ (.A(_11807_), .B(_11808_), .Y(_00105_));
NAND_g _17499_ (.A(_11540_), .B(_11769_), .Y(_11809_));
NAND_g _17500_ (.A(cpuregs_6[19]), .B(_11770_), .Y(_11810_));
NAND_g _17501_ (.A(_11809_), .B(_11810_), .Y(_00106_));
NAND_g _17502_ (.A(_11553_), .B(_11769_), .Y(_11811_));
NAND_g _17503_ (.A(cpuregs_6[20]), .B(_11770_), .Y(_11812_));
NAND_g _17504_ (.A(_11811_), .B(_11812_), .Y(_00107_));
NAND_g _17505_ (.A(_11566_), .B(_11769_), .Y(_11813_));
NAND_g _17506_ (.A(cpuregs_6[21]), .B(_11770_), .Y(_11814_));
NAND_g _17507_ (.A(_11813_), .B(_11814_), .Y(_00108_));
NAND_g _17508_ (.A(_11579_), .B(_11769_), .Y(_11815_));
NAND_g _17509_ (.A(cpuregs_6[22]), .B(_11770_), .Y(_11816_));
NAND_g _17510_ (.A(_11815_), .B(_11816_), .Y(_00109_));
NAND_g _17511_ (.A(_11592_), .B(_11769_), .Y(_11817_));
NAND_g _17512_ (.A(cpuregs_6[23]), .B(_11770_), .Y(_11818_));
NAND_g _17513_ (.A(_11817_), .B(_11818_), .Y(_00110_));
NAND_g _17514_ (.A(_11605_), .B(_11769_), .Y(_11819_));
NAND_g _17515_ (.A(cpuregs_6[24]), .B(_11770_), .Y(_11820_));
NAND_g _17516_ (.A(_11819_), .B(_11820_), .Y(_00111_));
NAND_g _17517_ (.A(_11618_), .B(_11769_), .Y(_11821_));
NAND_g _17518_ (.A(cpuregs_6[25]), .B(_11770_), .Y(_11822_));
NAND_g _17519_ (.A(_11821_), .B(_11822_), .Y(_00112_));
NAND_g _17520_ (.A(_11631_), .B(_11769_), .Y(_11823_));
NAND_g _17521_ (.A(cpuregs_6[26]), .B(_11770_), .Y(_11824_));
NAND_g _17522_ (.A(_11823_), .B(_11824_), .Y(_00113_));
NAND_g _17523_ (.A(_11644_), .B(_11769_), .Y(_11825_));
NAND_g _17524_ (.A(cpuregs_6[27]), .B(_11770_), .Y(_11826_));
NAND_g _17525_ (.A(_11825_), .B(_11826_), .Y(_00114_));
NAND_g _17526_ (.A(_11657_), .B(_11769_), .Y(_11827_));
NAND_g _17527_ (.A(cpuregs_6[28]), .B(_11770_), .Y(_11828_));
NAND_g _17528_ (.A(_11827_), .B(_11828_), .Y(_00115_));
NAND_g _17529_ (.A(_11670_), .B(_11769_), .Y(_11829_));
NAND_g _17530_ (.A(cpuregs_6[29]), .B(_11770_), .Y(_11830_));
NAND_g _17531_ (.A(_11829_), .B(_11830_), .Y(_00116_));
NAND_g _17532_ (.A(_11683_), .B(_11769_), .Y(_11831_));
NAND_g _17533_ (.A(cpuregs_6[30]), .B(_11770_), .Y(_11832_));
NAND_g _17534_ (.A(_11831_), .B(_11832_), .Y(_00117_));
NAND_g _17535_ (.A(_11695_), .B(_11769_), .Y(_11833_));
NAND_g _17536_ (.A(cpuregs_6[31]), .B(_11770_), .Y(_11834_));
NAND_g _17537_ (.A(_11833_), .B(_11834_), .Y(_00118_));
NAND_g _17538_ (.A(_11043_), .B(_11766_), .Y(_11835_));
NOR_g _17539_ (.A(latched_rd[2]), .B(_11835_), .Y(_11836_));
AND_g _17540_ (.A(_11765_), .B(_11836_), .Y(_11837_));
NAND_g _17541_ (.A(_11765_), .B(_11836_), .Y(_11838_));
NAND_g _17542_ (.A(_11301_), .B(_11837_), .Y(_11839_));
NAND_g _17543_ (.A(cpuregs_18[0]), .B(_11838_), .Y(_11840_));
NAND_g _17544_ (.A(_11839_), .B(_11840_), .Y(_00119_));
NAND_g _17545_ (.A(_11310_), .B(_11837_), .Y(_11841_));
NAND_g _17546_ (.A(cpuregs_18[1]), .B(_11838_), .Y(_11842_));
NAND_g _17547_ (.A(_11841_), .B(_11842_), .Y(_00120_));
NAND_g _17548_ (.A(_11319_), .B(_11837_), .Y(_11843_));
NAND_g _17549_ (.A(cpuregs_18[2]), .B(_11838_), .Y(_11844_));
NAND_g _17550_ (.A(_11843_), .B(_11844_), .Y(_00121_));
NAND_g _17551_ (.A(_11332_), .B(_11837_), .Y(_11845_));
NAND_g _17552_ (.A(cpuregs_18[3]), .B(_11838_), .Y(_11846_));
NAND_g _17553_ (.A(_11845_), .B(_11846_), .Y(_00122_));
NAND_g _17554_ (.A(_11345_), .B(_11837_), .Y(_11847_));
NAND_g _17555_ (.A(cpuregs_18[4]), .B(_11838_), .Y(_11848_));
NAND_g _17556_ (.A(_11847_), .B(_11848_), .Y(_00123_));
NAND_g _17557_ (.A(_11358_), .B(_11837_), .Y(_11849_));
NAND_g _17558_ (.A(cpuregs_18[5]), .B(_11838_), .Y(_11850_));
NAND_g _17559_ (.A(_11849_), .B(_11850_), .Y(_00124_));
NAND_g _17560_ (.A(_11371_), .B(_11837_), .Y(_11851_));
NAND_g _17561_ (.A(cpuregs_18[6]), .B(_11838_), .Y(_11852_));
NAND_g _17562_ (.A(_11851_), .B(_11852_), .Y(_00125_));
NAND_g _17563_ (.A(_11384_), .B(_11837_), .Y(_11853_));
NAND_g _17564_ (.A(cpuregs_18[7]), .B(_11838_), .Y(_11854_));
NAND_g _17565_ (.A(_11853_), .B(_11854_), .Y(_00126_));
NAND_g _17566_ (.A(_11397_), .B(_11837_), .Y(_11855_));
NAND_g _17567_ (.A(cpuregs_18[8]), .B(_11838_), .Y(_11856_));
NAND_g _17568_ (.A(_11855_), .B(_11856_), .Y(_00127_));
NAND_g _17569_ (.A(_11410_), .B(_11837_), .Y(_11857_));
NAND_g _17570_ (.A(cpuregs_18[9]), .B(_11838_), .Y(_11858_));
NAND_g _17571_ (.A(_11857_), .B(_11858_), .Y(_00128_));
NAND_g _17572_ (.A(_11423_), .B(_11837_), .Y(_11859_));
NAND_g _17573_ (.A(cpuregs_18[10]), .B(_11838_), .Y(_11860_));
NAND_g _17574_ (.A(_11859_), .B(_11860_), .Y(_00129_));
NAND_g _17575_ (.A(_11436_), .B(_11837_), .Y(_11861_));
NAND_g _17576_ (.A(cpuregs_18[11]), .B(_11838_), .Y(_11862_));
NAND_g _17577_ (.A(_11861_), .B(_11862_), .Y(_00130_));
NAND_g _17578_ (.A(_11449_), .B(_11837_), .Y(_11863_));
NAND_g _17579_ (.A(cpuregs_18[12]), .B(_11838_), .Y(_11864_));
NAND_g _17580_ (.A(_11863_), .B(_11864_), .Y(_00131_));
NAND_g _17581_ (.A(_11462_), .B(_11837_), .Y(_11865_));
NAND_g _17582_ (.A(cpuregs_18[13]), .B(_11838_), .Y(_11866_));
NAND_g _17583_ (.A(_11865_), .B(_11866_), .Y(_00132_));
NAND_g _17584_ (.A(_11475_), .B(_11837_), .Y(_11867_));
NAND_g _17585_ (.A(cpuregs_18[14]), .B(_11838_), .Y(_11868_));
NAND_g _17586_ (.A(_11867_), .B(_11868_), .Y(_00133_));
NAND_g _17587_ (.A(_11488_), .B(_11837_), .Y(_11869_));
NAND_g _17588_ (.A(cpuregs_18[15]), .B(_11838_), .Y(_11870_));
NAND_g _17589_ (.A(_11869_), .B(_11870_), .Y(_00134_));
NAND_g _17590_ (.A(_11501_), .B(_11837_), .Y(_11871_));
NAND_g _17591_ (.A(cpuregs_18[16]), .B(_11838_), .Y(_11872_));
NAND_g _17592_ (.A(_11871_), .B(_11872_), .Y(_00135_));
NOR_g _17593_ (.A(cpuregs_18[17]), .B(_11837_), .Y(_11873_));
NOR_g _17594_ (.A(_11514_), .B(_11838_), .Y(_11874_));
NOR_g _17595_ (.A(_11873_), .B(_11874_), .Y(_00136_));
NAND_g _17596_ (.A(_11527_), .B(_11837_), .Y(_11875_));
NAND_g _17597_ (.A(cpuregs_18[18]), .B(_11838_), .Y(_11876_));
NAND_g _17598_ (.A(_11875_), .B(_11876_), .Y(_00137_));
NAND_g _17599_ (.A(_11540_), .B(_11837_), .Y(_11877_));
NAND_g _17600_ (.A(cpuregs_18[19]), .B(_11838_), .Y(_11878_));
NAND_g _17601_ (.A(_11877_), .B(_11878_), .Y(_00138_));
NAND_g _17602_ (.A(_11553_), .B(_11837_), .Y(_11879_));
NAND_g _17603_ (.A(cpuregs_18[20]), .B(_11838_), .Y(_11880_));
NAND_g _17604_ (.A(_11879_), .B(_11880_), .Y(_00139_));
NAND_g _17605_ (.A(_11566_), .B(_11837_), .Y(_11881_));
NAND_g _17606_ (.A(cpuregs_18[21]), .B(_11838_), .Y(_11882_));
NAND_g _17607_ (.A(_11881_), .B(_11882_), .Y(_00140_));
NAND_g _17608_ (.A(_11579_), .B(_11837_), .Y(_11883_));
NAND_g _17609_ (.A(cpuregs_18[22]), .B(_11838_), .Y(_11884_));
NAND_g _17610_ (.A(_11883_), .B(_11884_), .Y(_00141_));
NAND_g _17611_ (.A(_11592_), .B(_11837_), .Y(_11885_));
NAND_g _17612_ (.A(cpuregs_18[23]), .B(_11838_), .Y(_11886_));
NAND_g _17613_ (.A(_11885_), .B(_11886_), .Y(_00142_));
NAND_g _17614_ (.A(_11605_), .B(_11837_), .Y(_11887_));
NAND_g _17615_ (.A(cpuregs_18[24]), .B(_11838_), .Y(_11888_));
NAND_g _17616_ (.A(_11887_), .B(_11888_), .Y(_00143_));
NAND_g _17617_ (.A(_11618_), .B(_11837_), .Y(_11889_));
NAND_g _17618_ (.A(cpuregs_18[25]), .B(_11838_), .Y(_11890_));
NAND_g _17619_ (.A(_11889_), .B(_11890_), .Y(_00144_));
NAND_g _17620_ (.A(_11631_), .B(_11837_), .Y(_11891_));
NAND_g _17621_ (.A(cpuregs_18[26]), .B(_11838_), .Y(_11892_));
NAND_g _17622_ (.A(_11891_), .B(_11892_), .Y(_00145_));
NAND_g _17623_ (.A(_11644_), .B(_11837_), .Y(_11893_));
NAND_g _17624_ (.A(cpuregs_18[27]), .B(_11838_), .Y(_11894_));
NAND_g _17625_ (.A(_11893_), .B(_11894_), .Y(_00146_));
NAND_g _17626_ (.A(_11657_), .B(_11837_), .Y(_11895_));
NAND_g _17627_ (.A(cpuregs_18[28]), .B(_11838_), .Y(_11896_));
NAND_g _17628_ (.A(_11895_), .B(_11896_), .Y(_00147_));
NAND_g _17629_ (.A(_11670_), .B(_11837_), .Y(_11897_));
NAND_g _17630_ (.A(cpuregs_18[29]), .B(_11838_), .Y(_11898_));
NAND_g _17631_ (.A(_11897_), .B(_11898_), .Y(_00148_));
NAND_g _17632_ (.A(_11683_), .B(_11837_), .Y(_11899_));
NAND_g _17633_ (.A(cpuregs_18[30]), .B(_11838_), .Y(_11900_));
NAND_g _17634_ (.A(_11899_), .B(_11900_), .Y(_00149_));
NAND_g _17635_ (.A(_11695_), .B(_11837_), .Y(_11901_));
NAND_g _17636_ (.A(cpuregs_18[31]), .B(_11838_), .Y(_11902_));
NAND_g _17637_ (.A(_11901_), .B(_11902_), .Y(_00150_));
AND_g _17638_ (.A(mem_state[0]), .B(mem_state[1]), .Y(_11903_));
AND_g _17639_ (.A(mem_do_rinst), .B(resetn), .Y(_11904_));
NAND_g _17640_ (.A(mem_do_rinst), .B(resetn), .Y(_11905_));
NAND_g _17641_ (.A(_11903_), .B(_11904_), .Y(_11906_));
NOR_g _17642_ (.A(mem_do_wdata), .B(mem_do_rdata), .Y(_11907_));
NOR_g _17643_ (.A(mem_do_rdata), .B(mem_do_rinst), .Y(_11908_));
NAND_g _17644_ (.A(_10893_), .B(_11908_), .Y(_11909_));
AND_g _17645_ (.A(mem_valid), .B(mem_ready), .Y(_11910_));
NAND_g _17646_ (.A(mem_valid), .B(mem_ready), .Y(_11911_));
NOR_g _17647_ (.A(mem_state[0]), .B(mem_state[1]), .Y(_11912_));
NAND_g _17648_ (.A(resetn), .B(_11910_), .Y(_11913_));
NOR_g _17649_ (.A(_11912_), .B(_11913_), .Y(_11914_));
NAND_g _17650_ (.A(_11909_), .B(_11914_), .Y(_11915_));
AND_g _17651_ (.A(_11906_), .B(_11915_), .Y(_11916_));
NOT_g _17652_ (.A(_11916_), .Y(_11917_));
NOR_g _17653_ (.A(_10898_), .B(_11916_), .Y(_11918_));
NAND_g _17654_ (.A(mem_do_rinst), .B(_11917_), .Y(_11919_));
NAND_g _17655_ (.A(mem_rdata[25]), .B(_11910_), .Y(_11920_));
NAND_g _17656_ (.A(mem_rdata_q[25]), .B(_11911_), .Y(_11921_));
NAND_g _17657_ (.A(_11920_), .B(_11921_), .Y(_00797_));
NAND_g _17658_ (.A(_11918_), .B(_00797_), .Y(_11922_));
NAND_g _17659_ (.A(decoded_imm_j[5]), .B(_11919_), .Y(_11923_));
NAND_g _17660_ (.A(_11922_), .B(_11923_), .Y(_00151_));
NAND_g _17661_ (.A(mem_rdata[28]), .B(_11910_), .Y(_11924_));
NAND_g _17662_ (.A(mem_rdata_q[28]), .B(_11911_), .Y(_11925_));
NAND_g _17663_ (.A(_11924_), .B(_11925_), .Y(_00800_));
NAND_g _17664_ (.A(_11918_), .B(_00800_), .Y(_11926_));
NAND_g _17665_ (.A(decoded_imm_j[8]), .B(_11919_), .Y(_11927_));
NAND_g _17666_ (.A(_11926_), .B(_11927_), .Y(_00152_));
NAND_g _17667_ (.A(mem_rdata[29]), .B(_11910_), .Y(_11928_));
NAND_g _17668_ (.A(mem_rdata_q[29]), .B(_11911_), .Y(_11929_));
NAND_g _17669_ (.A(_11928_), .B(_11929_), .Y(_00801_));
NAND_g _17670_ (.A(_11918_), .B(_00801_), .Y(_11930_));
NAND_g _17671_ (.A(decoded_imm_j[9]), .B(_11919_), .Y(_11931_));
NAND_g _17672_ (.A(_11930_), .B(_11931_), .Y(_00153_));
NOR_g _17673_ (.A(_11041_), .B(_11764_), .Y(_11932_));
AND_g _17674_ (.A(_11697_), .B(_11932_), .Y(_11933_));
NAND_g _17675_ (.A(_11697_), .B(_11932_), .Y(_11934_));
NAND_g _17676_ (.A(cpuregs_11[0]), .B(_11934_), .Y(_11935_));
NAND_g _17677_ (.A(_11301_), .B(_11933_), .Y(_11936_));
NAND_g _17678_ (.A(_11935_), .B(_11936_), .Y(_00154_));
NAND_g _17679_ (.A(cpuregs_11[1]), .B(_11934_), .Y(_11937_));
NAND_g _17680_ (.A(_11310_), .B(_11933_), .Y(_11938_));
NAND_g _17681_ (.A(_11937_), .B(_11938_), .Y(_00155_));
NAND_g _17682_ (.A(cpuregs_11[2]), .B(_11934_), .Y(_11939_));
NAND_g _17683_ (.A(_11319_), .B(_11933_), .Y(_11940_));
NAND_g _17684_ (.A(_11939_), .B(_11940_), .Y(_00156_));
NAND_g _17685_ (.A(cpuregs_11[3]), .B(_11934_), .Y(_11941_));
NAND_g _17686_ (.A(_11332_), .B(_11933_), .Y(_11942_));
NAND_g _17687_ (.A(_11941_), .B(_11942_), .Y(_00157_));
NAND_g _17688_ (.A(cpuregs_11[4]), .B(_11934_), .Y(_11943_));
NAND_g _17689_ (.A(_11345_), .B(_11933_), .Y(_11944_));
NAND_g _17690_ (.A(_11943_), .B(_11944_), .Y(_00158_));
NAND_g _17691_ (.A(cpuregs_11[5]), .B(_11934_), .Y(_11945_));
NAND_g _17692_ (.A(_11358_), .B(_11933_), .Y(_11946_));
NAND_g _17693_ (.A(_11945_), .B(_11946_), .Y(_00159_));
NAND_g _17694_ (.A(cpuregs_11[6]), .B(_11934_), .Y(_11947_));
NAND_g _17695_ (.A(_11371_), .B(_11933_), .Y(_11948_));
NAND_g _17696_ (.A(_11947_), .B(_11948_), .Y(_00160_));
NAND_g _17697_ (.A(cpuregs_11[7]), .B(_11934_), .Y(_11949_));
NAND_g _17698_ (.A(_11384_), .B(_11933_), .Y(_11950_));
NAND_g _17699_ (.A(_11949_), .B(_11950_), .Y(_00161_));
NAND_g _17700_ (.A(cpuregs_11[8]), .B(_11934_), .Y(_11951_));
NAND_g _17701_ (.A(_11397_), .B(_11933_), .Y(_11952_));
NAND_g _17702_ (.A(_11951_), .B(_11952_), .Y(_00162_));
NAND_g _17703_ (.A(cpuregs_11[9]), .B(_11934_), .Y(_11953_));
NAND_g _17704_ (.A(_11410_), .B(_11933_), .Y(_11954_));
NAND_g _17705_ (.A(_11953_), .B(_11954_), .Y(_00163_));
NAND_g _17706_ (.A(cpuregs_11[10]), .B(_11934_), .Y(_11955_));
NAND_g _17707_ (.A(_11423_), .B(_11933_), .Y(_11956_));
NAND_g _17708_ (.A(_11955_), .B(_11956_), .Y(_00164_));
NAND_g _17709_ (.A(cpuregs_11[11]), .B(_11934_), .Y(_11957_));
NAND_g _17710_ (.A(_11436_), .B(_11933_), .Y(_11958_));
NAND_g _17711_ (.A(_11957_), .B(_11958_), .Y(_00165_));
NAND_g _17712_ (.A(cpuregs_11[12]), .B(_11934_), .Y(_11959_));
NAND_g _17713_ (.A(_11449_), .B(_11933_), .Y(_11960_));
NAND_g _17714_ (.A(_11959_), .B(_11960_), .Y(_00166_));
NAND_g _17715_ (.A(cpuregs_11[13]), .B(_11934_), .Y(_11961_));
NAND_g _17716_ (.A(_11462_), .B(_11933_), .Y(_11962_));
NAND_g _17717_ (.A(_11961_), .B(_11962_), .Y(_00167_));
NAND_g _17718_ (.A(cpuregs_11[14]), .B(_11934_), .Y(_11963_));
NAND_g _17719_ (.A(_11475_), .B(_11933_), .Y(_11964_));
NAND_g _17720_ (.A(_11963_), .B(_11964_), .Y(_00168_));
NAND_g _17721_ (.A(cpuregs_11[15]), .B(_11934_), .Y(_11965_));
NAND_g _17722_ (.A(_11488_), .B(_11933_), .Y(_11966_));
NAND_g _17723_ (.A(_11965_), .B(_11966_), .Y(_00169_));
NOR_g _17724_ (.A(cpuregs_11[16]), .B(_11933_), .Y(_11967_));
NOR_g _17725_ (.A(_11501_), .B(_11934_), .Y(_11968_));
NOR_g _17726_ (.A(_11967_), .B(_11968_), .Y(_00170_));
NAND_g _17727_ (.A(_11514_), .B(_11933_), .Y(_11969_));
NAND_g _17728_ (.A(cpuregs_11[17]), .B(_11934_), .Y(_11970_));
NAND_g _17729_ (.A(_11969_), .B(_11970_), .Y(_00171_));
NAND_g _17730_ (.A(_11527_), .B(_11933_), .Y(_11971_));
NAND_g _17731_ (.A(cpuregs_11[18]), .B(_11934_), .Y(_11972_));
NAND_g _17732_ (.A(_11971_), .B(_11972_), .Y(_00172_));
NAND_g _17733_ (.A(_11540_), .B(_11933_), .Y(_11973_));
NAND_g _17734_ (.A(cpuregs_11[19]), .B(_11934_), .Y(_11974_));
NAND_g _17735_ (.A(_11973_), .B(_11974_), .Y(_00173_));
NAND_g _17736_ (.A(_11553_), .B(_11933_), .Y(_11975_));
NAND_g _17737_ (.A(cpuregs_11[20]), .B(_11934_), .Y(_11976_));
NAND_g _17738_ (.A(_11975_), .B(_11976_), .Y(_00174_));
NAND_g _17739_ (.A(_11566_), .B(_11933_), .Y(_11977_));
NAND_g _17740_ (.A(cpuregs_11[21]), .B(_11934_), .Y(_11978_));
NAND_g _17741_ (.A(_11977_), .B(_11978_), .Y(_00175_));
NAND_g _17742_ (.A(_11579_), .B(_11933_), .Y(_11979_));
NAND_g _17743_ (.A(cpuregs_11[22]), .B(_11934_), .Y(_11980_));
NAND_g _17744_ (.A(_11979_), .B(_11980_), .Y(_00176_));
NAND_g _17745_ (.A(_11592_), .B(_11933_), .Y(_11981_));
NAND_g _17746_ (.A(cpuregs_11[23]), .B(_11934_), .Y(_11982_));
NAND_g _17747_ (.A(_11981_), .B(_11982_), .Y(_00177_));
NAND_g _17748_ (.A(_11605_), .B(_11933_), .Y(_11983_));
NAND_g _17749_ (.A(cpuregs_11[24]), .B(_11934_), .Y(_11984_));
NAND_g _17750_ (.A(_11983_), .B(_11984_), .Y(_00178_));
NAND_g _17751_ (.A(_11618_), .B(_11933_), .Y(_11985_));
NAND_g _17752_ (.A(cpuregs_11[25]), .B(_11934_), .Y(_11986_));
NAND_g _17753_ (.A(_11985_), .B(_11986_), .Y(_00179_));
NAND_g _17754_ (.A(_11631_), .B(_11933_), .Y(_11987_));
NAND_g _17755_ (.A(cpuregs_11[26]), .B(_11934_), .Y(_11988_));
NAND_g _17756_ (.A(_11987_), .B(_11988_), .Y(_00180_));
NAND_g _17757_ (.A(_11644_), .B(_11933_), .Y(_11989_));
NAND_g _17758_ (.A(cpuregs_11[27]), .B(_11934_), .Y(_11990_));
NAND_g _17759_ (.A(_11989_), .B(_11990_), .Y(_00181_));
NAND_g _17760_ (.A(_11657_), .B(_11933_), .Y(_11991_));
NAND_g _17761_ (.A(cpuregs_11[28]), .B(_11934_), .Y(_11992_));
NAND_g _17762_ (.A(_11991_), .B(_11992_), .Y(_00182_));
NAND_g _17763_ (.A(_11670_), .B(_11933_), .Y(_11993_));
NAND_g _17764_ (.A(cpuregs_11[29]), .B(_11934_), .Y(_11994_));
NAND_g _17765_ (.A(_11993_), .B(_11994_), .Y(_00183_));
NAND_g _17766_ (.A(_11683_), .B(_11933_), .Y(_11995_));
NAND_g _17767_ (.A(cpuregs_11[30]), .B(_11934_), .Y(_11996_));
NAND_g _17768_ (.A(_11995_), .B(_11996_), .Y(_00184_));
NAND_g _17769_ (.A(_11695_), .B(_11933_), .Y(_11997_));
NAND_g _17770_ (.A(cpuregs_11[31]), .B(_11934_), .Y(_11998_));
NAND_g _17771_ (.A(_11997_), .B(_11998_), .Y(_00185_));
AND_g _17772_ (.A(_11042_), .B(latched_rd[3]), .Y(_11999_));
AND_g _17773_ (.A(_11766_), .B(_11999_), .Y(_12000_));
AND_g _17774_ (.A(latched_rd[3]), .B(_11766_), .Y(_12001_));
AND_g _17775_ (.A(_11042_), .B(_12001_), .Y(_12002_));
AND_g _17776_ (.A(_11289_), .B(_12002_), .Y(_12003_));
NAND_g _17777_ (.A(_11289_), .B(_12002_), .Y(_12004_));
NAND_g _17778_ (.A(cpuregs_25[0]), .B(_12004_), .Y(_12005_));
NAND_g _17779_ (.A(_11301_), .B(_12003_), .Y(_12006_));
AND_g _17780_ (.A(_11289_), .B(_12000_), .Y(_12007_));
NAND_g _17781_ (.A(_11289_), .B(_12000_), .Y(_12008_));
NAND_g _17782_ (.A(_12005_), .B(_12006_), .Y(_00186_));
NAND_g _17783_ (.A(cpuregs_25[1]), .B(_12004_), .Y(_12009_));
NAND_g _17784_ (.A(_11310_), .B(_12003_), .Y(_12010_));
NAND_g _17785_ (.A(_12009_), .B(_12010_), .Y(_00187_));
NAND_g _17786_ (.A(cpuregs_25[2]), .B(_12004_), .Y(_12011_));
NAND_g _17787_ (.A(_11319_), .B(_12003_), .Y(_12012_));
NAND_g _17788_ (.A(_12011_), .B(_12012_), .Y(_00188_));
NAND_g _17789_ (.A(cpuregs_25[3]), .B(_12004_), .Y(_12013_));
NAND_g _17790_ (.A(_11332_), .B(_12003_), .Y(_12014_));
NAND_g _17791_ (.A(_12013_), .B(_12014_), .Y(_00189_));
NAND_g _17792_ (.A(cpuregs_25[4]), .B(_12004_), .Y(_12015_));
NAND_g _17793_ (.A(_11345_), .B(_12003_), .Y(_12016_));
NAND_g _17794_ (.A(_12015_), .B(_12016_), .Y(_00190_));
NAND_g _17795_ (.A(cpuregs_25[5]), .B(_12004_), .Y(_12017_));
NAND_g _17796_ (.A(_11358_), .B(_12003_), .Y(_12018_));
NAND_g _17797_ (.A(_12017_), .B(_12018_), .Y(_00191_));
NAND_g _17798_ (.A(cpuregs_25[6]), .B(_12004_), .Y(_12019_));
NAND_g _17799_ (.A(_11371_), .B(_12003_), .Y(_12020_));
NAND_g _17800_ (.A(_12019_), .B(_12020_), .Y(_00192_));
NAND_g _17801_ (.A(cpuregs_25[7]), .B(_12004_), .Y(_12021_));
NAND_g _17802_ (.A(_11384_), .B(_12003_), .Y(_12022_));
NAND_g _17803_ (.A(_12021_), .B(_12022_), .Y(_00193_));
NAND_g _17804_ (.A(cpuregs_25[8]), .B(_12004_), .Y(_12023_));
NAND_g _17805_ (.A(_11397_), .B(_12003_), .Y(_12024_));
NAND_g _17806_ (.A(_12023_), .B(_12024_), .Y(_00194_));
NAND_g _17807_ (.A(cpuregs_25[9]), .B(_12004_), .Y(_12025_));
NAND_g _17808_ (.A(_11410_), .B(_12003_), .Y(_12026_));
NAND_g _17809_ (.A(_12025_), .B(_12026_), .Y(_00195_));
NAND_g _17810_ (.A(cpuregs_25[10]), .B(_12004_), .Y(_12027_));
NAND_g _17811_ (.A(_11423_), .B(_12003_), .Y(_12028_));
NAND_g _17812_ (.A(_12027_), .B(_12028_), .Y(_00196_));
NAND_g _17813_ (.A(cpuregs_25[11]), .B(_12004_), .Y(_12029_));
NAND_g _17814_ (.A(_11436_), .B(_12003_), .Y(_12030_));
NAND_g _17815_ (.A(_12029_), .B(_12030_), .Y(_00197_));
NAND_g _17816_ (.A(cpuregs_25[12]), .B(_12004_), .Y(_12031_));
NAND_g _17817_ (.A(_11449_), .B(_12003_), .Y(_12032_));
NAND_g _17818_ (.A(_12031_), .B(_12032_), .Y(_00198_));
NAND_g _17819_ (.A(cpuregs_25[13]), .B(_12004_), .Y(_12033_));
NAND_g _17820_ (.A(_11462_), .B(_12003_), .Y(_12034_));
NAND_g _17821_ (.A(_12033_), .B(_12034_), .Y(_00199_));
NAND_g _17822_ (.A(cpuregs_25[14]), .B(_12004_), .Y(_12035_));
NAND_g _17823_ (.A(_11475_), .B(_12003_), .Y(_12036_));
NAND_g _17824_ (.A(_12035_), .B(_12036_), .Y(_00200_));
NAND_g _17825_ (.A(cpuregs_25[15]), .B(_12004_), .Y(_12037_));
NAND_g _17826_ (.A(_11488_), .B(_12003_), .Y(_12038_));
NAND_g _17827_ (.A(_12037_), .B(_12038_), .Y(_00201_));
NAND_g _17828_ (.A(cpuregs_25[16]), .B(_12004_), .Y(_12039_));
NAND_g _17829_ (.A(_11501_), .B(_12003_), .Y(_12040_));
NAND_g _17830_ (.A(_12039_), .B(_12040_), .Y(_00202_));
NAND_g _17831_ (.A(cpuregs_25[17]), .B(_12008_), .Y(_12041_));
NAND_g _17832_ (.A(_11514_), .B(_12007_), .Y(_12042_));
NAND_g _17833_ (.A(_12041_), .B(_12042_), .Y(_00203_));
NAND_g _17834_ (.A(cpuregs_25[18]), .B(_12008_), .Y(_12043_));
NAND_g _17835_ (.A(_11527_), .B(_12007_), .Y(_12044_));
NAND_g _17836_ (.A(_12043_), .B(_12044_), .Y(_00204_));
NAND_g _17837_ (.A(cpuregs_25[19]), .B(_12008_), .Y(_12045_));
NAND_g _17838_ (.A(_11540_), .B(_12007_), .Y(_12046_));
NAND_g _17839_ (.A(_12045_), .B(_12046_), .Y(_00205_));
NAND_g _17840_ (.A(cpuregs_25[20]), .B(_12008_), .Y(_12047_));
NAND_g _17841_ (.A(_11553_), .B(_12007_), .Y(_12048_));
NAND_g _17842_ (.A(_12047_), .B(_12048_), .Y(_00206_));
NAND_g _17843_ (.A(cpuregs_25[21]), .B(_12008_), .Y(_12049_));
NAND_g _17844_ (.A(_11566_), .B(_12007_), .Y(_12050_));
NAND_g _17845_ (.A(_12049_), .B(_12050_), .Y(_00207_));
NAND_g _17846_ (.A(cpuregs_25[22]), .B(_12008_), .Y(_12051_));
NAND_g _17847_ (.A(_11579_), .B(_12007_), .Y(_12052_));
NAND_g _17848_ (.A(_12051_), .B(_12052_), .Y(_00208_));
NAND_g _17849_ (.A(cpuregs_25[23]), .B(_12008_), .Y(_12053_));
NAND_g _17850_ (.A(_11592_), .B(_12007_), .Y(_12054_));
NAND_g _17851_ (.A(_12053_), .B(_12054_), .Y(_00209_));
NAND_g _17852_ (.A(cpuregs_25[24]), .B(_12008_), .Y(_12055_));
NAND_g _17853_ (.A(_11605_), .B(_12007_), .Y(_12056_));
NAND_g _17854_ (.A(_12055_), .B(_12056_), .Y(_00210_));
NAND_g _17855_ (.A(cpuregs_25[25]), .B(_12008_), .Y(_12057_));
NAND_g _17856_ (.A(_11618_), .B(_12007_), .Y(_12058_));
NAND_g _17857_ (.A(_12057_), .B(_12058_), .Y(_00211_));
NAND_g _17858_ (.A(cpuregs_25[26]), .B(_12008_), .Y(_12059_));
NAND_g _17859_ (.A(_11631_), .B(_12007_), .Y(_12060_));
NAND_g _17860_ (.A(_12059_), .B(_12060_), .Y(_00212_));
NAND_g _17861_ (.A(cpuregs_25[27]), .B(_12008_), .Y(_12061_));
NAND_g _17862_ (.A(_11644_), .B(_12007_), .Y(_12062_));
NAND_g _17863_ (.A(_12061_), .B(_12062_), .Y(_00213_));
NAND_g _17864_ (.A(cpuregs_25[28]), .B(_12008_), .Y(_12063_));
NAND_g _17865_ (.A(_11657_), .B(_12007_), .Y(_12064_));
NAND_g _17866_ (.A(_12063_), .B(_12064_), .Y(_00214_));
NAND_g _17867_ (.A(cpuregs_25[29]), .B(_12008_), .Y(_12065_));
NAND_g _17868_ (.A(_11670_), .B(_12007_), .Y(_12066_));
NAND_g _17869_ (.A(_12065_), .B(_12066_), .Y(_00215_));
NAND_g _17870_ (.A(cpuregs_25[30]), .B(_12008_), .Y(_12067_));
NAND_g _17871_ (.A(_11683_), .B(_12007_), .Y(_12068_));
NAND_g _17872_ (.A(_12067_), .B(_12068_), .Y(_00216_));
NAND_g _17873_ (.A(cpuregs_25[31]), .B(_12008_), .Y(_12069_));
NAND_g _17874_ (.A(_11695_), .B(_12007_), .Y(_12070_));
NAND_g _17875_ (.A(_12069_), .B(_12070_), .Y(_00217_));
AND_g _17876_ (.A(_11278_), .B(_11768_), .Y(_12071_));
NAND_g _17877_ (.A(_11278_), .B(_11768_), .Y(_12072_));
NAND_g _17878_ (.A(_11301_), .B(_12071_), .Y(_12073_));
NAND_g _17879_ (.A(cpuregs_4[0]), .B(_12072_), .Y(_12074_));
AND_g _17880_ (.A(_11288_), .B(_11764_), .Y(_12075_));
NAND_g _17881_ (.A(_12073_), .B(_12074_), .Y(_00218_));
NAND_g _17882_ (.A(_11310_), .B(_12071_), .Y(_12076_));
NAND_g _17883_ (.A(cpuregs_4[1]), .B(_12072_), .Y(_12077_));
NAND_g _17884_ (.A(_12076_), .B(_12077_), .Y(_00219_));
NAND_g _17885_ (.A(_11319_), .B(_12071_), .Y(_12078_));
NAND_g _17886_ (.A(cpuregs_4[2]), .B(_12072_), .Y(_12079_));
NAND_g _17887_ (.A(_12078_), .B(_12079_), .Y(_00220_));
NAND_g _17888_ (.A(_11332_), .B(_12071_), .Y(_12080_));
NAND_g _17889_ (.A(cpuregs_4[3]), .B(_12072_), .Y(_12081_));
NAND_g _17890_ (.A(_12080_), .B(_12081_), .Y(_00221_));
NAND_g _17891_ (.A(_11345_), .B(_12071_), .Y(_12082_));
NAND_g _17892_ (.A(cpuregs_4[4]), .B(_12072_), .Y(_12083_));
NAND_g _17893_ (.A(_12082_), .B(_12083_), .Y(_00222_));
NAND_g _17894_ (.A(_11358_), .B(_12071_), .Y(_12084_));
NAND_g _17895_ (.A(cpuregs_4[5]), .B(_12072_), .Y(_12085_));
NAND_g _17896_ (.A(_12084_), .B(_12085_), .Y(_00223_));
NAND_g _17897_ (.A(_11371_), .B(_12071_), .Y(_12086_));
NAND_g _17898_ (.A(cpuregs_4[6]), .B(_12072_), .Y(_12087_));
NAND_g _17899_ (.A(_12086_), .B(_12087_), .Y(_00224_));
NAND_g _17900_ (.A(_11384_), .B(_12071_), .Y(_12088_));
NAND_g _17901_ (.A(cpuregs_4[7]), .B(_12072_), .Y(_12089_));
NAND_g _17902_ (.A(_12088_), .B(_12089_), .Y(_00225_));
NAND_g _17903_ (.A(_11397_), .B(_12071_), .Y(_12090_));
NAND_g _17904_ (.A(cpuregs_4[8]), .B(_12072_), .Y(_12091_));
NAND_g _17905_ (.A(_12090_), .B(_12091_), .Y(_00226_));
NAND_g _17906_ (.A(_11410_), .B(_12071_), .Y(_12092_));
NAND_g _17907_ (.A(cpuregs_4[9]), .B(_12072_), .Y(_12093_));
NAND_g _17908_ (.A(_12092_), .B(_12093_), .Y(_00227_));
NAND_g _17909_ (.A(_11423_), .B(_12071_), .Y(_12094_));
NAND_g _17910_ (.A(cpuregs_4[10]), .B(_12072_), .Y(_12095_));
NAND_g _17911_ (.A(_12094_), .B(_12095_), .Y(_00228_));
NAND_g _17912_ (.A(_11436_), .B(_12071_), .Y(_12096_));
NAND_g _17913_ (.A(cpuregs_4[11]), .B(_12072_), .Y(_12097_));
NAND_g _17914_ (.A(_12096_), .B(_12097_), .Y(_00229_));
NAND_g _17915_ (.A(_11449_), .B(_12071_), .Y(_12098_));
NAND_g _17916_ (.A(cpuregs_4[12]), .B(_12072_), .Y(_12099_));
NAND_g _17917_ (.A(_12098_), .B(_12099_), .Y(_00230_));
NAND_g _17918_ (.A(_11462_), .B(_12071_), .Y(_12100_));
NAND_g _17919_ (.A(cpuregs_4[13]), .B(_12072_), .Y(_12101_));
NAND_g _17920_ (.A(_12100_), .B(_12101_), .Y(_00231_));
NAND_g _17921_ (.A(_11475_), .B(_12071_), .Y(_12102_));
NAND_g _17922_ (.A(cpuregs_4[14]), .B(_12072_), .Y(_12103_));
NAND_g _17923_ (.A(_12102_), .B(_12103_), .Y(_00232_));
NAND_g _17924_ (.A(_11488_), .B(_12071_), .Y(_12104_));
NAND_g _17925_ (.A(cpuregs_4[15]), .B(_12072_), .Y(_12105_));
NAND_g _17926_ (.A(_12104_), .B(_12105_), .Y(_00233_));
NAND_g _17927_ (.A(_11501_), .B(_12071_), .Y(_12106_));
NAND_g _17928_ (.A(cpuregs_4[16]), .B(_12072_), .Y(_12107_));
NAND_g _17929_ (.A(_12106_), .B(_12107_), .Y(_00234_));
NOR_g _17930_ (.A(cpuregs_4[17]), .B(_12071_), .Y(_12108_));
NOR_g _17931_ (.A(_11514_), .B(_12072_), .Y(_12109_));
NOR_g _17932_ (.A(_12108_), .B(_12109_), .Y(_00235_));
NAND_g _17933_ (.A(cpuregs_4[18]), .B(_12072_), .Y(_12110_));
NAND_g _17934_ (.A(_11527_), .B(_12071_), .Y(_12111_));
NAND_g _17935_ (.A(_12110_), .B(_12111_), .Y(_00236_));
NAND_g _17936_ (.A(cpuregs_4[19]), .B(_12072_), .Y(_12112_));
NAND_g _17937_ (.A(_11540_), .B(_12071_), .Y(_12113_));
NAND_g _17938_ (.A(_12112_), .B(_12113_), .Y(_00237_));
NAND_g _17939_ (.A(cpuregs_4[20]), .B(_12072_), .Y(_12114_));
NAND_g _17940_ (.A(_11553_), .B(_12071_), .Y(_12115_));
NAND_g _17941_ (.A(_12114_), .B(_12115_), .Y(_00238_));
NAND_g _17942_ (.A(cpuregs_4[21]), .B(_12072_), .Y(_12116_));
NAND_g _17943_ (.A(_11566_), .B(_12071_), .Y(_12117_));
NAND_g _17944_ (.A(_12116_), .B(_12117_), .Y(_00239_));
NAND_g _17945_ (.A(cpuregs_4[22]), .B(_12072_), .Y(_12118_));
NAND_g _17946_ (.A(_11579_), .B(_12071_), .Y(_12119_));
NAND_g _17947_ (.A(_12118_), .B(_12119_), .Y(_00240_));
NAND_g _17948_ (.A(cpuregs_4[23]), .B(_12072_), .Y(_12120_));
NAND_g _17949_ (.A(_11592_), .B(_12071_), .Y(_12121_));
NAND_g _17950_ (.A(_12120_), .B(_12121_), .Y(_00241_));
NAND_g _17951_ (.A(cpuregs_4[24]), .B(_12072_), .Y(_12122_));
NAND_g _17952_ (.A(_11605_), .B(_12071_), .Y(_12123_));
NAND_g _17953_ (.A(_12122_), .B(_12123_), .Y(_00242_));
NAND_g _17954_ (.A(cpuregs_4[25]), .B(_12072_), .Y(_12124_));
NAND_g _17955_ (.A(_11618_), .B(_12071_), .Y(_12125_));
NAND_g _17956_ (.A(_12124_), .B(_12125_), .Y(_00243_));
NAND_g _17957_ (.A(cpuregs_4[26]), .B(_12072_), .Y(_12126_));
NAND_g _17958_ (.A(_11631_), .B(_12071_), .Y(_12127_));
NAND_g _17959_ (.A(_12126_), .B(_12127_), .Y(_00244_));
NAND_g _17960_ (.A(cpuregs_4[27]), .B(_12072_), .Y(_12128_));
NAND_g _17961_ (.A(_11644_), .B(_12071_), .Y(_12129_));
NAND_g _17962_ (.A(_12128_), .B(_12129_), .Y(_00245_));
NAND_g _17963_ (.A(cpuregs_4[28]), .B(_12072_), .Y(_12130_));
NAND_g _17964_ (.A(_11657_), .B(_12071_), .Y(_12131_));
NAND_g _17965_ (.A(_12130_), .B(_12131_), .Y(_00246_));
NAND_g _17966_ (.A(cpuregs_4[29]), .B(_12072_), .Y(_12132_));
NAND_g _17967_ (.A(_11670_), .B(_12071_), .Y(_12133_));
NAND_g _17968_ (.A(_12132_), .B(_12133_), .Y(_00247_));
NAND_g _17969_ (.A(cpuregs_4[30]), .B(_12072_), .Y(_12134_));
NAND_g _17970_ (.A(_11683_), .B(_12071_), .Y(_12135_));
NAND_g _17971_ (.A(_12134_), .B(_12135_), .Y(_00248_));
NAND_g _17972_ (.A(cpuregs_4[31]), .B(_12072_), .Y(_12136_));
NAND_g _17973_ (.A(_11695_), .B(_12071_), .Y(_12137_));
NAND_g _17974_ (.A(_12136_), .B(_12137_), .Y(_00249_));
AND_g _17975_ (.A(_11289_), .B(_11836_), .Y(_12138_));
NAND_g _17976_ (.A(_11289_), .B(_11836_), .Y(_12139_));
NAND_g _17977_ (.A(cpuregs_17[0]), .B(_12139_), .Y(_12140_));
NAND_g _17978_ (.A(_11301_), .B(_12138_), .Y(_12141_));
NAND_g _17979_ (.A(_12140_), .B(_12141_), .Y(_00250_));
NAND_g _17980_ (.A(cpuregs_17[1]), .B(_12139_), .Y(_12142_));
NAND_g _17981_ (.A(_11310_), .B(_12138_), .Y(_12143_));
NAND_g _17982_ (.A(_12142_), .B(_12143_), .Y(_00251_));
NAND_g _17983_ (.A(cpuregs_17[2]), .B(_12139_), .Y(_12144_));
NAND_g _17984_ (.A(_11319_), .B(_12138_), .Y(_12145_));
NAND_g _17985_ (.A(_12144_), .B(_12145_), .Y(_00252_));
NAND_g _17986_ (.A(cpuregs_17[3]), .B(_12139_), .Y(_12146_));
NAND_g _17987_ (.A(_11332_), .B(_12138_), .Y(_12147_));
NAND_g _17988_ (.A(_12146_), .B(_12147_), .Y(_00253_));
NAND_g _17989_ (.A(cpuregs_17[4]), .B(_12139_), .Y(_12148_));
NAND_g _17990_ (.A(_11345_), .B(_12138_), .Y(_12149_));
NAND_g _17991_ (.A(_12148_), .B(_12149_), .Y(_00254_));
NAND_g _17992_ (.A(cpuregs_17[5]), .B(_12139_), .Y(_12150_));
NAND_g _17993_ (.A(_11358_), .B(_12138_), .Y(_12151_));
NAND_g _17994_ (.A(_12150_), .B(_12151_), .Y(_00255_));
NAND_g _17995_ (.A(cpuregs_17[6]), .B(_12139_), .Y(_12152_));
NAND_g _17996_ (.A(_11371_), .B(_12138_), .Y(_12153_));
NAND_g _17997_ (.A(_12152_), .B(_12153_), .Y(_00256_));
NAND_g _17998_ (.A(cpuregs_17[7]), .B(_12139_), .Y(_12154_));
NAND_g _17999_ (.A(_11384_), .B(_12138_), .Y(_12155_));
NAND_g _18000_ (.A(_12154_), .B(_12155_), .Y(_00257_));
NAND_g _18001_ (.A(cpuregs_17[8]), .B(_12139_), .Y(_12156_));
NAND_g _18002_ (.A(_11397_), .B(_12138_), .Y(_12157_));
NAND_g _18003_ (.A(_12156_), .B(_12157_), .Y(_00258_));
NAND_g _18004_ (.A(cpuregs_17[9]), .B(_12139_), .Y(_12158_));
NAND_g _18005_ (.A(_11410_), .B(_12138_), .Y(_12159_));
NAND_g _18006_ (.A(_12158_), .B(_12159_), .Y(_00259_));
NAND_g _18007_ (.A(cpuregs_17[10]), .B(_12139_), .Y(_12160_));
NAND_g _18008_ (.A(_11423_), .B(_12138_), .Y(_12161_));
NAND_g _18009_ (.A(_12160_), .B(_12161_), .Y(_00260_));
NAND_g _18010_ (.A(cpuregs_17[11]), .B(_12139_), .Y(_12162_));
NAND_g _18011_ (.A(_11436_), .B(_12138_), .Y(_12163_));
NAND_g _18012_ (.A(_12162_), .B(_12163_), .Y(_00261_));
NAND_g _18013_ (.A(cpuregs_17[12]), .B(_12139_), .Y(_12164_));
NAND_g _18014_ (.A(_11449_), .B(_12138_), .Y(_12165_));
NAND_g _18015_ (.A(_12164_), .B(_12165_), .Y(_00262_));
NAND_g _18016_ (.A(cpuregs_17[13]), .B(_12139_), .Y(_12166_));
NAND_g _18017_ (.A(_11462_), .B(_12138_), .Y(_12167_));
NAND_g _18018_ (.A(_12166_), .B(_12167_), .Y(_00263_));
NAND_g _18019_ (.A(cpuregs_17[14]), .B(_12139_), .Y(_12168_));
NAND_g _18020_ (.A(_11475_), .B(_12138_), .Y(_12169_));
NAND_g _18021_ (.A(_12168_), .B(_12169_), .Y(_00264_));
NAND_g _18022_ (.A(cpuregs_17[15]), .B(_12139_), .Y(_12170_));
NAND_g _18023_ (.A(_11488_), .B(_12138_), .Y(_12171_));
NAND_g _18024_ (.A(_12170_), .B(_12171_), .Y(_00265_));
NAND_g _18025_ (.A(cpuregs_17[16]), .B(_12139_), .Y(_12172_));
NAND_g _18026_ (.A(_11501_), .B(_12138_), .Y(_12173_));
NAND_g _18027_ (.A(_12172_), .B(_12173_), .Y(_00266_));
NOR_g _18028_ (.A(cpuregs_17[17]), .B(_12138_), .Y(_12174_));
NOR_g _18029_ (.A(_11514_), .B(_12139_), .Y(_12175_));
NOR_g _18030_ (.A(_12174_), .B(_12175_), .Y(_00267_));
NAND_g _18031_ (.A(cpuregs_17[18]), .B(_12139_), .Y(_12176_));
NAND_g _18032_ (.A(_11527_), .B(_12138_), .Y(_12177_));
NAND_g _18033_ (.A(_12176_), .B(_12177_), .Y(_00268_));
NAND_g _18034_ (.A(cpuregs_17[19]), .B(_12139_), .Y(_12178_));
NAND_g _18035_ (.A(_11540_), .B(_12138_), .Y(_12179_));
NAND_g _18036_ (.A(_12178_), .B(_12179_), .Y(_00269_));
NAND_g _18037_ (.A(cpuregs_17[20]), .B(_12139_), .Y(_12180_));
NAND_g _18038_ (.A(_11553_), .B(_12138_), .Y(_12181_));
NAND_g _18039_ (.A(_12180_), .B(_12181_), .Y(_00270_));
NAND_g _18040_ (.A(cpuregs_17[21]), .B(_12139_), .Y(_12182_));
NAND_g _18041_ (.A(_11566_), .B(_12138_), .Y(_12183_));
NAND_g _18042_ (.A(_12182_), .B(_12183_), .Y(_00271_));
NAND_g _18043_ (.A(cpuregs_17[22]), .B(_12139_), .Y(_12184_));
NAND_g _18044_ (.A(_11579_), .B(_12138_), .Y(_12185_));
NAND_g _18045_ (.A(_12184_), .B(_12185_), .Y(_00272_));
NAND_g _18046_ (.A(cpuregs_17[23]), .B(_12139_), .Y(_12186_));
NAND_g _18047_ (.A(_11592_), .B(_12138_), .Y(_12187_));
NAND_g _18048_ (.A(_12186_), .B(_12187_), .Y(_00273_));
NAND_g _18049_ (.A(cpuregs_17[24]), .B(_12139_), .Y(_12188_));
NAND_g _18050_ (.A(_11605_), .B(_12138_), .Y(_12189_));
NAND_g _18051_ (.A(_12188_), .B(_12189_), .Y(_00274_));
NAND_g _18052_ (.A(cpuregs_17[25]), .B(_12139_), .Y(_12190_));
NAND_g _18053_ (.A(_11618_), .B(_12138_), .Y(_12191_));
NAND_g _18054_ (.A(_12190_), .B(_12191_), .Y(_00275_));
NAND_g _18055_ (.A(cpuregs_17[26]), .B(_12139_), .Y(_12192_));
NAND_g _18056_ (.A(_11631_), .B(_12138_), .Y(_12193_));
NAND_g _18057_ (.A(_12192_), .B(_12193_), .Y(_00276_));
NAND_g _18058_ (.A(cpuregs_17[27]), .B(_12139_), .Y(_12194_));
NAND_g _18059_ (.A(_11644_), .B(_12138_), .Y(_12195_));
NAND_g _18060_ (.A(_12194_), .B(_12195_), .Y(_00277_));
NAND_g _18061_ (.A(cpuregs_17[28]), .B(_12139_), .Y(_12196_));
NAND_g _18062_ (.A(_11657_), .B(_12138_), .Y(_12197_));
NAND_g _18063_ (.A(_12196_), .B(_12197_), .Y(_00278_));
NAND_g _18064_ (.A(cpuregs_17[29]), .B(_12139_), .Y(_12198_));
NAND_g _18065_ (.A(_11670_), .B(_12138_), .Y(_12199_));
NAND_g _18066_ (.A(_12198_), .B(_12199_), .Y(_00279_));
NAND_g _18067_ (.A(cpuregs_17[30]), .B(_12139_), .Y(_12200_));
NAND_g _18068_ (.A(_11683_), .B(_12138_), .Y(_12201_));
NAND_g _18069_ (.A(_12200_), .B(_12201_), .Y(_00280_));
NAND_g _18070_ (.A(cpuregs_17[31]), .B(_12139_), .Y(_12202_));
NAND_g _18071_ (.A(_11695_), .B(_12138_), .Y(_12203_));
NAND_g _18072_ (.A(_12202_), .B(_12203_), .Y(_00281_));
AND_g _18073_ (.A(_11932_), .B(_12000_), .Y(_12204_));
NAND_g _18074_ (.A(_11932_), .B(_12000_), .Y(_12205_));
NAND_g _18075_ (.A(cpuregs_27[0]), .B(_12205_), .Y(_12206_));
NAND_g _18076_ (.A(_11301_), .B(_12204_), .Y(_12207_));
NAND_g _18077_ (.A(_12206_), .B(_12207_), .Y(_00282_));
NAND_g _18078_ (.A(cpuregs_27[1]), .B(_12205_), .Y(_12208_));
NAND_g _18079_ (.A(_11310_), .B(_12204_), .Y(_12209_));
NAND_g _18080_ (.A(_12208_), .B(_12209_), .Y(_00283_));
NAND_g _18081_ (.A(cpuregs_27[2]), .B(_12205_), .Y(_12210_));
NAND_g _18082_ (.A(_11319_), .B(_12204_), .Y(_12211_));
NAND_g _18083_ (.A(_12210_), .B(_12211_), .Y(_00284_));
NAND_g _18084_ (.A(cpuregs_27[3]), .B(_12205_), .Y(_12212_));
NAND_g _18085_ (.A(_11332_), .B(_12204_), .Y(_12213_));
NAND_g _18086_ (.A(_12212_), .B(_12213_), .Y(_00285_));
NAND_g _18087_ (.A(cpuregs_27[4]), .B(_12205_), .Y(_12214_));
NAND_g _18088_ (.A(_11345_), .B(_12204_), .Y(_12215_));
NAND_g _18089_ (.A(_12214_), .B(_12215_), .Y(_00286_));
NAND_g _18090_ (.A(cpuregs_27[5]), .B(_12205_), .Y(_12216_));
NAND_g _18091_ (.A(_11358_), .B(_12204_), .Y(_12217_));
NAND_g _18092_ (.A(_12216_), .B(_12217_), .Y(_00287_));
NAND_g _18093_ (.A(cpuregs_27[6]), .B(_12205_), .Y(_12218_));
NAND_g _18094_ (.A(_11371_), .B(_12204_), .Y(_12219_));
NAND_g _18095_ (.A(_12218_), .B(_12219_), .Y(_00288_));
NAND_g _18096_ (.A(cpuregs_27[7]), .B(_12205_), .Y(_12220_));
NAND_g _18097_ (.A(_11384_), .B(_12204_), .Y(_12221_));
NAND_g _18098_ (.A(_12220_), .B(_12221_), .Y(_00289_));
NAND_g _18099_ (.A(cpuregs_27[8]), .B(_12205_), .Y(_12222_));
NAND_g _18100_ (.A(_11397_), .B(_12204_), .Y(_12223_));
NAND_g _18101_ (.A(_12222_), .B(_12223_), .Y(_00290_));
NAND_g _18102_ (.A(cpuregs_27[9]), .B(_12205_), .Y(_12224_));
NAND_g _18103_ (.A(_11410_), .B(_12204_), .Y(_12225_));
NAND_g _18104_ (.A(_12224_), .B(_12225_), .Y(_00291_));
NAND_g _18105_ (.A(cpuregs_27[10]), .B(_12205_), .Y(_12226_));
NAND_g _18106_ (.A(_11423_), .B(_12204_), .Y(_12227_));
NAND_g _18107_ (.A(_12226_), .B(_12227_), .Y(_00292_));
NAND_g _18108_ (.A(cpuregs_27[11]), .B(_12205_), .Y(_12228_));
NAND_g _18109_ (.A(_11436_), .B(_12204_), .Y(_12229_));
NAND_g _18110_ (.A(_12228_), .B(_12229_), .Y(_00293_));
NAND_g _18111_ (.A(cpuregs_27[12]), .B(_12205_), .Y(_12230_));
NAND_g _18112_ (.A(_11449_), .B(_12204_), .Y(_12231_));
NAND_g _18113_ (.A(_12230_), .B(_12231_), .Y(_00294_));
NAND_g _18114_ (.A(cpuregs_27[13]), .B(_12205_), .Y(_12232_));
NAND_g _18115_ (.A(_11462_), .B(_12204_), .Y(_12233_));
NAND_g _18116_ (.A(_12232_), .B(_12233_), .Y(_00295_));
NAND_g _18117_ (.A(cpuregs_27[14]), .B(_12205_), .Y(_12234_));
NAND_g _18118_ (.A(_11475_), .B(_12204_), .Y(_12235_));
NAND_g _18119_ (.A(_12234_), .B(_12235_), .Y(_00296_));
NAND_g _18120_ (.A(cpuregs_27[15]), .B(_12205_), .Y(_12236_));
NAND_g _18121_ (.A(_11488_), .B(_12204_), .Y(_12237_));
NAND_g _18122_ (.A(_12236_), .B(_12237_), .Y(_00297_));
NAND_g _18123_ (.A(cpuregs_27[16]), .B(_12205_), .Y(_12238_));
NAND_g _18124_ (.A(_11501_), .B(_12204_), .Y(_12239_));
NAND_g _18125_ (.A(_12238_), .B(_12239_), .Y(_00298_));
NAND_g _18126_ (.A(_11514_), .B(_12204_), .Y(_12240_));
NAND_g _18127_ (.A(cpuregs_27[17]), .B(_12205_), .Y(_12241_));
NAND_g _18128_ (.A(_12240_), .B(_12241_), .Y(_00299_));
NAND_g _18129_ (.A(_11527_), .B(_12204_), .Y(_12242_));
NAND_g _18130_ (.A(cpuregs_27[18]), .B(_12205_), .Y(_12243_));
NAND_g _18131_ (.A(_12242_), .B(_12243_), .Y(_00300_));
NAND_g _18132_ (.A(_11540_), .B(_12204_), .Y(_12244_));
NAND_g _18133_ (.A(cpuregs_27[19]), .B(_12205_), .Y(_12245_));
NAND_g _18134_ (.A(_12244_), .B(_12245_), .Y(_00301_));
NAND_g _18135_ (.A(_11553_), .B(_12204_), .Y(_12246_));
NAND_g _18136_ (.A(cpuregs_27[20]), .B(_12205_), .Y(_12247_));
NAND_g _18137_ (.A(_12246_), .B(_12247_), .Y(_00302_));
NAND_g _18138_ (.A(_11566_), .B(_12204_), .Y(_12248_));
NAND_g _18139_ (.A(cpuregs_27[21]), .B(_12205_), .Y(_12249_));
NAND_g _18140_ (.A(_12248_), .B(_12249_), .Y(_00303_));
NAND_g _18141_ (.A(_11579_), .B(_12204_), .Y(_12250_));
NAND_g _18142_ (.A(cpuregs_27[22]), .B(_12205_), .Y(_12251_));
NAND_g _18143_ (.A(_12250_), .B(_12251_), .Y(_00304_));
NAND_g _18144_ (.A(_11592_), .B(_12204_), .Y(_12252_));
NAND_g _18145_ (.A(cpuregs_27[23]), .B(_12205_), .Y(_12253_));
NAND_g _18146_ (.A(_12252_), .B(_12253_), .Y(_00305_));
NAND_g _18147_ (.A(_11605_), .B(_12204_), .Y(_12254_));
NAND_g _18148_ (.A(cpuregs_27[24]), .B(_12205_), .Y(_12255_));
NAND_g _18149_ (.A(_12254_), .B(_12255_), .Y(_00306_));
NAND_g _18150_ (.A(_11618_), .B(_12204_), .Y(_12256_));
NAND_g _18151_ (.A(cpuregs_27[25]), .B(_12205_), .Y(_12257_));
NAND_g _18152_ (.A(_12256_), .B(_12257_), .Y(_00307_));
NAND_g _18153_ (.A(_11631_), .B(_12204_), .Y(_12258_));
NAND_g _18154_ (.A(cpuregs_27[26]), .B(_12205_), .Y(_12259_));
NAND_g _18155_ (.A(_12258_), .B(_12259_), .Y(_00308_));
NAND_g _18156_ (.A(_11644_), .B(_12204_), .Y(_12260_));
NAND_g _18157_ (.A(cpuregs_27[27]), .B(_12205_), .Y(_12261_));
NAND_g _18158_ (.A(_12260_), .B(_12261_), .Y(_00309_));
NAND_g _18159_ (.A(_11657_), .B(_12204_), .Y(_12262_));
NAND_g _18160_ (.A(cpuregs_27[28]), .B(_12205_), .Y(_12263_));
NAND_g _18161_ (.A(_12262_), .B(_12263_), .Y(_00310_));
NAND_g _18162_ (.A(_11670_), .B(_12204_), .Y(_12264_));
NAND_g _18163_ (.A(cpuregs_27[29]), .B(_12205_), .Y(_12265_));
NAND_g _18164_ (.A(_12264_), .B(_12265_), .Y(_00311_));
NAND_g _18165_ (.A(_11683_), .B(_12204_), .Y(_12266_));
NAND_g _18166_ (.A(cpuregs_27[30]), .B(_12205_), .Y(_12267_));
NAND_g _18167_ (.A(_12266_), .B(_12267_), .Y(_00312_));
NAND_g _18168_ (.A(_11695_), .B(_12204_), .Y(_12268_));
NAND_g _18169_ (.A(cpuregs_27[31]), .B(_12205_), .Y(_12269_));
NAND_g _18170_ (.A(_12268_), .B(_12269_), .Y(_00313_));
NAND_g _18171_ (.A(instr_jalr), .B(_11919_), .Y(_12270_));
NAND_g _18172_ (.A(mem_rdata[14]), .B(_11910_), .Y(_12271_));
NAND_g _18173_ (.A(mem_rdata_q[14]), .B(_11911_), .Y(_12272_));
NAND_g _18174_ (.A(_12271_), .B(_12272_), .Y(_00786_));
NOR_g _18175_ (.A(_11919_), .B(_00786_), .Y(_12273_));
NAND_g _18176_ (.A(mem_rdata[0]), .B(_11910_), .Y(_12274_));
NAND_g _18177_ (.A(mem_rdata_q[0]), .B(_11911_), .Y(_12275_));
NAND_g _18178_ (.A(_12274_), .B(_12275_), .Y(_00872_));
NAND_g _18179_ (.A(mem_rdata[1]), .B(_11910_), .Y(_12276_));
NAND_g _18180_ (.A(mem_rdata_q[1]), .B(_11911_), .Y(_12277_));
NAND_g _18181_ (.A(_12276_), .B(_12277_), .Y(_00873_));
AND_g _18182_ (.A(_00872_), .B(_00873_), .Y(_12278_));
NAND_g _18183_ (.A(mem_rdata[2]), .B(_11910_), .Y(_12279_));
NAND_g _18184_ (.A(mem_rdata_q[2]), .B(_11911_), .Y(_12280_));
NAND_g _18185_ (.A(_12279_), .B(_12280_), .Y(_00874_));
AND_g _18186_ (.A(_12278_), .B(_00874_), .Y(_12281_));
NAND_g _18187_ (.A(mem_rdata[3]), .B(_11910_), .Y(_12282_));
NAND_g _18188_ (.A(mem_rdata_q[3]), .B(_11911_), .Y(_12283_));
NAND_g _18189_ (.A(_12282_), .B(_12283_), .Y(_00875_));
NOT_g _18190_ (.A(_00875_), .Y(_12284_));
AND_g _18191_ (.A(_12281_), .B(_12284_), .Y(_12285_));
NAND_g _18192_ (.A(mem_rdata[4]), .B(_11910_), .Y(_12286_));
NAND_g _18193_ (.A(mem_rdata_q[4]), .B(_11911_), .Y(_12287_));
AND_g _18194_ (.A(_12286_), .B(_12287_), .Y(_12288_));
NOT_g _18195_ (.A(_12288_), .Y(_00876_));
NAND_g _18196_ (.A(mem_rdata[5]), .B(_11910_), .Y(_12289_));
NAND_g _18197_ (.A(mem_rdata_q[5]), .B(_11911_), .Y(_12290_));
NAND_g _18198_ (.A(_12289_), .B(_12290_), .Y(_00877_));
NOT_g _18199_ (.A(_00877_), .Y(_12291_));
AND_g _18200_ (.A(_12288_), .B(_00877_), .Y(_12292_));
NAND_g _18201_ (.A(mem_rdata[6]), .B(_11910_), .Y(_12293_));
NAND_g _18202_ (.A(mem_rdata_q[6]), .B(_11911_), .Y(_12294_));
NAND_g _18203_ (.A(_12293_), .B(_12294_), .Y(_00878_));
NOT_g _18204_ (.A(_00878_), .Y(_12295_));
AND_g _18205_ (.A(_12292_), .B(_00878_), .Y(_12296_));
NAND_g _18206_ (.A(mem_rdata[13]), .B(_11910_), .Y(_12297_));
NAND_g _18207_ (.A(mem_rdata_q[13]), .B(_11911_), .Y(_12298_));
NAND_g _18208_ (.A(_12297_), .B(_12298_), .Y(_00785_));
NAND_g _18209_ (.A(mem_rdata[12]), .B(_11910_), .Y(_12299_));
NAND_g _18210_ (.A(mem_rdata_q[12]), .B(_11911_), .Y(_12300_));
NAND_g _18211_ (.A(_12299_), .B(_12300_), .Y(_00784_));
NOR_g _18212_ (.A(_00785_), .B(_00784_), .Y(_12301_));
AND_g _18213_ (.A(_12296_), .B(_12301_), .Y(_12302_));
AND_g _18214_ (.A(_12285_), .B(_12302_), .Y(_12303_));
NAND_g _18215_ (.A(_12273_), .B(_12303_), .Y(_12304_));
NAND_g _18216_ (.A(_12270_), .B(_12304_), .Y(_00314_));
NAND_g _18217_ (.A(instr_auipc), .B(_11919_), .Y(_12305_));
NOR_g _18218_ (.A(_12288_), .B(_00878_), .Y(_12306_));
AND_g _18219_ (.A(_12291_), .B(_12306_), .Y(_12307_));
AND_g _18220_ (.A(_11918_), .B(_12285_), .Y(_12308_));
NAND_g _18221_ (.A(_12307_), .B(_12308_), .Y(_12309_));
NAND_g _18222_ (.A(_12305_), .B(_12309_), .Y(_00315_));
AND_g _18223_ (.A(_12281_), .B(_00875_), .Y(_12310_));
AND_g _18224_ (.A(_12296_), .B(_12310_), .Y(_12311_));
NAND_g _18225_ (.A(instr_jal), .B(_11919_), .Y(_12312_));
NAND_g _18226_ (.A(_11918_), .B(_12311_), .Y(_12313_));
NAND_g _18227_ (.A(_12312_), .B(_12313_), .Y(_00316_));
AND_g _18228_ (.A(decoder_trigger), .B(_11211_), .Y(_12314_));
NAND_g _18229_ (.A(decoder_trigger), .B(_11211_), .Y(_12315_));
AND_g _18230_ (.A(resetn), .B(_12315_), .Y(_12316_));
NAND_g _18231_ (.A(instr_beq), .B(_12316_), .Y(_12317_));
NOR_g _18232_ (.A(mem_rdata_q[12]), .B(mem_rdata_q[13]), .Y(_12318_));
AND_g _18233_ (.A(_11079_), .B(_12318_), .Y(_12319_));
AND_g _18234_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(resetn), .Y(_12320_));
AND_g _18235_ (.A(_12314_), .B(_12320_), .Y(_12321_));
NAND_g _18236_ (.A(_12319_), .B(_12321_), .Y(_12322_));
NAND_g _18237_ (.A(_12317_), .B(_12322_), .Y(_00317_));
AND_g _18238_ (.A(mem_rdata_q[12]), .B(_11078_), .Y(_12323_));
NAND_g _18239_ (.A(mem_rdata_q[12]), .B(_11078_), .Y(_12324_));
AND_g _18240_ (.A(_11079_), .B(_12323_), .Y(_12325_));
NAND_g _18241_ (.A(_12321_), .B(_12325_), .Y(_12326_));
NAND_g _18242_ (.A(instr_bne), .B(_12316_), .Y(_12327_));
NAND_g _18243_ (.A(_12326_), .B(_12327_), .Y(_00318_));
AND_g _18244_ (.A(mem_rdata_q[14]), .B(_12318_), .Y(_12328_));
NAND_g _18245_ (.A(_12321_), .B(_12328_), .Y(_12329_));
NAND_g _18246_ (.A(instr_blt), .B(_12316_), .Y(_12330_));
NAND_g _18247_ (.A(_12329_), .B(_12330_), .Y(_00319_));
AND_g _18248_ (.A(mem_rdata_q[14]), .B(_12323_), .Y(_12331_));
NAND_g _18249_ (.A(_12321_), .B(_12331_), .Y(_12332_));
NAND_g _18250_ (.A(instr_bge), .B(_12316_), .Y(_12333_));
NAND_g _18251_ (.A(_12332_), .B(_12333_), .Y(_00320_));
AND_g _18252_ (.A(_11077_), .B(mem_rdata_q[13]), .Y(_12334_));
AND_g _18253_ (.A(mem_rdata_q[14]), .B(_12334_), .Y(_12335_));
NAND_g _18254_ (.A(_12321_), .B(_12335_), .Y(_12336_));
NAND_g _18255_ (.A(instr_bltu), .B(_12316_), .Y(_12337_));
NAND_g _18256_ (.A(_12336_), .B(_12337_), .Y(_00321_));
AND_g _18257_ (.A(mem_rdata_q[12]), .B(mem_rdata_q[13]), .Y(_12338_));
AND_g _18258_ (.A(mem_rdata_q[14]), .B(_12338_), .Y(_12339_));
NAND_g _18259_ (.A(_12321_), .B(_12339_), .Y(_12340_));
NAND_g _18260_ (.A(instr_bgeu), .B(_12316_), .Y(_12341_));
NAND_g _18261_ (.A(_12340_), .B(_12341_), .Y(_00322_));
NAND_g _18262_ (.A(is_sll_srl_sra), .B(_12315_), .Y(_12342_));
NOR_g _18263_ (.A(mem_rdata_q[25]), .B(mem_rdata_q[26]), .Y(_12343_));
NOR_g _18264_ (.A(mem_rdata_q[27]), .B(mem_rdata_q[28]), .Y(_12344_));
AND_g _18265_ (.A(_11083_), .B(_12344_), .Y(_12345_));
AND_g _18266_ (.A(_12343_), .B(_12345_), .Y(_12346_));
NOR_g _18267_ (.A(mem_rdata_q[29]), .B(mem_rdata_q[30]), .Y(_12347_));
AND_g _18268_ (.A(_12346_), .B(_12347_), .Y(_12348_));
NAND_g _18269_ (.A(_12323_), .B(_12348_), .Y(_12349_));
AND_g _18270_ (.A(_11082_), .B(mem_rdata_q[30]), .Y(_12350_));
AND_g _18271_ (.A(_12346_), .B(_12350_), .Y(_12351_));
AND_g _18272_ (.A(_12331_), .B(_12351_), .Y(_12352_));
NOT_g _18273_ (.A(_12352_), .Y(_12353_));
NAND_g _18274_ (.A(_12349_), .B(_12353_), .Y(_12354_));
AND_g _18275_ (.A(is_alu_reg_reg), .B(_12314_), .Y(_12355_));
NAND_g _18276_ (.A(_12354_), .B(_12355_), .Y(_12356_));
NAND_g _18277_ (.A(_12342_), .B(_12356_), .Y(_00323_));
NAND_g _18278_ (.A(instr_lb), .B(_12315_), .Y(_12357_));
AND_g _18279_ (.A(is_lb_lh_lw_lbu_lhu), .B(_12314_), .Y(_12358_));
NAND_g _18280_ (.A(_12319_), .B(_12358_), .Y(_12359_));
NAND_g _18281_ (.A(_12357_), .B(_12359_), .Y(_00324_));
NAND_g _18282_ (.A(instr_lh), .B(_12315_), .Y(_12360_));
NAND_g _18283_ (.A(_12325_), .B(_12358_), .Y(_12361_));
NAND_g _18284_ (.A(_12360_), .B(_12361_), .Y(_00325_));
NAND_g _18285_ (.A(instr_lw), .B(_12315_), .Y(_12362_));
AND_g _18286_ (.A(_11079_), .B(_12334_), .Y(_12363_));
NAND_g _18287_ (.A(_12358_), .B(_12363_), .Y(_12364_));
NAND_g _18288_ (.A(_12362_), .B(_12364_), .Y(_00326_));
NAND_g _18289_ (.A(instr_lbu), .B(_12315_), .Y(_12365_));
NAND_g _18290_ (.A(_12328_), .B(_12358_), .Y(_12366_));
NAND_g _18291_ (.A(_12365_), .B(_12366_), .Y(_00327_));
NAND_g _18292_ (.A(instr_lhu), .B(_12315_), .Y(_12367_));
NAND_g _18293_ (.A(_12331_), .B(_12358_), .Y(_12368_));
NAND_g _18294_ (.A(_12367_), .B(_12368_), .Y(_00328_));
NAND_g _18295_ (.A(instr_sb), .B(_12315_), .Y(_12369_));
AND_g _18296_ (.A(is_sb_sh_sw), .B(_12314_), .Y(_12370_));
NAND_g _18297_ (.A(_12319_), .B(_12370_), .Y(_12371_));
NAND_g _18298_ (.A(_12369_), .B(_12371_), .Y(_00329_));
NAND_g _18299_ (.A(instr_sh), .B(_12315_), .Y(_12372_));
NAND_g _18300_ (.A(_12325_), .B(_12370_), .Y(_12373_));
NAND_g _18301_ (.A(_12372_), .B(_12373_), .Y(_00330_));
NAND_g _18302_ (.A(instr_addi), .B(_12316_), .Y(_12374_));
AND_g _18303_ (.A(is_alu_reg_imm), .B(_12314_), .Y(_12375_));
AND_g _18304_ (.A(resetn), .B(_12375_), .Y(_12376_));
NAND_g _18305_ (.A(_12319_), .B(_12376_), .Y(_12377_));
NAND_g _18306_ (.A(_12374_), .B(_12377_), .Y(_00331_));
NAND_g _18307_ (.A(instr_slti), .B(_12316_), .Y(_12378_));
NAND_g _18308_ (.A(_12363_), .B(_12376_), .Y(_12379_));
NAND_g _18309_ (.A(_12378_), .B(_12379_), .Y(_00332_));
AND_g _18310_ (.A(_11079_), .B(_12338_), .Y(_12380_));
NAND_g _18311_ (.A(_12376_), .B(_12380_), .Y(_12381_));
NAND_g _18312_ (.A(instr_sltiu), .B(_12316_), .Y(_12382_));
NAND_g _18313_ (.A(_12381_), .B(_12382_), .Y(_00333_));
NAND_g _18314_ (.A(instr_xori), .B(_12316_), .Y(_12383_));
NAND_g _18315_ (.A(_12328_), .B(_12376_), .Y(_12384_));
NAND_g _18316_ (.A(_12383_), .B(_12384_), .Y(_00334_));
NAND_g _18317_ (.A(instr_ori), .B(_12316_), .Y(_12385_));
NAND_g _18318_ (.A(_12335_), .B(_12376_), .Y(_12386_));
NAND_g _18319_ (.A(_12385_), .B(_12386_), .Y(_00335_));
NAND_g _18320_ (.A(instr_andi), .B(_12316_), .Y(_12387_));
NAND_g _18321_ (.A(_12339_), .B(_12376_), .Y(_12388_));
NAND_g _18322_ (.A(_12387_), .B(_12388_), .Y(_00336_));
NAND_g _18323_ (.A(instr_sw), .B(_12315_), .Y(_12389_));
NAND_g _18324_ (.A(_12363_), .B(_12370_), .Y(_12390_));
NAND_g _18325_ (.A(_12389_), .B(_12390_), .Y(_00337_));
NAND_g _18326_ (.A(instr_slli), .B(_12315_), .Y(_12391_));
AND_g _18327_ (.A(_12325_), .B(_12348_), .Y(_12392_));
NAND_g _18328_ (.A(_12375_), .B(_12392_), .Y(_12393_));
NAND_g _18329_ (.A(_12391_), .B(_12393_), .Y(_00338_));
NAND_g _18330_ (.A(instr_srli), .B(_12315_), .Y(_12394_));
AND_g _18331_ (.A(_12331_), .B(_12375_), .Y(_12395_));
NAND_g _18332_ (.A(_12348_), .B(_12395_), .Y(_12396_));
NAND_g _18333_ (.A(_12394_), .B(_12396_), .Y(_00339_));
NAND_g _18334_ (.A(instr_add), .B(_12316_), .Y(_12397_));
AND_g _18335_ (.A(resetn), .B(_12355_), .Y(_12398_));
AND_g _18336_ (.A(_12319_), .B(_12398_), .Y(_12399_));
NAND_g _18337_ (.A(_12348_), .B(_12399_), .Y(_12400_));
NAND_g _18338_ (.A(_12397_), .B(_12400_), .Y(_00340_));
NAND_g _18339_ (.A(instr_sub), .B(_12316_), .Y(_12401_));
NAND_g _18340_ (.A(_12351_), .B(_12399_), .Y(_12402_));
NAND_g _18341_ (.A(_12401_), .B(_12402_), .Y(_00341_));
NAND_g _18342_ (.A(instr_sll), .B(_12316_), .Y(_12403_));
AND_g _18343_ (.A(_12348_), .B(_12398_), .Y(_12404_));
NAND_g _18344_ (.A(_12325_), .B(_12404_), .Y(_12405_));
NAND_g _18345_ (.A(_12403_), .B(_12405_), .Y(_00342_));
NAND_g _18346_ (.A(_12363_), .B(_12404_), .Y(_12406_));
NAND_g _18347_ (.A(instr_slt), .B(_12316_), .Y(_12407_));
NAND_g _18348_ (.A(_12406_), .B(_12407_), .Y(_00343_));
NAND_g _18349_ (.A(instr_sltu), .B(_12316_), .Y(_12408_));
NAND_g _18350_ (.A(_12380_), .B(_12404_), .Y(_12409_));
NAND_g _18351_ (.A(_12408_), .B(_12409_), .Y(_00344_));
NAND_g _18352_ (.A(_12328_), .B(_12404_), .Y(_12410_));
NAND_g _18353_ (.A(instr_xor), .B(_12316_), .Y(_12411_));
NAND_g _18354_ (.A(_12410_), .B(_12411_), .Y(_00345_));
NAND_g _18355_ (.A(instr_srl), .B(_12316_), .Y(_12412_));
NAND_g _18356_ (.A(_12331_), .B(_12404_), .Y(_12413_));
NAND_g _18357_ (.A(_12412_), .B(_12413_), .Y(_00346_));
NAND_g _18358_ (.A(instr_sra), .B(_12316_), .Y(_12414_));
NAND_g _18359_ (.A(_12352_), .B(_12398_), .Y(_12415_));
NAND_g _18360_ (.A(_12414_), .B(_12415_), .Y(_00347_));
NAND_g _18361_ (.A(instr_or), .B(_12316_), .Y(_12416_));
NAND_g _18362_ (.A(_12335_), .B(_12404_), .Y(_12417_));
NAND_g _18363_ (.A(_12416_), .B(_12417_), .Y(_00348_));
NAND_g _18364_ (.A(instr_and), .B(_12316_), .Y(_12418_));
NAND_g _18365_ (.A(_12339_), .B(_12404_), .Y(_12419_));
NAND_g _18366_ (.A(_12418_), .B(_12419_), .Y(_00349_));
NAND_g _18367_ (.A(instr_srai), .B(_12315_), .Y(_12420_));
NAND_g _18368_ (.A(_12352_), .B(_12375_), .Y(_12421_));
NAND_g _18369_ (.A(_12420_), .B(_12421_), .Y(_00350_));
NAND_g _18370_ (.A(instr_rdcycle), .B(_12315_), .Y(_12422_));
NOR_g _18371_ (.A(mem_rdata_q[24]), .B(_12315_), .Y(_12423_));
NAND_g _18372_ (.A(_12343_), .B(_12423_), .Y(_12424_));
NOR_g _18373_ (.A(mem_rdata_q[27]), .B(_12424_), .Y(_12425_));
NOR_g _18374_ (.A(mem_rdata_q[15]), .B(mem_rdata_q[16]), .Y(_12426_));
AND_g _18375_ (.A(mem_rdata_q[31]), .B(mem_rdata_q[0]), .Y(_12427_));
AND_g _18376_ (.A(mem_rdata_q[1]), .B(_11085_), .Y(_12428_));
AND_g _18377_ (.A(_12427_), .B(_12428_), .Y(_12429_));
AND_g _18378_ (.A(_11086_), .B(mem_rdata_q[4]), .Y(_12430_));
AND_g _18379_ (.A(mem_rdata_q[5]), .B(mem_rdata_q[6]), .Y(_12431_));
AND_g _18380_ (.A(_12430_), .B(_12431_), .Y(_12432_));
NOR_g _18381_ (.A(mem_rdata_q[22]), .B(mem_rdata_q[23]), .Y(_12433_));
AND_g _18382_ (.A(_12429_), .B(_12432_), .Y(_12434_));
NOR_g _18383_ (.A(mem_rdata_q[18]), .B(mem_rdata_q[19]), .Y(_12435_));
NOR_g _18384_ (.A(mem_rdata_q[17]), .B(mem_rdata_q[28]), .Y(_12436_));
AND_g _18385_ (.A(_12435_), .B(_12436_), .Y(_12437_));
AND_g _18386_ (.A(_12350_), .B(_12426_), .Y(_12438_));
AND_g _18387_ (.A(_12437_), .B(_12438_), .Y(_12439_));
AND_g _18388_ (.A(_12363_), .B(_12439_), .Y(_12440_));
AND_g _18389_ (.A(_12434_), .B(_12440_), .Y(_12441_));
NAND_g _18390_ (.A(_12433_), .B(_12441_), .Y(_12442_));
NOR_g _18391_ (.A(mem_rdata_q[21]), .B(_12442_), .Y(_12443_));
NAND_g _18392_ (.A(_12425_), .B(_12443_), .Y(_12444_));
NAND_g _18393_ (.A(_12422_), .B(_12444_), .Y(_00351_));
NAND_g _18394_ (.A(instr_rdcycleh), .B(_12315_), .Y(_12445_));
NOR_g _18395_ (.A(_11081_), .B(_12424_), .Y(_12446_));
NAND_g _18396_ (.A(_12443_), .B(_12446_), .Y(_12447_));
NAND_g _18397_ (.A(_12445_), .B(_12447_), .Y(_00352_));
NAND_g _18398_ (.A(instr_rdinstr), .B(_12315_), .Y(_12448_));
NAND_g _18399_ (.A(_11080_), .B(mem_rdata_q[21]), .Y(_12449_));
NOR_g _18400_ (.A(_12442_), .B(_12449_), .Y(_12450_));
NAND_g _18401_ (.A(_12425_), .B(_12450_), .Y(_12451_));
NAND_g _18402_ (.A(_12448_), .B(_12451_), .Y(_00353_));
NAND_g _18403_ (.A(instr_rdinstrh), .B(_12315_), .Y(_12452_));
NAND_g _18404_ (.A(_12446_), .B(_12450_), .Y(_12453_));
NAND_g _18405_ (.A(_12452_), .B(_12453_), .Y(_00354_));
NAND_g _18406_ (.A(mem_rdata[7]), .B(_11910_), .Y(_12454_));
NAND_g _18407_ (.A(mem_rdata_q[7]), .B(_11911_), .Y(_12455_));
NAND_g _18408_ (.A(_12454_), .B(_12455_), .Y(_00779_));
NAND_g _18409_ (.A(_11918_), .B(_00779_), .Y(_12456_));
NAND_g _18410_ (.A(decoded_rd[0]), .B(_11919_), .Y(_12457_));
NAND_g _18411_ (.A(_12456_), .B(_12457_), .Y(_00355_));
NAND_g _18412_ (.A(mem_rdata[8]), .B(_11910_), .Y(_12458_));
NAND_g _18413_ (.A(mem_rdata_q[8]), .B(_11911_), .Y(_12459_));
NAND_g _18414_ (.A(_12458_), .B(_12459_), .Y(_00780_));
NAND_g _18415_ (.A(_11918_), .B(_00780_), .Y(_12460_));
NAND_g _18416_ (.A(decoded_rd[1]), .B(_11919_), .Y(_12461_));
NAND_g _18417_ (.A(_12460_), .B(_12461_), .Y(_00356_));
NAND_g _18418_ (.A(mem_rdata[9]), .B(_11910_), .Y(_12462_));
NAND_g _18419_ (.A(mem_rdata_q[9]), .B(_11911_), .Y(_12463_));
NAND_g _18420_ (.A(_12462_), .B(_12463_), .Y(_00781_));
NAND_g _18421_ (.A(_11918_), .B(_00781_), .Y(_12464_));
NAND_g _18422_ (.A(decoded_rd[2]), .B(_11919_), .Y(_12465_));
NAND_g _18423_ (.A(_12464_), .B(_12465_), .Y(_00357_));
NAND_g _18424_ (.A(mem_rdata[10]), .B(_11910_), .Y(_12466_));
NAND_g _18425_ (.A(mem_rdata_q[10]), .B(_11911_), .Y(_12467_));
NAND_g _18426_ (.A(_12466_), .B(_12467_), .Y(_00782_));
NAND_g _18427_ (.A(_11918_), .B(_00782_), .Y(_12468_));
NAND_g _18428_ (.A(decoded_rd[3]), .B(_11919_), .Y(_12469_));
NAND_g _18429_ (.A(_12468_), .B(_12469_), .Y(_00358_));
NAND_g _18430_ (.A(mem_rdata[11]), .B(_11910_), .Y(_12470_));
NAND_g _18431_ (.A(mem_rdata_q[11]), .B(_11911_), .Y(_12471_));
NAND_g _18432_ (.A(_12470_), .B(_12471_), .Y(_00783_));
NAND_g _18433_ (.A(_11918_), .B(_00783_), .Y(_12472_));
NAND_g _18434_ (.A(decoded_rd[4]), .B(_11919_), .Y(_12473_));
NAND_g _18435_ (.A(_12472_), .B(_12473_), .Y(_00359_));
NAND_g _18436_ (.A(mem_rdata[20]), .B(_11910_), .Y(_12474_));
NAND_g _18437_ (.A(mem_rdata_q[20]), .B(_11911_), .Y(_12475_));
NAND_g _18438_ (.A(_12474_), .B(_12475_), .Y(_00792_));
NAND_g _18439_ (.A(_11918_), .B(_00792_), .Y(_12476_));
NAND_g _18440_ (.A(decoded_imm_j[11]), .B(_11919_), .Y(_12477_));
NAND_g _18441_ (.A(_12476_), .B(_12477_), .Y(_00360_));
NAND_g _18442_ (.A(mem_rdata[23]), .B(_11910_), .Y(_12478_));
NAND_g _18443_ (.A(mem_rdata_q[23]), .B(_11911_), .Y(_12479_));
NAND_g _18444_ (.A(_12478_), .B(_12479_), .Y(_00795_));
NAND_g _18445_ (.A(_11918_), .B(_00795_), .Y(_12480_));
NAND_g _18446_ (.A(decoded_imm_j[3]), .B(_11919_), .Y(_12481_));
NAND_g _18447_ (.A(_12480_), .B(_12481_), .Y(_00361_));
NAND_g _18448_ (.A(mem_rdata_q[7]), .B(_12370_), .Y(_12482_));
NOR_g _18449_ (.A(instr_jalr), .B(is_lb_lh_lw_lbu_lhu), .Y(_12483_));
NAND_g _18450_ (.A(_10981_), .B(_12483_), .Y(_12484_));
NOT_g _18451_ (.A(_12484_), .Y(_12485_));
AND_g _18452_ (.A(mem_rdata_q[20]), .B(_12314_), .Y(_12486_));
NAND_g _18453_ (.A(_12484_), .B(_12486_), .Y(_12487_));
NAND_g _18454_ (.A(decoded_imm[0]), .B(_12315_), .Y(_12488_));
AND_g _18455_ (.A(_12482_), .B(_12487_), .Y(_12489_));
NAND_g _18456_ (.A(_12488_), .B(_12489_), .Y(_00362_));
NAND_g _18457_ (.A(mem_rdata[21]), .B(_11910_), .Y(_12490_));
NAND_g _18458_ (.A(mem_rdata_q[21]), .B(_11911_), .Y(_12491_));
NAND_g _18459_ (.A(_12490_), .B(_12491_), .Y(_00793_));
NAND_g _18460_ (.A(_11918_), .B(_00793_), .Y(_12492_));
NAND_g _18461_ (.A(decoded_imm_j[1]), .B(_11919_), .Y(_12493_));
NAND_g _18462_ (.A(_12492_), .B(_12493_), .Y(_00363_));
NAND_g _18463_ (.A(mem_rdata[22]), .B(_11910_), .Y(_12494_));
NAND_g _18464_ (.A(mem_rdata_q[22]), .B(_11911_), .Y(_12495_));
NAND_g _18465_ (.A(_12494_), .B(_12495_), .Y(_00794_));
NAND_g _18466_ (.A(_11918_), .B(_00794_), .Y(_12496_));
NAND_g _18467_ (.A(decoded_imm_j[2]), .B(_11919_), .Y(_12497_));
NAND_g _18468_ (.A(_12496_), .B(_12497_), .Y(_00364_));
NAND_g _18469_ (.A(is_lb_lh_lw_lbu_lhu), .B(_11919_), .Y(_12498_));
NOR_g _18470_ (.A(_00877_), .B(_00878_), .Y(_12499_));
NOR_g _18471_ (.A(_00874_), .B(_00875_), .Y(_12500_));
AND_g _18472_ (.A(_12278_), .B(_12500_), .Y(_12501_));
AND_g _18473_ (.A(_11918_), .B(_12501_), .Y(_12502_));
AND_g _18474_ (.A(_12499_), .B(_12502_), .Y(_12503_));
NAND_g _18475_ (.A(_12288_), .B(_12503_), .Y(_12504_));
NAND_g _18476_ (.A(_12498_), .B(_12504_), .Y(_00365_));
NAND_g _18477_ (.A(is_slli_srli_srai), .B(_12315_), .Y(_12505_));
NAND_g _18478_ (.A(_12354_), .B(_12375_), .Y(_12506_));
NAND_g _18479_ (.A(_12505_), .B(_12506_), .Y(_00366_));
NAND_g _18480_ (.A(is_alu_reg_imm), .B(_12324_), .Y(_12507_));
NAND_g _18481_ (.A(_10978_), .B(_12315_), .Y(_12508_));
NOR_g _18482_ (.A(instr_jalr), .B(_12315_), .Y(_12509_));
NAND_g _18483_ (.A(_12507_), .B(_12509_), .Y(_12510_));
AND_g _18484_ (.A(_12508_), .B(_12510_), .Y(_00367_));
NAND_g _18485_ (.A(instr_lui), .B(_11919_), .Y(_12511_));
AND_g _18486_ (.A(_00877_), .B(_12306_), .Y(_12512_));
NAND_g _18487_ (.A(_12308_), .B(_12512_), .Y(_12513_));
NAND_g _18488_ (.A(_12511_), .B(_12513_), .Y(_00368_));
NAND_g _18489_ (.A(is_sb_sh_sw), .B(_11919_), .Y(_12514_));
AND_g _18490_ (.A(_12292_), .B(_12295_), .Y(_12515_));
NAND_g _18491_ (.A(_12502_), .B(_12515_), .Y(_12516_));
NAND_g _18492_ (.A(_12514_), .B(_12516_), .Y(_00369_));
NAND_g _18493_ (.A(_11919_), .B(_12320_), .Y(_12517_));
NAND_g _18494_ (.A(_12296_), .B(_12502_), .Y(_12518_));
NAND_g _18495_ (.A(_12517_), .B(_12518_), .Y(_00370_));
NOR_g _18496_ (.A(instr_auipc), .B(instr_lui), .Y(_12519_));
NAND_g _18497_ (.A(_10961_), .B(_10979_), .Y(_12520_));
AND_g _18498_ (.A(_10962_), .B(_12519_), .Y(_12521_));
NOT_g _18499_ (.A(_12521_), .Y(_00006_));
NOR_g _18500_ (.A(instr_sub), .B(instr_add), .Y(_12522_));
NOR_g _18501_ (.A(instr_addi), .B(instr_jalr), .Y(_12523_));
AND_g _18502_ (.A(_12522_), .B(_12523_), .Y(_12524_));
NAND_g _18503_ (.A(_12521_), .B(_12524_), .Y(_12525_));
AND_g _18504_ (.A(_12315_), .B(_12525_), .Y(_00371_));
NAND_g _18505_ (.A(is_alu_reg_imm), .B(_11919_), .Y(_12526_));
NAND_g _18506_ (.A(_12307_), .B(_12502_), .Y(_12527_));
NAND_g _18507_ (.A(_12526_), .B(_12527_), .Y(_00372_));
NAND_g _18508_ (.A(_12502_), .B(_12512_), .Y(_12528_));
NAND_g _18509_ (.A(is_alu_reg_reg), .B(_11919_), .Y(_12529_));
NAND_g _18510_ (.A(_12528_), .B(_12529_), .Y(_00373_));
NOR_g _18511_ (.A(instr_sltiu), .B(instr_slti), .Y(_12530_));
NOR_g _18512_ (.A(instr_sltu), .B(instr_slt), .Y(_12531_));
AND_g _18513_ (.A(_12530_), .B(_12531_), .Y(_12532_));
NAND_g _18514_ (.A(_10902_), .B(_12532_), .Y(_12533_));
AND_g _18515_ (.A(_12316_), .B(_12533_), .Y(_00374_));
AND_g _18516_ (.A(resetn), .B(_11916_), .Y(_12534_));
NAND_g _18517_ (.A(resetn), .B(_11916_), .Y(_12535_));
NAND_g _18518_ (.A(_10962_), .B(decoder_trigger), .Y(_12536_));
AND_g _18519_ (.A(_10962_), .B(launch_next_insn), .Y(_12537_));
NOR_g _18520_ (.A(mem_do_prefetch), .B(_12537_), .Y(_12538_));
NOR_g _18521_ (.A(_12535_), .B(_12538_), .Y(_12539_));
AND_g _18522_ (.A(instr_jalr), .B(_12537_), .Y(_12540_));
NAND_g _18523_ (.A(resetn), .B(_12540_), .Y(_12541_));
AND_g _18524_ (.A(_12539_), .B(_12541_), .Y(_00375_));
AND_g _18525_ (.A(latched_branch), .B(latched_store), .Y(_12542_));
NAND_g _18526_ (.A(latched_branch), .B(latched_store), .Y(_12543_));
NAND_g _18527_ (.A(_11306_), .B(_12542_), .Y(_12544_));
NAND_g _18528_ (.A(reg_next_pc[1]), .B(_12543_), .Y(_12545_));
NAND_g _18529_ (.A(_12544_), .B(_12545_), .Y(_12546_));
AND_g _18530_ (.A(_11275_), .B(_12546_), .Y(_12547_));
NOT_g _18531_ (.A(_12547_), .Y(_12548_));
AND_g _18532_ (.A(resetn), .B(_11263_), .Y(_12549_));
NAND_g _18533_ (.A(reg_pc[1]), .B(_12549_), .Y(_12550_));
NAND_g _18534_ (.A(_12548_), .B(_12550_), .Y(_00376_));
NAND_g _18535_ (.A(reg_next_pc[2]), .B(_12543_), .Y(_12551_));
NAND_g _18536_ (.A(_11315_), .B(_12542_), .Y(_12552_));
NAND_g _18537_ (.A(_12551_), .B(_12552_), .Y(_12553_));
AND_g _18538_ (.A(_11275_), .B(_12553_), .Y(_12554_));
NAND_g _18539_ (.A(_11275_), .B(_12553_), .Y(_12555_));
NAND_g _18540_ (.A(reg_pc[2]), .B(_12549_), .Y(_12556_));
NAND_g _18541_ (.A(_12555_), .B(_12556_), .Y(_00377_));
NAND_g _18542_ (.A(reg_next_pc[3]), .B(_12543_), .Y(_12557_));
NAND_g _18543_ (.A(_11324_), .B(_12542_), .Y(_12558_));
NAND_g _18544_ (.A(_12557_), .B(_12558_), .Y(_12559_));
AND_g _18545_ (.A(_11275_), .B(_12559_), .Y(_12560_));
NAND_g _18546_ (.A(_11275_), .B(_12559_), .Y(_12561_));
NAND_g _18547_ (.A(reg_pc[3]), .B(_12549_), .Y(_12562_));
NAND_g _18548_ (.A(_12561_), .B(_12562_), .Y(_00378_));
NAND_g _18549_ (.A(reg_next_pc[4]), .B(_12543_), .Y(_12563_));
NAND_g _18550_ (.A(_11337_), .B(_12542_), .Y(_12564_));
NAND_g _18551_ (.A(_12563_), .B(_12564_), .Y(_12565_));
NAND_g _18552_ (.A(_11275_), .B(_12565_), .Y(_12566_));
NOT_g _18553_ (.A(_12566_), .Y(_12567_));
NAND_g _18554_ (.A(reg_pc[4]), .B(_12549_), .Y(_12568_));
NAND_g _18555_ (.A(_12566_), .B(_12568_), .Y(_00379_));
NAND_g _18556_ (.A(reg_next_pc[5]), .B(_12543_), .Y(_12569_));
NAND_g _18557_ (.A(_11350_), .B(_12542_), .Y(_12570_));
NAND_g _18558_ (.A(_12569_), .B(_12570_), .Y(_12571_));
AND_g _18559_ (.A(_11275_), .B(_12571_), .Y(_12572_));
NOT_g _18560_ (.A(_12572_), .Y(_12573_));
NAND_g _18561_ (.A(reg_pc[5]), .B(_12549_), .Y(_12574_));
NAND_g _18562_ (.A(_12573_), .B(_12574_), .Y(_00380_));
NAND_g _18563_ (.A(reg_next_pc[6]), .B(_12543_), .Y(_12575_));
NAND_g _18564_ (.A(_11363_), .B(_12542_), .Y(_12576_));
NAND_g _18565_ (.A(_12575_), .B(_12576_), .Y(_12577_));
NAND_g _18566_ (.A(_11275_), .B(_12577_), .Y(_12578_));
NOT_g _18567_ (.A(_12578_), .Y(_12579_));
NAND_g _18568_ (.A(reg_pc[6]), .B(_12549_), .Y(_12580_));
NAND_g _18569_ (.A(_12578_), .B(_12580_), .Y(_00381_));
NAND_g _18570_ (.A(reg_next_pc[7]), .B(_12543_), .Y(_12581_));
NAND_g _18571_ (.A(_11376_), .B(_12542_), .Y(_12582_));
NAND_g _18572_ (.A(_12581_), .B(_12582_), .Y(_12583_));
NAND_g _18573_ (.A(_11275_), .B(_12583_), .Y(_12584_));
NOT_g _18574_ (.A(_12584_), .Y(_12585_));
NAND_g _18575_ (.A(reg_pc[7]), .B(_12549_), .Y(_12586_));
NAND_g _18576_ (.A(_12584_), .B(_12586_), .Y(_00382_));
NAND_g _18577_ (.A(reg_next_pc[8]), .B(_12543_), .Y(_12587_));
NAND_g _18578_ (.A(_11389_), .B(_12542_), .Y(_12588_));
NAND_g _18579_ (.A(_12587_), .B(_12588_), .Y(_12589_));
AND_g _18580_ (.A(_11275_), .B(_12589_), .Y(_12590_));
NAND_g _18581_ (.A(_11275_), .B(_12589_), .Y(_12591_));
NAND_g _18582_ (.A(reg_pc[8]), .B(_12549_), .Y(_12592_));
NAND_g _18583_ (.A(_12591_), .B(_12592_), .Y(_00383_));
NAND_g _18584_ (.A(reg_next_pc[9]), .B(_12543_), .Y(_12593_));
NAND_g _18585_ (.A(_11402_), .B(_12542_), .Y(_12594_));
NAND_g _18586_ (.A(_12593_), .B(_12594_), .Y(_12595_));
AND_g _18587_ (.A(_11275_), .B(_12595_), .Y(_12596_));
NAND_g _18588_ (.A(_11275_), .B(_12595_), .Y(_12597_));
NAND_g _18589_ (.A(reg_pc[9]), .B(_12549_), .Y(_12598_));
NAND_g _18590_ (.A(_12597_), .B(_12598_), .Y(_00384_));
NAND_g _18591_ (.A(reg_next_pc[10]), .B(_12543_), .Y(_12599_));
NAND_g _18592_ (.A(_11415_), .B(_12542_), .Y(_12600_));
NAND_g _18593_ (.A(_12599_), .B(_12600_), .Y(_12601_));
AND_g _18594_ (.A(_11275_), .B(_12601_), .Y(_12602_));
NAND_g _18595_ (.A(_11275_), .B(_12601_), .Y(_12603_));
NAND_g _18596_ (.A(reg_pc[10]), .B(_12549_), .Y(_12604_));
NAND_g _18597_ (.A(_12603_), .B(_12604_), .Y(_00385_));
NAND_g _18598_ (.A(reg_next_pc[11]), .B(_12543_), .Y(_12605_));
NAND_g _18599_ (.A(_11428_), .B(_12542_), .Y(_12606_));
NAND_g _18600_ (.A(_12605_), .B(_12606_), .Y(_12607_));
AND_g _18601_ (.A(_11275_), .B(_12607_), .Y(_12608_));
NAND_g _18602_ (.A(_11275_), .B(_12607_), .Y(_12609_));
NAND_g _18603_ (.A(reg_pc[11]), .B(_12549_), .Y(_12610_));
NAND_g _18604_ (.A(_12609_), .B(_12610_), .Y(_00386_));
NAND_g _18605_ (.A(reg_next_pc[12]), .B(_12543_), .Y(_12611_));
NAND_g _18606_ (.A(_11441_), .B(_12542_), .Y(_12612_));
NAND_g _18607_ (.A(_12611_), .B(_12612_), .Y(_12613_));
AND_g _18608_ (.A(_11275_), .B(_12613_), .Y(_12614_));
NAND_g _18609_ (.A(_11275_), .B(_12613_), .Y(_12615_));
NAND_g _18610_ (.A(reg_pc[12]), .B(_12549_), .Y(_12616_));
NAND_g _18611_ (.A(_12615_), .B(_12616_), .Y(_00387_));
NAND_g _18612_ (.A(reg_next_pc[13]), .B(_12543_), .Y(_12617_));
NAND_g _18613_ (.A(_11454_), .B(_12542_), .Y(_12618_));
NAND_g _18614_ (.A(_12617_), .B(_12618_), .Y(_12619_));
NAND_g _18615_ (.A(_11275_), .B(_12619_), .Y(_12620_));
NOT_g _18616_ (.A(_12620_), .Y(_12621_));
NAND_g _18617_ (.A(reg_pc[13]), .B(_12549_), .Y(_12622_));
NAND_g _18618_ (.A(_12620_), .B(_12622_), .Y(_00388_));
NAND_g _18619_ (.A(reg_next_pc[14]), .B(_12543_), .Y(_12623_));
NAND_g _18620_ (.A(_11467_), .B(_12542_), .Y(_12624_));
NAND_g _18621_ (.A(_12623_), .B(_12624_), .Y(_12625_));
AND_g _18622_ (.A(_11275_), .B(_12625_), .Y(_12626_));
NAND_g _18623_ (.A(_11275_), .B(_12625_), .Y(_12627_));
NAND_g _18624_ (.A(reg_pc[14]), .B(_12549_), .Y(_12628_));
NAND_g _18625_ (.A(_12627_), .B(_12628_), .Y(_00389_));
NAND_g _18626_ (.A(reg_next_pc[15]), .B(_12543_), .Y(_12629_));
NAND_g _18627_ (.A(_11480_), .B(_12542_), .Y(_12630_));
NAND_g _18628_ (.A(_12629_), .B(_12630_), .Y(_12631_));
NAND_g _18629_ (.A(_11275_), .B(_12631_), .Y(_12632_));
NOT_g _18630_ (.A(_12632_), .Y(_12633_));
NAND_g _18631_ (.A(reg_pc[15]), .B(_12549_), .Y(_12634_));
NAND_g _18632_ (.A(_12632_), .B(_12634_), .Y(_00390_));
NAND_g _18633_ (.A(reg_next_pc[16]), .B(_12543_), .Y(_12635_));
NAND_g _18634_ (.A(_11493_), .B(_12542_), .Y(_12636_));
NAND_g _18635_ (.A(_12635_), .B(_12636_), .Y(_12637_));
AND_g _18636_ (.A(_11275_), .B(_12637_), .Y(_12638_));
NAND_g _18637_ (.A(_11275_), .B(_12637_), .Y(_12639_));
NAND_g _18638_ (.A(reg_pc[16]), .B(_12549_), .Y(_12640_));
NAND_g _18639_ (.A(_12639_), .B(_12640_), .Y(_00391_));
NAND_g _18640_ (.A(reg_next_pc[17]), .B(_12543_), .Y(_12641_));
NAND_g _18641_ (.A(_11506_), .B(_12542_), .Y(_12642_));
NAND_g _18642_ (.A(_12641_), .B(_12642_), .Y(_12643_));
NAND_g _18643_ (.A(_11275_), .B(_12643_), .Y(_12644_));
NOT_g _18644_ (.A(_12644_), .Y(_12645_));
NAND_g _18645_ (.A(reg_pc[17]), .B(_12549_), .Y(_12646_));
NAND_g _18646_ (.A(_12644_), .B(_12646_), .Y(_00392_));
NAND_g _18647_ (.A(reg_next_pc[18]), .B(_12543_), .Y(_12647_));
NAND_g _18648_ (.A(_11519_), .B(_12542_), .Y(_12648_));
NAND_g _18649_ (.A(_12647_), .B(_12648_), .Y(_12649_));
AND_g _18650_ (.A(_11275_), .B(_12649_), .Y(_12650_));
NAND_g _18651_ (.A(_11275_), .B(_12649_), .Y(_12651_));
NAND_g _18652_ (.A(reg_pc[18]), .B(_12549_), .Y(_12652_));
NAND_g _18653_ (.A(_12651_), .B(_12652_), .Y(_00393_));
NAND_g _18654_ (.A(reg_next_pc[19]), .B(_12543_), .Y(_12653_));
NAND_g _18655_ (.A(_11532_), .B(_12542_), .Y(_12654_));
NAND_g _18656_ (.A(_12653_), .B(_12654_), .Y(_12655_));
NAND_g _18657_ (.A(_11275_), .B(_12655_), .Y(_12656_));
NOT_g _18658_ (.A(_12656_), .Y(_12657_));
NAND_g _18659_ (.A(reg_pc[19]), .B(_12549_), .Y(_12658_));
NAND_g _18660_ (.A(_12656_), .B(_12658_), .Y(_00394_));
NAND_g _18661_ (.A(reg_next_pc[20]), .B(_12543_), .Y(_12659_));
NAND_g _18662_ (.A(_11545_), .B(_12542_), .Y(_12660_));
NAND_g _18663_ (.A(_12659_), .B(_12660_), .Y(_12661_));
AND_g _18664_ (.A(_11275_), .B(_12661_), .Y(_12662_));
NAND_g _18665_ (.A(_11275_), .B(_12661_), .Y(_12663_));
NAND_g _18666_ (.A(reg_pc[20]), .B(_12549_), .Y(_12664_));
NAND_g _18667_ (.A(_12663_), .B(_12664_), .Y(_00395_));
NAND_g _18668_ (.A(reg_next_pc[21]), .B(_12543_), .Y(_12665_));
NAND_g _18669_ (.A(_11558_), .B(_12542_), .Y(_12666_));
NAND_g _18670_ (.A(_12665_), .B(_12666_), .Y(_12667_));
NAND_g _18671_ (.A(_11275_), .B(_12667_), .Y(_12668_));
NOT_g _18672_ (.A(_12668_), .Y(_12669_));
NAND_g _18673_ (.A(reg_pc[21]), .B(_12549_), .Y(_12670_));
NAND_g _18674_ (.A(_12668_), .B(_12670_), .Y(_00396_));
NAND_g _18675_ (.A(reg_next_pc[22]), .B(_12543_), .Y(_12671_));
NAND_g _18676_ (.A(_11571_), .B(_12542_), .Y(_12672_));
NAND_g _18677_ (.A(_12671_), .B(_12672_), .Y(_12673_));
AND_g _18678_ (.A(_11275_), .B(_12673_), .Y(_12674_));
NAND_g _18679_ (.A(_11275_), .B(_12673_), .Y(_12675_));
NAND_g _18680_ (.A(reg_pc[22]), .B(_12549_), .Y(_12676_));
NAND_g _18681_ (.A(_12675_), .B(_12676_), .Y(_00397_));
NAND_g _18682_ (.A(reg_next_pc[23]), .B(_12543_), .Y(_12677_));
NAND_g _18683_ (.A(_11584_), .B(_12542_), .Y(_12678_));
NAND_g _18684_ (.A(_12677_), .B(_12678_), .Y(_12679_));
NAND_g _18685_ (.A(_11275_), .B(_12679_), .Y(_12680_));
NAND_g _18686_ (.A(reg_pc[23]), .B(_12549_), .Y(_12681_));
NAND_g _18687_ (.A(_12680_), .B(_12681_), .Y(_00398_));
NAND_g _18688_ (.A(reg_next_pc[24]), .B(_12543_), .Y(_12682_));
NAND_g _18689_ (.A(_11597_), .B(_12542_), .Y(_12683_));
NAND_g _18690_ (.A(_12682_), .B(_12683_), .Y(_12684_));
AND_g _18691_ (.A(_11275_), .B(_12684_), .Y(_12685_));
NAND_g _18692_ (.A(_11275_), .B(_12684_), .Y(_12686_));
NAND_g _18693_ (.A(reg_pc[24]), .B(_12549_), .Y(_12687_));
NAND_g _18694_ (.A(_12686_), .B(_12687_), .Y(_00399_));
NAND_g _18695_ (.A(reg_next_pc[25]), .B(_12543_), .Y(_12688_));
NAND_g _18696_ (.A(_11610_), .B(_12542_), .Y(_12689_));
NAND_g _18697_ (.A(_12688_), .B(_12689_), .Y(_12690_));
NAND_g _18698_ (.A(_11275_), .B(_12690_), .Y(_12691_));
NAND_g _18699_ (.A(reg_pc[25]), .B(_12549_), .Y(_12692_));
NAND_g _18700_ (.A(_12691_), .B(_12692_), .Y(_00400_));
NAND_g _18701_ (.A(reg_next_pc[26]), .B(_12543_), .Y(_12693_));
NAND_g _18702_ (.A(_11623_), .B(_12542_), .Y(_12694_));
NAND_g _18703_ (.A(_12693_), .B(_12694_), .Y(_12695_));
NAND_g _18704_ (.A(_11275_), .B(_12695_), .Y(_12696_));
NOT_g _18705_ (.A(_12696_), .Y(_12697_));
NAND_g _18706_ (.A(reg_pc[26]), .B(_12549_), .Y(_12698_));
NAND_g _18707_ (.A(_12696_), .B(_12698_), .Y(_00401_));
NAND_g _18708_ (.A(reg_next_pc[27]), .B(_12543_), .Y(_12699_));
NAND_g _18709_ (.A(_11636_), .B(_12542_), .Y(_12700_));
NAND_g _18710_ (.A(_12699_), .B(_12700_), .Y(_12701_));
NAND_g _18711_ (.A(_11275_), .B(_12701_), .Y(_12702_));
NAND_g _18712_ (.A(reg_pc[27]), .B(_12549_), .Y(_12703_));
NAND_g _18713_ (.A(_12702_), .B(_12703_), .Y(_00402_));
NAND_g _18714_ (.A(reg_next_pc[28]), .B(_12543_), .Y(_12704_));
NAND_g _18715_ (.A(_11649_), .B(_12542_), .Y(_12705_));
NAND_g _18716_ (.A(_12704_), .B(_12705_), .Y(_12706_));
NAND_g _18717_ (.A(_11275_), .B(_12706_), .Y(_12707_));
NOT_g _18718_ (.A(_12707_), .Y(_12708_));
NAND_g _18719_ (.A(reg_pc[28]), .B(_12549_), .Y(_12709_));
NAND_g _18720_ (.A(_12707_), .B(_12709_), .Y(_00403_));
NAND_g _18721_ (.A(reg_next_pc[29]), .B(_12543_), .Y(_12710_));
NAND_g _18722_ (.A(_11662_), .B(_12542_), .Y(_12711_));
NAND_g _18723_ (.A(_12710_), .B(_12711_), .Y(_12712_));
AND_g _18724_ (.A(_11275_), .B(_12712_), .Y(_12713_));
NAND_g _18725_ (.A(_11275_), .B(_12712_), .Y(_12714_));
NAND_g _18726_ (.A(reg_pc[29]), .B(_12549_), .Y(_12715_));
NAND_g _18727_ (.A(_12714_), .B(_12715_), .Y(_00404_));
NAND_g _18728_ (.A(reg_next_pc[30]), .B(_12543_), .Y(_12716_));
NAND_g _18729_ (.A(_11675_), .B(_12542_), .Y(_12717_));
NAND_g _18730_ (.A(_12716_), .B(_12717_), .Y(_12718_));
NAND_g _18731_ (.A(_11275_), .B(_12718_), .Y(_12719_));
NAND_g _18732_ (.A(reg_pc[30]), .B(_12549_), .Y(_12720_));
NAND_g _18733_ (.A(_12719_), .B(_12720_), .Y(_00405_));
NAND_g _18734_ (.A(reg_next_pc[31]), .B(_12543_), .Y(_12721_));
NAND_g _18735_ (.A(_11688_), .B(_12542_), .Y(_12722_));
NAND_g _18736_ (.A(_12721_), .B(_12722_), .Y(_12723_));
NAND_g _18737_ (.A(_11275_), .B(_12723_), .Y(_12724_));
NAND_g _18738_ (.A(reg_pc[31]), .B(_12549_), .Y(_12725_));
NAND_g _18739_ (.A(_12724_), .B(_12725_), .Y(_00406_));
NAND_g _18740_ (.A(reg_next_pc[1]), .B(_12549_), .Y(_12726_));
AND_g _18741_ (.A(instr_jal), .B(decoded_imm_j[1]), .Y(_12727_));
NAND_g _18742_ (.A(decoder_trigger), .B(_12727_), .Y(_12728_));
XNOR_g _18743_ (.A(_12546_), .B(_12728_), .Y(_12729_));
NAND_g _18744_ (.A(_11275_), .B(_12729_), .Y(_12730_));
NAND_g _18745_ (.A(_12726_), .B(_12730_), .Y(_00407_));
NAND_g _18746_ (.A(reg_next_pc[2]), .B(_12549_), .Y(_12731_));
AND_g _18747_ (.A(decoded_imm_j[1]), .B(_12547_), .Y(_12732_));
NAND_g _18748_ (.A(decoded_imm_j[2]), .B(_12554_), .Y(_12733_));
XNOR_g _18749_ (.A(decoded_imm_j[2]), .B(_12555_), .Y(_12734_));
NAND_g _18750_ (.A(_12732_), .B(_12734_), .Y(_12735_));
XOR_g _18751_ (.A(_12732_), .B(_12734_), .Y(_12736_));
NAND_g _18752_ (.A(instr_jal), .B(_12736_), .Y(_12737_));
NAND_g _18753_ (.A(_10962_), .B(_12555_), .Y(_12738_));
AND_g _18754_ (.A(decoder_trigger), .B(_12738_), .Y(_12739_));
NAND_g _18755_ (.A(_12737_), .B(_12739_), .Y(_12740_));
NAND_g _18756_ (.A(resetn), .B(launch_next_insn), .Y(_12741_));
NAND_g _18757_ (.A(_12555_), .B(_12741_), .Y(_12742_));
NAND_g _18758_ (.A(_12740_), .B(_12742_), .Y(_12743_));
NAND_g _18759_ (.A(_12731_), .B(_12743_), .Y(_00408_));
NAND_g _18760_ (.A(reg_next_pc[3]), .B(_12549_), .Y(_12744_));
NAND_g _18761_ (.A(_12733_), .B(_12735_), .Y(_12745_));
NAND_g _18762_ (.A(decoded_imm_j[3]), .B(_12560_), .Y(_12746_));
NAND_g _18763_ (.A(_10976_), .B(_12561_), .Y(_12747_));
XNOR_g _18764_ (.A(decoded_imm_j[3]), .B(_12560_), .Y(_12748_));
XNOR_g _18765_ (.A(_12745_), .B(_12748_), .Y(_12749_));
NAND_g _18766_ (.A(instr_jal), .B(_12749_), .Y(_12750_));
AND_g _18767_ (.A(_12553_), .B(_12560_), .Y(_12751_));
NAND_g _18768_ (.A(_12554_), .B(_12559_), .Y(_12752_));
NAND_g _18769_ (.A(_10962_), .B(_12752_), .Y(_12753_));
AND_g _18770_ (.A(decoder_trigger), .B(_12753_), .Y(_12754_));
NAND_g _18771_ (.A(_12750_), .B(_12754_), .Y(_12755_));
NAND_g _18772_ (.A(_11275_), .B(_12739_), .Y(_12756_));
NAND_g _18773_ (.A(_12561_), .B(_12756_), .Y(_12757_));
NAND_g _18774_ (.A(_12755_), .B(_12757_), .Y(_12758_));
NAND_g _18775_ (.A(_12744_), .B(_12758_), .Y(_00409_));
NAND_g _18776_ (.A(reg_next_pc[4]), .B(_12549_), .Y(_12759_));
NAND_g _18777_ (.A(decoded_imm_j[4]), .B(_12567_), .Y(_12760_));
XNOR_g _18778_ (.A(decoded_imm_j[4]), .B(_12566_), .Y(_12761_));
NAND_g _18779_ (.A(_12745_), .B(_12747_), .Y(_12762_));
NAND_g _18780_ (.A(_12746_), .B(_12762_), .Y(_12763_));
NAND_g _18781_ (.A(_12761_), .B(_12763_), .Y(_12764_));
XOR_g _18782_ (.A(_12761_), .B(_12763_), .Y(_12765_));
AND_g _18783_ (.A(_12566_), .B(_12752_), .Y(_12766_));
AND_g _18784_ (.A(_12565_), .B(_12751_), .Y(_12767_));
NOR_g _18785_ (.A(_12766_), .B(_12767_), .Y(_12768_));
NAND_g _18786_ (.A(instr_jal), .B(_12765_), .Y(_12769_));
NAND_g _18787_ (.A(_10962_), .B(_12768_), .Y(_12770_));
AND_g _18788_ (.A(decoder_trigger), .B(_12770_), .Y(_12771_));
NAND_g _18789_ (.A(_12769_), .B(_12771_), .Y(_12772_));
NAND_g _18790_ (.A(_12566_), .B(_12741_), .Y(_12773_));
NAND_g _18791_ (.A(_12772_), .B(_12773_), .Y(_12774_));
NAND_g _18792_ (.A(_12759_), .B(_12774_), .Y(_00410_));
NAND_g _18793_ (.A(reg_next_pc[5]), .B(_12549_), .Y(_12775_));
NAND_g _18794_ (.A(_12760_), .B(_12764_), .Y(_12776_));
NAND_g _18795_ (.A(decoded_imm_j[5]), .B(_12572_), .Y(_12777_));
XOR_g _18796_ (.A(decoded_imm_j[5]), .B(_12572_), .Y(_12778_));
NAND_g _18797_ (.A(_12776_), .B(_12778_), .Y(_12779_));
XNOR_g _18798_ (.A(_12776_), .B(_12778_), .Y(_12780_));
NAND_g _18799_ (.A(instr_jal), .B(_12780_), .Y(_12781_));
AND_g _18800_ (.A(_12572_), .B(_12767_), .Y(_12782_));
XNOR_g _18801_ (.A(_12572_), .B(_12767_), .Y(_12783_));
NAND_g _18802_ (.A(_10962_), .B(_12783_), .Y(_12784_));
NAND_g _18803_ (.A(_12781_), .B(_12784_), .Y(_12785_));
NAND_g _18804_ (.A(decoder_trigger), .B(_12785_), .Y(_12786_));
NAND_g _18805_ (.A(_12573_), .B(_12741_), .Y(_12787_));
NAND_g _18806_ (.A(_12786_), .B(_12787_), .Y(_12788_));
NAND_g _18807_ (.A(_12775_), .B(_12788_), .Y(_00411_));
NAND_g _18808_ (.A(reg_next_pc[6]), .B(_12549_), .Y(_12789_));
NAND_g _18809_ (.A(_12777_), .B(_12779_), .Y(_12790_));
NAND_g _18810_ (.A(decoded_imm_j[6]), .B(_12579_), .Y(_12791_));
XNOR_g _18811_ (.A(decoded_imm_j[6]), .B(_12578_), .Y(_12792_));
NAND_g _18812_ (.A(_12790_), .B(_12792_), .Y(_12793_));
XOR_g _18813_ (.A(_12790_), .B(_12792_), .Y(_12794_));
NAND_g _18814_ (.A(instr_jal), .B(_12794_), .Y(_12795_));
AND_g _18815_ (.A(_12577_), .B(_12782_), .Y(_12796_));
NOR_g _18816_ (.A(_12579_), .B(_12782_), .Y(_12797_));
NOR_g _18817_ (.A(_12796_), .B(_12797_), .Y(_12798_));
NAND_g _18818_ (.A(_10962_), .B(_12798_), .Y(_12799_));
AND_g _18819_ (.A(decoder_trigger), .B(_12799_), .Y(_12800_));
NAND_g _18820_ (.A(_12795_), .B(_12800_), .Y(_12801_));
NAND_g _18821_ (.A(_12578_), .B(_12741_), .Y(_12802_));
NAND_g _18822_ (.A(_12801_), .B(_12802_), .Y(_12803_));
NAND_g _18823_ (.A(_12789_), .B(_12803_), .Y(_00412_));
NAND_g _18824_ (.A(reg_next_pc[7]), .B(_12549_), .Y(_12804_));
NAND_g _18825_ (.A(_12791_), .B(_12793_), .Y(_12805_));
NAND_g _18826_ (.A(decoded_imm_j[7]), .B(_12585_), .Y(_12806_));
NAND_g _18827_ (.A(_11137_), .B(_12584_), .Y(_12807_));
XNOR_g _18828_ (.A(_11137_), .B(_12584_), .Y(_12808_));
XNOR_g _18829_ (.A(_12805_), .B(_12808_), .Y(_12809_));
NAND_g _18830_ (.A(instr_jal), .B(_12809_), .Y(_12810_));
AND_g _18831_ (.A(_12585_), .B(_12796_), .Y(_12811_));
XNOR_g _18832_ (.A(_12584_), .B(_12796_), .Y(_12812_));
NAND_g _18833_ (.A(_10962_), .B(_12812_), .Y(_12813_));
AND_g _18834_ (.A(decoder_trigger), .B(_12810_), .Y(_12814_));
NAND_g _18835_ (.A(_12813_), .B(_12814_), .Y(_12815_));
NAND_g _18836_ (.A(_12584_), .B(_12741_), .Y(_12816_));
NAND_g _18837_ (.A(_12815_), .B(_12816_), .Y(_12817_));
NAND_g _18838_ (.A(_12804_), .B(_12817_), .Y(_00413_));
NAND_g _18839_ (.A(reg_next_pc[8]), .B(_12549_), .Y(_12818_));
NAND_g _18840_ (.A(decoded_imm_j[8]), .B(_12590_), .Y(_12819_));
XNOR_g _18841_ (.A(decoded_imm_j[8]), .B(_12591_), .Y(_12820_));
NAND_g _18842_ (.A(_12805_), .B(_12807_), .Y(_12821_));
NAND_g _18843_ (.A(_12806_), .B(_12821_), .Y(_12822_));
NAND_g _18844_ (.A(_12820_), .B(_12822_), .Y(_12823_));
XOR_g _18845_ (.A(_12820_), .B(_12822_), .Y(_12824_));
NAND_g _18846_ (.A(instr_jal), .B(_12824_), .Y(_12825_));
AND_g _18847_ (.A(_12589_), .B(_12811_), .Y(_12826_));
NOR_g _18848_ (.A(_12590_), .B(_12811_), .Y(_12827_));
NOR_g _18849_ (.A(_12826_), .B(_12827_), .Y(_12828_));
NAND_g _18850_ (.A(_10962_), .B(_12828_), .Y(_12829_));
AND_g _18851_ (.A(decoder_trigger), .B(_12829_), .Y(_12830_));
NAND_g _18852_ (.A(_12825_), .B(_12830_), .Y(_12831_));
NAND_g _18853_ (.A(_12591_), .B(_12741_), .Y(_12832_));
NAND_g _18854_ (.A(_12831_), .B(_12832_), .Y(_12833_));
NAND_g _18855_ (.A(_12818_), .B(_12833_), .Y(_00414_));
NAND_g _18856_ (.A(reg_next_pc[9]), .B(_12549_), .Y(_12834_));
NAND_g _18857_ (.A(_12819_), .B(_12823_), .Y(_12835_));
NAND_g _18858_ (.A(decoded_imm_j[9]), .B(_12596_), .Y(_12836_));
NOR_g _18859_ (.A(decoded_imm_j[9]), .B(_12596_), .Y(_12837_));
NOT_g _18860_ (.A(_12837_), .Y(_12838_));
XNOR_g _18861_ (.A(decoded_imm_j[9]), .B(_12596_), .Y(_12839_));
XNOR_g _18862_ (.A(_12835_), .B(_12839_), .Y(_12840_));
NAND_g _18863_ (.A(instr_jal), .B(_12840_), .Y(_12841_));
AND_g _18864_ (.A(_12596_), .B(_12826_), .Y(_12842_));
XNOR_g _18865_ (.A(_12597_), .B(_12826_), .Y(_12843_));
NAND_g _18866_ (.A(_10962_), .B(_12843_), .Y(_12844_));
AND_g _18867_ (.A(decoder_trigger), .B(_12841_), .Y(_12845_));
NAND_g _18868_ (.A(_12844_), .B(_12845_), .Y(_12846_));
NAND_g _18869_ (.A(_12597_), .B(_12741_), .Y(_12847_));
NAND_g _18870_ (.A(_12846_), .B(_12847_), .Y(_12848_));
NAND_g _18871_ (.A(_12834_), .B(_12848_), .Y(_00415_));
NAND_g _18872_ (.A(reg_next_pc[10]), .B(_12549_), .Y(_12849_));
NAND_g _18873_ (.A(decoded_imm_j[10]), .B(_12602_), .Y(_12850_));
XNOR_g _18874_ (.A(decoded_imm_j[10]), .B(_12603_), .Y(_12851_));
NAND_g _18875_ (.A(_12835_), .B(_12838_), .Y(_12852_));
NAND_g _18876_ (.A(_12836_), .B(_12852_), .Y(_12853_));
NAND_g _18877_ (.A(_12851_), .B(_12853_), .Y(_12854_));
XOR_g _18878_ (.A(_12851_), .B(_12853_), .Y(_12855_));
NAND_g _18879_ (.A(instr_jal), .B(_12855_), .Y(_12856_));
AND_g _18880_ (.A(_12601_), .B(_12842_), .Y(_12857_));
NOR_g _18881_ (.A(_12602_), .B(_12842_), .Y(_12858_));
NOR_g _18882_ (.A(_12857_), .B(_12858_), .Y(_12859_));
NAND_g _18883_ (.A(_10962_), .B(_12859_), .Y(_12860_));
AND_g _18884_ (.A(decoder_trigger), .B(_12860_), .Y(_12861_));
NAND_g _18885_ (.A(_12856_), .B(_12861_), .Y(_12862_));
NAND_g _18886_ (.A(_12603_), .B(_12741_), .Y(_12863_));
NAND_g _18887_ (.A(_12862_), .B(_12863_), .Y(_12864_));
NAND_g _18888_ (.A(_12849_), .B(_12864_), .Y(_00416_));
NAND_g _18889_ (.A(reg_next_pc[11]), .B(_12549_), .Y(_12865_));
AND_g _18890_ (.A(_12850_), .B(_12854_), .Y(_12866_));
NAND_g _18891_ (.A(decoded_imm_j[11]), .B(_12608_), .Y(_12867_));
NOR_g _18892_ (.A(decoded_imm_j[11]), .B(_12608_), .Y(_12868_));
XNOR_g _18893_ (.A(decoded_imm_j[11]), .B(_12609_), .Y(_12869_));
XNOR_g _18894_ (.A(_12866_), .B(_12869_), .Y(_12870_));
NAND_g _18895_ (.A(instr_jal), .B(_12870_), .Y(_12871_));
AND_g _18896_ (.A(_12608_), .B(_12857_), .Y(_12872_));
XNOR_g _18897_ (.A(_12609_), .B(_12857_), .Y(_12873_));
NAND_g _18898_ (.A(_10962_), .B(_12873_), .Y(_12874_));
AND_g _18899_ (.A(decoder_trigger), .B(_12874_), .Y(_12875_));
NAND_g _18900_ (.A(_12871_), .B(_12875_), .Y(_12876_));
NAND_g _18901_ (.A(_12609_), .B(_12741_), .Y(_12877_));
NAND_g _18902_ (.A(_12876_), .B(_12877_), .Y(_12878_));
NAND_g _18903_ (.A(_12865_), .B(_12878_), .Y(_00417_));
NAND_g _18904_ (.A(reg_next_pc[12]), .B(_12549_), .Y(_12879_));
NAND_g _18905_ (.A(decoded_imm_j[12]), .B(_12614_), .Y(_12880_));
XNOR_g _18906_ (.A(decoded_imm_j[12]), .B(_12615_), .Y(_12881_));
AND_g _18907_ (.A(_12866_), .B(_12867_), .Y(_12882_));
NOR_g _18908_ (.A(_12868_), .B(_12882_), .Y(_12883_));
NAND_g _18909_ (.A(_12881_), .B(_12883_), .Y(_12884_));
XOR_g _18910_ (.A(_12881_), .B(_12883_), .Y(_12885_));
NAND_g _18911_ (.A(instr_jal), .B(_12885_), .Y(_12886_));
AND_g _18912_ (.A(_12613_), .B(_12872_), .Y(_12887_));
NOR_g _18913_ (.A(_12614_), .B(_12872_), .Y(_12888_));
NOR_g _18914_ (.A(_12887_), .B(_12888_), .Y(_12889_));
NAND_g _18915_ (.A(_10962_), .B(_12889_), .Y(_12890_));
AND_g _18916_ (.A(decoder_trigger), .B(_12890_), .Y(_12891_));
NAND_g _18917_ (.A(_12886_), .B(_12891_), .Y(_12892_));
NAND_g _18918_ (.A(_12615_), .B(_12741_), .Y(_12893_));
NAND_g _18919_ (.A(_12892_), .B(_12893_), .Y(_12894_));
NAND_g _18920_ (.A(_12879_), .B(_12894_), .Y(_00418_));
NAND_g _18921_ (.A(reg_next_pc[13]), .B(_12549_), .Y(_12895_));
NAND_g _18922_ (.A(_12880_), .B(_12884_), .Y(_12896_));
NAND_g _18923_ (.A(decoded_imm_j[13]), .B(_12621_), .Y(_12897_));
NAND_g _18924_ (.A(_11155_), .B(_12620_), .Y(_12898_));
XNOR_g _18925_ (.A(_11155_), .B(_12620_), .Y(_12899_));
XNOR_g _18926_ (.A(_12896_), .B(_12899_), .Y(_12900_));
NAND_g _18927_ (.A(instr_jal), .B(_12900_), .Y(_12901_));
AND_g _18928_ (.A(_12621_), .B(_12887_), .Y(_12902_));
XNOR_g _18929_ (.A(_12620_), .B(_12887_), .Y(_12903_));
NAND_g _18930_ (.A(_10962_), .B(_12903_), .Y(_12904_));
AND_g _18931_ (.A(decoder_trigger), .B(_12901_), .Y(_12905_));
NAND_g _18932_ (.A(_12904_), .B(_12905_), .Y(_12906_));
NAND_g _18933_ (.A(_12620_), .B(_12741_), .Y(_12907_));
NAND_g _18934_ (.A(_12906_), .B(_12907_), .Y(_12908_));
NAND_g _18935_ (.A(_12895_), .B(_12908_), .Y(_00419_));
NAND_g _18936_ (.A(reg_next_pc[14]), .B(_12549_), .Y(_12909_));
NAND_g _18937_ (.A(decoded_imm_j[14]), .B(_12626_), .Y(_12910_));
XNOR_g _18938_ (.A(decoded_imm_j[14]), .B(_12627_), .Y(_12911_));
NAND_g _18939_ (.A(_12896_), .B(_12898_), .Y(_12912_));
NAND_g _18940_ (.A(_12897_), .B(_12912_), .Y(_12913_));
NAND_g _18941_ (.A(_12911_), .B(_12913_), .Y(_12914_));
XOR_g _18942_ (.A(_12911_), .B(_12913_), .Y(_12915_));
NAND_g _18943_ (.A(instr_jal), .B(_12915_), .Y(_12916_));
AND_g _18944_ (.A(_12625_), .B(_12902_), .Y(_12917_));
NOR_g _18945_ (.A(_12626_), .B(_12902_), .Y(_12918_));
NOR_g _18946_ (.A(_12917_), .B(_12918_), .Y(_12919_));
NAND_g _18947_ (.A(_10962_), .B(_12919_), .Y(_12920_));
AND_g _18948_ (.A(decoder_trigger), .B(_12920_), .Y(_12921_));
NAND_g _18949_ (.A(_12916_), .B(_12921_), .Y(_12922_));
NAND_g _18950_ (.A(_12627_), .B(_12741_), .Y(_12923_));
NAND_g _18951_ (.A(_12922_), .B(_12923_), .Y(_12924_));
NAND_g _18952_ (.A(_12909_), .B(_12924_), .Y(_00420_));
NAND_g _18953_ (.A(reg_next_pc[15]), .B(_12549_), .Y(_12925_));
NAND_g _18954_ (.A(decoded_imm_j[15]), .B(_12633_), .Y(_12926_));
NAND_g _18955_ (.A(_11046_), .B(_12632_), .Y(_12927_));
XNOR_g _18956_ (.A(_11046_), .B(_12632_), .Y(_12928_));
NAND_g _18957_ (.A(_12910_), .B(_12914_), .Y(_12929_));
XNOR_g _18958_ (.A(_12928_), .B(_12929_), .Y(_12930_));
NAND_g _18959_ (.A(instr_jal), .B(_12930_), .Y(_12931_));
AND_g _18960_ (.A(_12633_), .B(_12917_), .Y(_12932_));
XNOR_g _18961_ (.A(_12632_), .B(_12917_), .Y(_12933_));
NAND_g _18962_ (.A(_10962_), .B(_12933_), .Y(_12934_));
AND_g _18963_ (.A(decoder_trigger), .B(_12931_), .Y(_12935_));
NAND_g _18964_ (.A(_12934_), .B(_12935_), .Y(_12936_));
NAND_g _18965_ (.A(_12632_), .B(_12741_), .Y(_12937_));
NAND_g _18966_ (.A(_12936_), .B(_12937_), .Y(_12938_));
NAND_g _18967_ (.A(_12925_), .B(_12938_), .Y(_00421_));
NAND_g _18968_ (.A(reg_next_pc[16]), .B(_12549_), .Y(_12939_));
NAND_g _18969_ (.A(decoded_imm_j[16]), .B(_12638_), .Y(_12940_));
XNOR_g _18970_ (.A(decoded_imm_j[16]), .B(_12639_), .Y(_12941_));
NAND_g _18971_ (.A(_12927_), .B(_12929_), .Y(_12942_));
NAND_g _18972_ (.A(_12926_), .B(_12942_), .Y(_12943_));
NAND_g _18973_ (.A(_12941_), .B(_12943_), .Y(_12944_));
XOR_g _18974_ (.A(_12941_), .B(_12943_), .Y(_12945_));
NAND_g _18975_ (.A(instr_jal), .B(_12945_), .Y(_12946_));
AND_g _18976_ (.A(_12637_), .B(_12932_), .Y(_12947_));
NOR_g _18977_ (.A(_12638_), .B(_12932_), .Y(_12948_));
NOR_g _18978_ (.A(_12947_), .B(_12948_), .Y(_12949_));
NAND_g _18979_ (.A(_10962_), .B(_12949_), .Y(_12950_));
AND_g _18980_ (.A(decoder_trigger), .B(_12950_), .Y(_12951_));
NAND_g _18981_ (.A(_12946_), .B(_12951_), .Y(_12952_));
NAND_g _18982_ (.A(_12639_), .B(_12741_), .Y(_12953_));
NAND_g _18983_ (.A(_12952_), .B(_12953_), .Y(_12954_));
NAND_g _18984_ (.A(_12939_), .B(_12954_), .Y(_00422_));
NAND_g _18985_ (.A(reg_next_pc[17]), .B(_12549_), .Y(_12955_));
NAND_g _18986_ (.A(decoded_imm_j[17]), .B(_12645_), .Y(_12956_));
NAND_g _18987_ (.A(_11047_), .B(_12644_), .Y(_12957_));
XNOR_g _18988_ (.A(_11047_), .B(_12644_), .Y(_12958_));
NAND_g _18989_ (.A(_12940_), .B(_12944_), .Y(_12959_));
XNOR_g _18990_ (.A(_12958_), .B(_12959_), .Y(_12960_));
NAND_g _18991_ (.A(instr_jal), .B(_12960_), .Y(_12961_));
AND_g _18992_ (.A(_12645_), .B(_12947_), .Y(_12962_));
XNOR_g _18993_ (.A(_12644_), .B(_12947_), .Y(_12963_));
NAND_g _18994_ (.A(_10962_), .B(_12963_), .Y(_12964_));
AND_g _18995_ (.A(decoder_trigger), .B(_12964_), .Y(_12965_));
NAND_g _18996_ (.A(_12961_), .B(_12965_), .Y(_12966_));
NAND_g _18997_ (.A(_12644_), .B(_12741_), .Y(_12967_));
NAND_g _18998_ (.A(_12966_), .B(_12967_), .Y(_12968_));
NAND_g _18999_ (.A(_12955_), .B(_12968_), .Y(_00423_));
NAND_g _19000_ (.A(reg_next_pc[18]), .B(_12549_), .Y(_12969_));
NAND_g _19001_ (.A(decoded_imm_j[18]), .B(_12650_), .Y(_12970_));
XNOR_g _19002_ (.A(decoded_imm_j[18]), .B(_12651_), .Y(_12971_));
NAND_g _19003_ (.A(_12957_), .B(_12959_), .Y(_12972_));
NAND_g _19004_ (.A(_12956_), .B(_12972_), .Y(_12973_));
NAND_g _19005_ (.A(_12971_), .B(_12973_), .Y(_12974_));
XOR_g _19006_ (.A(_12971_), .B(_12973_), .Y(_12975_));
NAND_g _19007_ (.A(instr_jal), .B(_12975_), .Y(_12976_));
NAND_g _19008_ (.A(_12649_), .B(_12962_), .Y(_12977_));
NOT_g _19009_ (.A(_12977_), .Y(_12978_));
NOR_g _19010_ (.A(_12650_), .B(_12962_), .Y(_12979_));
NOR_g _19011_ (.A(instr_jal), .B(_12979_), .Y(_12980_));
NAND_g _19012_ (.A(_12977_), .B(_12980_), .Y(_12981_));
AND_g _19013_ (.A(decoder_trigger), .B(_12981_), .Y(_12982_));
NAND_g _19014_ (.A(_12976_), .B(_12982_), .Y(_12983_));
NAND_g _19015_ (.A(_12651_), .B(_12741_), .Y(_12984_));
NAND_g _19016_ (.A(_12983_), .B(_12984_), .Y(_12985_));
NAND_g _19017_ (.A(_12969_), .B(_12985_), .Y(_00424_));
NAND_g _19018_ (.A(reg_next_pc[19]), .B(_12549_), .Y(_12986_));
NAND_g _19019_ (.A(_12970_), .B(_12974_), .Y(_12987_));
NOT_g _19020_ (.A(_12987_), .Y(_12988_));
NAND_g _19021_ (.A(decoded_imm_j[19]), .B(_12657_), .Y(_12989_));
NAND_g _19022_ (.A(_11048_), .B(_12656_), .Y(_12990_));
XNOR_g _19023_ (.A(_11048_), .B(_12656_), .Y(_12991_));
XNOR_g _19024_ (.A(_12987_), .B(_12991_), .Y(_12992_));
NAND_g _19025_ (.A(instr_jal), .B(_12992_), .Y(_12993_));
NAND_g _19026_ (.A(_12656_), .B(_12977_), .Y(_12994_));
AND_g _19027_ (.A(_12655_), .B(_12978_), .Y(_12995_));
NOR_g _19028_ (.A(instr_jal), .B(_12995_), .Y(_12996_));
NAND_g _19029_ (.A(_12994_), .B(_12996_), .Y(_12997_));
AND_g _19030_ (.A(decoder_trigger), .B(_12997_), .Y(_12998_));
NAND_g _19031_ (.A(_12993_), .B(_12998_), .Y(_12999_));
NAND_g _19032_ (.A(_12656_), .B(_12741_), .Y(_13000_));
NAND_g _19033_ (.A(_12999_), .B(_13000_), .Y(_13001_));
NAND_g _19034_ (.A(_12986_), .B(_13001_), .Y(_00425_));
NAND_g _19035_ (.A(reg_next_pc[20]), .B(_12549_), .Y(_13002_));
AND_g _19036_ (.A(decoded_imm_j[31]), .B(_12662_), .Y(_13003_));
XNOR_g _19037_ (.A(decoded_imm_j[31]), .B(_12662_), .Y(_13004_));
NAND_g _19038_ (.A(_12988_), .B(_12989_), .Y(_13005_));
NAND_g _19039_ (.A(_12990_), .B(_13005_), .Y(_13006_));
NAND_g _19040_ (.A(_12987_), .B(_12990_), .Y(_13007_));
NAND_g _19041_ (.A(_12989_), .B(_13007_), .Y(_13008_));
NOR_g _19042_ (.A(_13004_), .B(_13006_), .Y(_13009_));
XNOR_g _19043_ (.A(_13004_), .B(_13008_), .Y(_13010_));
NAND_g _19044_ (.A(instr_jal), .B(_13010_), .Y(_13011_));
AND_g _19045_ (.A(_12662_), .B(_12995_), .Y(_13012_));
XNOR_g _19046_ (.A(_12663_), .B(_12995_), .Y(_13013_));
NAND_g _19047_ (.A(_10962_), .B(_13013_), .Y(_13014_));
AND_g _19048_ (.A(decoder_trigger), .B(_13014_), .Y(_13015_));
NAND_g _19049_ (.A(_13011_), .B(_13015_), .Y(_13016_));
NAND_g _19050_ (.A(_12663_), .B(_12741_), .Y(_13017_));
NAND_g _19051_ (.A(_13016_), .B(_13017_), .Y(_13018_));
NAND_g _19052_ (.A(_13002_), .B(_13018_), .Y(_00426_));
NAND_g _19053_ (.A(reg_next_pc[21]), .B(_12549_), .Y(_13019_));
NOR_g _19054_ (.A(_13003_), .B(_13009_), .Y(_13020_));
NOR_g _19055_ (.A(_11138_), .B(_12668_), .Y(_13021_));
XNOR_g _19056_ (.A(decoded_imm_j[31]), .B(_12668_), .Y(_13022_));
XNOR_g _19057_ (.A(_13020_), .B(_13022_), .Y(_13023_));
NAND_g _19058_ (.A(instr_jal), .B(_13023_), .Y(_13024_));
NOR_g _19059_ (.A(_12669_), .B(_13012_), .Y(_13025_));
AND_g _19060_ (.A(_12667_), .B(_13012_), .Y(_13026_));
NOR_g _19061_ (.A(_13025_), .B(_13026_), .Y(_13027_));
NAND_g _19062_ (.A(_10962_), .B(_13027_), .Y(_13028_));
AND_g _19063_ (.A(decoder_trigger), .B(_13028_), .Y(_13029_));
NAND_g _19064_ (.A(_13024_), .B(_13029_), .Y(_13030_));
NAND_g _19065_ (.A(_12668_), .B(_12741_), .Y(_13031_));
NAND_g _19066_ (.A(_13030_), .B(_13031_), .Y(_13032_));
NAND_g _19067_ (.A(_13019_), .B(_13032_), .Y(_00427_));
NAND_g _19068_ (.A(reg_next_pc[22]), .B(_12549_), .Y(_13033_));
NAND_g _19069_ (.A(_13009_), .B(_13022_), .Y(_13034_));
NOR_g _19070_ (.A(_13003_), .B(_13021_), .Y(_13035_));
NAND_g _19071_ (.A(_13034_), .B(_13035_), .Y(_13036_));
NAND_g _19072_ (.A(decoded_imm_j[31]), .B(_12674_), .Y(_13037_));
XNOR_g _19073_ (.A(_11138_), .B(_12674_), .Y(_13038_));
NAND_g _19074_ (.A(_13036_), .B(_13038_), .Y(_13039_));
XOR_g _19075_ (.A(_13036_), .B(_13038_), .Y(_13040_));
NAND_g _19076_ (.A(instr_jal), .B(_13040_), .Y(_13041_));
AND_g _19077_ (.A(_12674_), .B(_13026_), .Y(_13042_));
NAND_g _19078_ (.A(_12674_), .B(_13026_), .Y(_13043_));
XNOR_g _19079_ (.A(_12675_), .B(_13026_), .Y(_13044_));
NAND_g _19080_ (.A(_10962_), .B(_13044_), .Y(_13045_));
AND_g _19081_ (.A(decoder_trigger), .B(_13045_), .Y(_13046_));
NAND_g _19082_ (.A(_13041_), .B(_13046_), .Y(_13047_));
NAND_g _19083_ (.A(_12675_), .B(_12741_), .Y(_13048_));
NAND_g _19084_ (.A(_13047_), .B(_13048_), .Y(_13049_));
NAND_g _19085_ (.A(_13033_), .B(_13049_), .Y(_00428_));
NAND_g _19086_ (.A(reg_next_pc[23]), .B(_12549_), .Y(_13050_));
NAND_g _19087_ (.A(_13037_), .B(_13039_), .Y(_13051_));
XNOR_g _19088_ (.A(_11138_), .B(_12680_), .Y(_13052_));
XNOR_g _19089_ (.A(_13051_), .B(_13052_), .Y(_13053_));
NAND_g _19090_ (.A(instr_jal), .B(_13053_), .Y(_13054_));
AND_g _19091_ (.A(_12680_), .B(_13043_), .Y(_13055_));
AND_g _19092_ (.A(_12679_), .B(_13042_), .Y(_13056_));
NOR_g _19093_ (.A(_13055_), .B(_13056_), .Y(_13057_));
NAND_g _19094_ (.A(_10962_), .B(_13057_), .Y(_13058_));
AND_g _19095_ (.A(decoder_trigger), .B(_13058_), .Y(_13059_));
NAND_g _19096_ (.A(_13054_), .B(_13059_), .Y(_13060_));
NAND_g _19097_ (.A(_12680_), .B(_12741_), .Y(_13061_));
NAND_g _19098_ (.A(_13060_), .B(_13061_), .Y(_13062_));
NAND_g _19099_ (.A(_13050_), .B(_13062_), .Y(_00429_));
NAND_g _19100_ (.A(reg_next_pc[24]), .B(_12549_), .Y(_13063_));
AND_g _19101_ (.A(_12663_), .B(_12668_), .Y(_13064_));
AND_g _19102_ (.A(_12675_), .B(_12680_), .Y(_13065_));
NAND_g _19103_ (.A(_13064_), .B(_13065_), .Y(_13066_));
NAND_g _19104_ (.A(decoded_imm_j[31]), .B(_13066_), .Y(_13067_));
NOR_g _19105_ (.A(_13034_), .B(_13052_), .Y(_13068_));
NAND_g _19106_ (.A(_13038_), .B(_13068_), .Y(_13069_));
AND_g _19107_ (.A(_13067_), .B(_13069_), .Y(_13070_));
AND_g _19108_ (.A(decoded_imm_j[31]), .B(_12685_), .Y(_13071_));
XNOR_g _19109_ (.A(decoded_imm_j[31]), .B(_12685_), .Y(_13072_));
NOR_g _19110_ (.A(_13070_), .B(_13072_), .Y(_13073_));
XOR_g _19111_ (.A(_13070_), .B(_13072_), .Y(_13074_));
NAND_g _19112_ (.A(instr_jal), .B(_13074_), .Y(_13075_));
AND_g _19113_ (.A(_12685_), .B(_13056_), .Y(_13076_));
NAND_g _19114_ (.A(_12685_), .B(_13056_), .Y(_13077_));
XNOR_g _19115_ (.A(_12686_), .B(_13056_), .Y(_13078_));
NAND_g _19116_ (.A(_10962_), .B(_13078_), .Y(_13079_));
AND_g _19117_ (.A(decoder_trigger), .B(_13079_), .Y(_13080_));
NAND_g _19118_ (.A(_13075_), .B(_13080_), .Y(_13081_));
NAND_g _19119_ (.A(_12686_), .B(_12741_), .Y(_13082_));
NAND_g _19120_ (.A(_13081_), .B(_13082_), .Y(_13083_));
NAND_g _19121_ (.A(_13063_), .B(_13083_), .Y(_00430_));
NOR_g _19122_ (.A(_13071_), .B(_13073_), .Y(_13084_));
NOR_g _19123_ (.A(_11138_), .B(_12691_), .Y(_13085_));
XNOR_g _19124_ (.A(decoded_imm_j[31]), .B(_12691_), .Y(_13086_));
XNOR_g _19125_ (.A(_13084_), .B(_13086_), .Y(_13087_));
NAND_g _19126_ (.A(instr_jal), .B(_13087_), .Y(_13088_));
AND_g _19127_ (.A(_12691_), .B(_13077_), .Y(_13089_));
AND_g _19128_ (.A(_12690_), .B(_13076_), .Y(_13090_));
NOR_g _19129_ (.A(_13089_), .B(_13090_), .Y(_13091_));
NAND_g _19130_ (.A(_10962_), .B(_13091_), .Y(_13092_));
AND_g _19131_ (.A(decoder_trigger), .B(_13092_), .Y(_13093_));
NAND_g _19132_ (.A(_13088_), .B(_13093_), .Y(_13094_));
NAND_g _19133_ (.A(_12691_), .B(_12741_), .Y(_13095_));
NAND_g _19134_ (.A(_13094_), .B(_13095_), .Y(_13096_));
NAND_g _19135_ (.A(reg_next_pc[25]), .B(_12549_), .Y(_13097_));
NAND_g _19136_ (.A(_13096_), .B(_13097_), .Y(_00431_));
NAND_g _19137_ (.A(reg_next_pc[26]), .B(_12549_), .Y(_13098_));
NAND_g _19138_ (.A(_13073_), .B(_13086_), .Y(_13099_));
NOR_g _19139_ (.A(_13071_), .B(_13085_), .Y(_13100_));
NAND_g _19140_ (.A(_13099_), .B(_13100_), .Y(_13101_));
NAND_g _19141_ (.A(decoded_imm_j[31]), .B(_12697_), .Y(_13102_));
XNOR_g _19142_ (.A(decoded_imm_j[31]), .B(_12696_), .Y(_13103_));
NAND_g _19143_ (.A(_13101_), .B(_13103_), .Y(_13104_));
XOR_g _19144_ (.A(_13101_), .B(_13103_), .Y(_13105_));
NAND_g _19145_ (.A(instr_jal), .B(_13105_), .Y(_13106_));
AND_g _19146_ (.A(_12697_), .B(_13090_), .Y(_13107_));
NOT_g _19147_ (.A(_13107_), .Y(_13108_));
XNOR_g _19148_ (.A(_12696_), .B(_13090_), .Y(_13109_));
NAND_g _19149_ (.A(_10962_), .B(_13109_), .Y(_13110_));
AND_g _19150_ (.A(decoder_trigger), .B(_13110_), .Y(_13111_));
NAND_g _19151_ (.A(_13106_), .B(_13111_), .Y(_13112_));
NAND_g _19152_ (.A(_12696_), .B(_12741_), .Y(_13113_));
NAND_g _19153_ (.A(_13112_), .B(_13113_), .Y(_13114_));
NAND_g _19154_ (.A(_13098_), .B(_13114_), .Y(_00432_));
NAND_g _19155_ (.A(reg_next_pc[27]), .B(_12549_), .Y(_13115_));
NAND_g _19156_ (.A(_13102_), .B(_13104_), .Y(_13116_));
XNOR_g _19157_ (.A(_11138_), .B(_12702_), .Y(_13117_));
XNOR_g _19158_ (.A(_13116_), .B(_13117_), .Y(_13118_));
NAND_g _19159_ (.A(instr_jal), .B(_13118_), .Y(_13119_));
AND_g _19160_ (.A(_12701_), .B(_13107_), .Y(_13120_));
AND_g _19161_ (.A(_12702_), .B(_13108_), .Y(_13121_));
NOR_g _19162_ (.A(_13120_), .B(_13121_), .Y(_13122_));
NAND_g _19163_ (.A(_10962_), .B(_13122_), .Y(_13123_));
AND_g _19164_ (.A(decoder_trigger), .B(_13123_), .Y(_13124_));
NAND_g _19165_ (.A(_13119_), .B(_13124_), .Y(_13125_));
NAND_g _19166_ (.A(_12702_), .B(_12741_), .Y(_13126_));
NAND_g _19167_ (.A(_13125_), .B(_13126_), .Y(_13127_));
NAND_g _19168_ (.A(_13115_), .B(_13127_), .Y(_00433_));
NAND_g _19169_ (.A(reg_next_pc[28]), .B(_12549_), .Y(_13128_));
AND_g _19170_ (.A(_12686_), .B(_12691_), .Y(_13129_));
AND_g _19171_ (.A(_12696_), .B(_12702_), .Y(_13130_));
NAND_g _19172_ (.A(_13129_), .B(_13130_), .Y(_13131_));
NAND_g _19173_ (.A(decoded_imm_j[31]), .B(_13131_), .Y(_13132_));
NOR_g _19174_ (.A(_13099_), .B(_13117_), .Y(_13133_));
NAND_g _19175_ (.A(_13103_), .B(_13133_), .Y(_13134_));
NAND_g _19176_ (.A(_13132_), .B(_13134_), .Y(_13135_));
NAND_g _19177_ (.A(decoded_imm_j[31]), .B(_12708_), .Y(_13136_));
XNOR_g _19178_ (.A(decoded_imm_j[31]), .B(_12707_), .Y(_13137_));
NAND_g _19179_ (.A(_13135_), .B(_13137_), .Y(_13138_));
XOR_g _19180_ (.A(_13135_), .B(_13137_), .Y(_13139_));
NAND_g _19181_ (.A(instr_jal), .B(_13139_), .Y(_13140_));
AND_g _19182_ (.A(_12708_), .B(_13120_), .Y(_13141_));
XNOR_g _19183_ (.A(_12707_), .B(_13120_), .Y(_13142_));
NAND_g _19184_ (.A(_10962_), .B(_13142_), .Y(_13143_));
AND_g _19185_ (.A(decoder_trigger), .B(_13143_), .Y(_13144_));
NAND_g _19186_ (.A(_13140_), .B(_13144_), .Y(_13145_));
NAND_g _19187_ (.A(_12707_), .B(_12741_), .Y(_13146_));
NAND_g _19188_ (.A(_13145_), .B(_13146_), .Y(_13147_));
NAND_g _19189_ (.A(_13128_), .B(_13147_), .Y(_00434_));
NAND_g _19190_ (.A(reg_next_pc[29]), .B(_12549_), .Y(_13148_));
NAND_g _19191_ (.A(_13136_), .B(_13138_), .Y(_13149_));
AND_g _19192_ (.A(decoded_imm_j[31]), .B(_12713_), .Y(_13150_));
XNOR_g _19193_ (.A(decoded_imm_j[31]), .B(_12713_), .Y(_13151_));
XNOR_g _19194_ (.A(_13149_), .B(_13151_), .Y(_13152_));
NAND_g _19195_ (.A(instr_jal), .B(_13152_), .Y(_13153_));
NAND_g _19196_ (.A(_12712_), .B(_13141_), .Y(_13154_));
NOR_g _19197_ (.A(_12713_), .B(_13141_), .Y(_13155_));
NOR_g _19198_ (.A(instr_jal), .B(_13155_), .Y(_13156_));
NAND_g _19199_ (.A(_13154_), .B(_13156_), .Y(_13157_));
AND_g _19200_ (.A(decoder_trigger), .B(_13157_), .Y(_13158_));
NAND_g _19201_ (.A(_13153_), .B(_13158_), .Y(_13159_));
NAND_g _19202_ (.A(_12714_), .B(_12741_), .Y(_13160_));
NAND_g _19203_ (.A(_13159_), .B(_13160_), .Y(_13161_));
NAND_g _19204_ (.A(_13148_), .B(_13161_), .Y(_00435_));
NAND_g _19205_ (.A(reg_next_pc[30]), .B(_12549_), .Y(_13162_));
NOR_g _19206_ (.A(_12719_), .B(_13154_), .Y(_13163_));
NOT_g _19207_ (.A(_13163_), .Y(_13164_));
NAND_g _19208_ (.A(_10962_), .B(_13164_), .Y(_13165_));
NAND_g _19209_ (.A(decoder_trigger), .B(_13165_), .Y(_13166_));
AND_g _19210_ (.A(decoder_trigger), .B(_12719_), .Y(_13167_));
NAND_g _19211_ (.A(_13154_), .B(_13167_), .Y(_13168_));
NAND_g _19212_ (.A(_13166_), .B(_13168_), .Y(_13169_));
AND_g _19213_ (.A(decoded_imm_j[31]), .B(_12719_), .Y(_13170_));
NOR_g _19214_ (.A(decoded_imm_j[31]), .B(_12719_), .Y(_13171_));
XNOR_g _19215_ (.A(decoded_imm_j[31]), .B(_12719_), .Y(_13172_));
NAND_g _19216_ (.A(_13136_), .B(_13151_), .Y(_13173_));
AND_g _19217_ (.A(_13149_), .B(_13173_), .Y(_13174_));
NOR_g _19218_ (.A(_13150_), .B(_13174_), .Y(_13175_));
XNOR_g _19219_ (.A(_13172_), .B(_13175_), .Y(_13176_));
NAND_g _19220_ (.A(instr_jal), .B(_13176_), .Y(_13177_));
NAND_g _19221_ (.A(_13169_), .B(_13177_), .Y(_13178_));
NAND_g _19222_ (.A(_12719_), .B(_12741_), .Y(_13179_));
NAND_g _19223_ (.A(_13178_), .B(_13179_), .Y(_13180_));
NAND_g _19224_ (.A(_13162_), .B(_13180_), .Y(_00436_));
NAND_g _19225_ (.A(_13170_), .B(_13175_), .Y(_13181_));
NAND_g _19226_ (.A(_13171_), .B(_13174_), .Y(_13182_));
AND_g _19227_ (.A(instr_jal), .B(_13182_), .Y(_13183_));
AND_g _19228_ (.A(_13181_), .B(_13183_), .Y(_13184_));
NOR_g _19229_ (.A(_13166_), .B(_13184_), .Y(_13185_));
NOR_g _19230_ (.A(_12724_), .B(_13185_), .Y(_13186_));
AND_g _19231_ (.A(reg_next_pc[31]), .B(_11263_), .Y(_13187_));
NOR_g _19232_ (.A(_13186_), .B(_13187_), .Y(_13188_));
AND_g _19233_ (.A(_12724_), .B(_13185_), .Y(_13189_));
NAND_g _19234_ (.A(_11262_), .B(_13189_), .Y(_13190_));
NAND_g _19235_ (.A(_13188_), .B(_13190_), .Y(_13191_));
AND_g _19236_ (.A(resetn), .B(_13191_), .Y(_00437_));
NOR_g _19237_ (.A(_10963_), .B(count_cycle[0]), .Y(_00438_));
NAND_g _19238_ (.A(count_cycle[0]), .B(count_cycle[1]), .Y(_13192_));
NOR_g _19239_ (.A(count_cycle[0]), .B(count_cycle[1]), .Y(_13193_));
NOR_g _19240_ (.A(_10963_), .B(_13193_), .Y(_13194_));
AND_g _19241_ (.A(_13192_), .B(_13194_), .Y(_00439_));
NOR_g _19242_ (.A(_11224_), .B(_13192_), .Y(_13195_));
NAND_g _19243_ (.A(_11224_), .B(_13192_), .Y(_13196_));
NAND_g _19244_ (.A(resetn), .B(_13196_), .Y(_13197_));
NOR_g _19245_ (.A(_13195_), .B(_13197_), .Y(_00440_));
NAND_g _19246_ (.A(count_cycle[3]), .B(_13195_), .Y(_13198_));
NOR_g _19247_ (.A(count_cycle[3]), .B(_13195_), .Y(_13199_));
NOR_g _19248_ (.A(_10963_), .B(_13199_), .Y(_13200_));
AND_g _19249_ (.A(_13198_), .B(_13200_), .Y(_00441_));
NOR_g _19250_ (.A(_11225_), .B(_13198_), .Y(_13201_));
NAND_g _19251_ (.A(_11225_), .B(_13198_), .Y(_13202_));
NAND_g _19252_ (.A(resetn), .B(_13202_), .Y(_13203_));
NOR_g _19253_ (.A(_13201_), .B(_13203_), .Y(_00442_));
NAND_g _19254_ (.A(count_cycle[5]), .B(_13201_), .Y(_13204_));
NOR_g _19255_ (.A(count_cycle[5]), .B(_13201_), .Y(_13205_));
NOR_g _19256_ (.A(_10963_), .B(_13205_), .Y(_13206_));
AND_g _19257_ (.A(_13204_), .B(_13206_), .Y(_00443_));
NOR_g _19258_ (.A(_11226_), .B(_13204_), .Y(_13207_));
NAND_g _19259_ (.A(_11226_), .B(_13204_), .Y(_13208_));
NAND_g _19260_ (.A(resetn), .B(_13208_), .Y(_13209_));
NOR_g _19261_ (.A(_13207_), .B(_13209_), .Y(_00444_));
NAND_g _19262_ (.A(count_cycle[7]), .B(_13207_), .Y(_13210_));
NOR_g _19263_ (.A(count_cycle[7]), .B(_13207_), .Y(_13211_));
NOR_g _19264_ (.A(_10963_), .B(_13211_), .Y(_13212_));
AND_g _19265_ (.A(_13210_), .B(_13212_), .Y(_00445_));
NOR_g _19266_ (.A(_11227_), .B(_13210_), .Y(_13213_));
NAND_g _19267_ (.A(_11227_), .B(_13210_), .Y(_13214_));
NAND_g _19268_ (.A(resetn), .B(_13214_), .Y(_13215_));
NOR_g _19269_ (.A(_13213_), .B(_13215_), .Y(_00446_));
NAND_g _19270_ (.A(count_cycle[9]), .B(_13213_), .Y(_13216_));
NOR_g _19271_ (.A(count_cycle[9]), .B(_13213_), .Y(_13217_));
NOR_g _19272_ (.A(_10963_), .B(_13217_), .Y(_13218_));
AND_g _19273_ (.A(_13216_), .B(_13218_), .Y(_00447_));
NOR_g _19274_ (.A(_11228_), .B(_13216_), .Y(_13219_));
NAND_g _19275_ (.A(_11228_), .B(_13216_), .Y(_13220_));
NAND_g _19276_ (.A(resetn), .B(_13220_), .Y(_13221_));
NOR_g _19277_ (.A(_13219_), .B(_13221_), .Y(_00448_));
NAND_g _19278_ (.A(count_cycle[11]), .B(_13219_), .Y(_13222_));
NOR_g _19279_ (.A(count_cycle[11]), .B(_13219_), .Y(_13223_));
NOR_g _19280_ (.A(_10963_), .B(_13223_), .Y(_13224_));
AND_g _19281_ (.A(_13222_), .B(_13224_), .Y(_00449_));
NOR_g _19282_ (.A(_11229_), .B(_13222_), .Y(_13225_));
NAND_g _19283_ (.A(_11229_), .B(_13222_), .Y(_13226_));
NAND_g _19284_ (.A(resetn), .B(_13226_), .Y(_13227_));
NOR_g _19285_ (.A(_13225_), .B(_13227_), .Y(_00450_));
NAND_g _19286_ (.A(count_cycle[13]), .B(_13225_), .Y(_13228_));
NOR_g _19287_ (.A(count_cycle[13]), .B(_13225_), .Y(_13229_));
NOR_g _19288_ (.A(_10963_), .B(_13229_), .Y(_13230_));
AND_g _19289_ (.A(_13228_), .B(_13230_), .Y(_00451_));
NOR_g _19290_ (.A(_11230_), .B(_13228_), .Y(_13231_));
NAND_g _19291_ (.A(_11230_), .B(_13228_), .Y(_13232_));
NAND_g _19292_ (.A(resetn), .B(_13232_), .Y(_13233_));
NOR_g _19293_ (.A(_13231_), .B(_13233_), .Y(_00452_));
NAND_g _19294_ (.A(count_cycle[15]), .B(_13231_), .Y(_13234_));
NOR_g _19295_ (.A(count_cycle[15]), .B(_13231_), .Y(_13235_));
NOR_g _19296_ (.A(_10963_), .B(_13235_), .Y(_13236_));
AND_g _19297_ (.A(_13234_), .B(_13236_), .Y(_00453_));
NOR_g _19298_ (.A(_11231_), .B(_13234_), .Y(_13237_));
NAND_g _19299_ (.A(_11231_), .B(_13234_), .Y(_13238_));
NAND_g _19300_ (.A(resetn), .B(_13238_), .Y(_13239_));
NOR_g _19301_ (.A(_13237_), .B(_13239_), .Y(_00454_));
NAND_g _19302_ (.A(count_cycle[17]), .B(_13237_), .Y(_13240_));
NOR_g _19303_ (.A(count_cycle[17]), .B(_13237_), .Y(_13241_));
NOR_g _19304_ (.A(_10963_), .B(_13241_), .Y(_13242_));
AND_g _19305_ (.A(_13240_), .B(_13242_), .Y(_00455_));
NOR_g _19306_ (.A(_11232_), .B(_13240_), .Y(_13243_));
NAND_g _19307_ (.A(_11232_), .B(_13240_), .Y(_13244_));
NAND_g _19308_ (.A(resetn), .B(_13244_), .Y(_13245_));
NOR_g _19309_ (.A(_13243_), .B(_13245_), .Y(_00456_));
NAND_g _19310_ (.A(count_cycle[19]), .B(_13243_), .Y(_13246_));
NOR_g _19311_ (.A(count_cycle[19]), .B(_13243_), .Y(_13247_));
NOR_g _19312_ (.A(_10963_), .B(_13247_), .Y(_13248_));
AND_g _19313_ (.A(_13246_), .B(_13248_), .Y(_00457_));
NOR_g _19314_ (.A(_11233_), .B(_13246_), .Y(_13249_));
NAND_g _19315_ (.A(_11233_), .B(_13246_), .Y(_13250_));
NAND_g _19316_ (.A(resetn), .B(_13250_), .Y(_13251_));
NOR_g _19317_ (.A(_13249_), .B(_13251_), .Y(_00458_));
NAND_g _19318_ (.A(count_cycle[21]), .B(_13249_), .Y(_13252_));
NOR_g _19319_ (.A(count_cycle[21]), .B(_13249_), .Y(_13253_));
NOR_g _19320_ (.A(_10963_), .B(_13253_), .Y(_13254_));
AND_g _19321_ (.A(_13252_), .B(_13254_), .Y(_00459_));
NOR_g _19322_ (.A(_11234_), .B(_13252_), .Y(_13255_));
NAND_g _19323_ (.A(_11234_), .B(_13252_), .Y(_13256_));
NAND_g _19324_ (.A(resetn), .B(_13256_), .Y(_13257_));
NOR_g _19325_ (.A(_13255_), .B(_13257_), .Y(_00460_));
NAND_g _19326_ (.A(count_cycle[23]), .B(_13255_), .Y(_13258_));
NOR_g _19327_ (.A(count_cycle[23]), .B(_13255_), .Y(_13259_));
NOR_g _19328_ (.A(_10963_), .B(_13259_), .Y(_13260_));
AND_g _19329_ (.A(_13258_), .B(_13260_), .Y(_00461_));
NOR_g _19330_ (.A(_11235_), .B(_13258_), .Y(_13261_));
NAND_g _19331_ (.A(_11235_), .B(_13258_), .Y(_13262_));
NAND_g _19332_ (.A(resetn), .B(_13262_), .Y(_13263_));
NOR_g _19333_ (.A(_13261_), .B(_13263_), .Y(_00462_));
NAND_g _19334_ (.A(count_cycle[25]), .B(_13261_), .Y(_13264_));
NOR_g _19335_ (.A(count_cycle[25]), .B(_13261_), .Y(_13265_));
NOR_g _19336_ (.A(_10963_), .B(_13265_), .Y(_13266_));
AND_g _19337_ (.A(_13264_), .B(_13266_), .Y(_00463_));
NOR_g _19338_ (.A(_11236_), .B(_13264_), .Y(_13267_));
NAND_g _19339_ (.A(_11236_), .B(_13264_), .Y(_13268_));
NAND_g _19340_ (.A(resetn), .B(_13268_), .Y(_13269_));
NOR_g _19341_ (.A(_13267_), .B(_13269_), .Y(_00464_));
NAND_g _19342_ (.A(count_cycle[27]), .B(_13267_), .Y(_13270_));
NOR_g _19343_ (.A(count_cycle[27]), .B(_13267_), .Y(_13271_));
NOR_g _19344_ (.A(_10963_), .B(_13271_), .Y(_13272_));
AND_g _19345_ (.A(_13270_), .B(_13272_), .Y(_00465_));
NOR_g _19346_ (.A(_11237_), .B(_13270_), .Y(_13273_));
NAND_g _19347_ (.A(_11237_), .B(_13270_), .Y(_13274_));
NAND_g _19348_ (.A(resetn), .B(_13274_), .Y(_13275_));
NOR_g _19349_ (.A(_13273_), .B(_13275_), .Y(_00466_));
NAND_g _19350_ (.A(count_cycle[29]), .B(_13273_), .Y(_13276_));
NOR_g _19351_ (.A(count_cycle[29]), .B(_13273_), .Y(_13277_));
NOR_g _19352_ (.A(_10963_), .B(_13277_), .Y(_13278_));
AND_g _19353_ (.A(_13276_), .B(_13278_), .Y(_00467_));
NOR_g _19354_ (.A(_11238_), .B(_13276_), .Y(_13279_));
NAND_g _19355_ (.A(_11238_), .B(_13276_), .Y(_13280_));
NAND_g _19356_ (.A(resetn), .B(_13280_), .Y(_13281_));
NOR_g _19357_ (.A(_13279_), .B(_13281_), .Y(_00468_));
NAND_g _19358_ (.A(count_cycle[31]), .B(_13279_), .Y(_13282_));
NOR_g _19359_ (.A(count_cycle[31]), .B(_13279_), .Y(_13283_));
NOR_g _19360_ (.A(_10963_), .B(_13283_), .Y(_13284_));
AND_g _19361_ (.A(_13282_), .B(_13284_), .Y(_00469_));
NOR_g _19362_ (.A(_11239_), .B(_13282_), .Y(_13285_));
NAND_g _19363_ (.A(_11239_), .B(_13282_), .Y(_13286_));
NAND_g _19364_ (.A(resetn), .B(_13286_), .Y(_13287_));
NOR_g _19365_ (.A(_13285_), .B(_13287_), .Y(_00470_));
NAND_g _19366_ (.A(count_cycle[33]), .B(_13285_), .Y(_13288_));
NOR_g _19367_ (.A(count_cycle[33]), .B(_13285_), .Y(_13289_));
NOR_g _19368_ (.A(_10963_), .B(_13289_), .Y(_13290_));
AND_g _19369_ (.A(_13288_), .B(_13290_), .Y(_00471_));
NOR_g _19370_ (.A(_11240_), .B(_13288_), .Y(_13291_));
NAND_g _19371_ (.A(_11240_), .B(_13288_), .Y(_13292_));
NAND_g _19372_ (.A(resetn), .B(_13292_), .Y(_13293_));
NOR_g _19373_ (.A(_13291_), .B(_13293_), .Y(_00472_));
NAND_g _19374_ (.A(count_cycle[35]), .B(_13291_), .Y(_13294_));
NOR_g _19375_ (.A(count_cycle[35]), .B(_13291_), .Y(_13295_));
NOR_g _19376_ (.A(_10963_), .B(_13295_), .Y(_13296_));
AND_g _19377_ (.A(_13294_), .B(_13296_), .Y(_00473_));
NOR_g _19378_ (.A(_11241_), .B(_13294_), .Y(_13297_));
NAND_g _19379_ (.A(_11241_), .B(_13294_), .Y(_13298_));
NAND_g _19380_ (.A(resetn), .B(_13298_), .Y(_13299_));
NOR_g _19381_ (.A(_13297_), .B(_13299_), .Y(_00474_));
NAND_g _19382_ (.A(count_cycle[37]), .B(_13297_), .Y(_13300_));
NOR_g _19383_ (.A(count_cycle[37]), .B(_13297_), .Y(_13301_));
NOR_g _19384_ (.A(_10963_), .B(_13301_), .Y(_13302_));
AND_g _19385_ (.A(_13300_), .B(_13302_), .Y(_00475_));
NOR_g _19386_ (.A(_11242_), .B(_13300_), .Y(_13303_));
NAND_g _19387_ (.A(_11242_), .B(_13300_), .Y(_13304_));
NAND_g _19388_ (.A(resetn), .B(_13304_), .Y(_13305_));
NOR_g _19389_ (.A(_13303_), .B(_13305_), .Y(_00476_));
NAND_g _19390_ (.A(count_cycle[39]), .B(_13303_), .Y(_13306_));
NOR_g _19391_ (.A(count_cycle[39]), .B(_13303_), .Y(_13307_));
NOR_g _19392_ (.A(_10963_), .B(_13307_), .Y(_13308_));
AND_g _19393_ (.A(_13306_), .B(_13308_), .Y(_00477_));
NOR_g _19394_ (.A(_11243_), .B(_13306_), .Y(_13309_));
NAND_g _19395_ (.A(_11243_), .B(_13306_), .Y(_13310_));
NAND_g _19396_ (.A(resetn), .B(_13310_), .Y(_13311_));
NOR_g _19397_ (.A(_13309_), .B(_13311_), .Y(_00478_));
NAND_g _19398_ (.A(count_cycle[41]), .B(_13309_), .Y(_13312_));
NOR_g _19399_ (.A(count_cycle[41]), .B(_13309_), .Y(_13313_));
NOR_g _19400_ (.A(_10963_), .B(_13313_), .Y(_13314_));
AND_g _19401_ (.A(_13312_), .B(_13314_), .Y(_00479_));
NOR_g _19402_ (.A(_11244_), .B(_13312_), .Y(_13315_));
NAND_g _19403_ (.A(_11244_), .B(_13312_), .Y(_13316_));
NAND_g _19404_ (.A(resetn), .B(_13316_), .Y(_13317_));
NOR_g _19405_ (.A(_13315_), .B(_13317_), .Y(_00480_));
NAND_g _19406_ (.A(count_cycle[43]), .B(_13315_), .Y(_13318_));
NOR_g _19407_ (.A(count_cycle[43]), .B(_13315_), .Y(_13319_));
NOR_g _19408_ (.A(_10963_), .B(_13319_), .Y(_13320_));
AND_g _19409_ (.A(_13318_), .B(_13320_), .Y(_00481_));
NOR_g _19410_ (.A(_11245_), .B(_13318_), .Y(_13321_));
NAND_g _19411_ (.A(_11245_), .B(_13318_), .Y(_13322_));
NAND_g _19412_ (.A(resetn), .B(_13322_), .Y(_13323_));
NOR_g _19413_ (.A(_13321_), .B(_13323_), .Y(_00482_));
NAND_g _19414_ (.A(count_cycle[45]), .B(_13321_), .Y(_13324_));
NOR_g _19415_ (.A(count_cycle[45]), .B(_13321_), .Y(_13325_));
NOR_g _19416_ (.A(_10963_), .B(_13325_), .Y(_13326_));
AND_g _19417_ (.A(_13324_), .B(_13326_), .Y(_00483_));
NOR_g _19418_ (.A(_11246_), .B(_13324_), .Y(_13327_));
NAND_g _19419_ (.A(_11246_), .B(_13324_), .Y(_13328_));
NAND_g _19420_ (.A(resetn), .B(_13328_), .Y(_13329_));
NOR_g _19421_ (.A(_13327_), .B(_13329_), .Y(_00484_));
NAND_g _19422_ (.A(count_cycle[47]), .B(_13327_), .Y(_13330_));
NOR_g _19423_ (.A(count_cycle[47]), .B(_13327_), .Y(_13331_));
NOR_g _19424_ (.A(_10963_), .B(_13331_), .Y(_13332_));
AND_g _19425_ (.A(_13330_), .B(_13332_), .Y(_00485_));
NOR_g _19426_ (.A(_11247_), .B(_13330_), .Y(_13333_));
NAND_g _19427_ (.A(_11247_), .B(_13330_), .Y(_13334_));
NAND_g _19428_ (.A(resetn), .B(_13334_), .Y(_13335_));
NOR_g _19429_ (.A(_13333_), .B(_13335_), .Y(_00486_));
NAND_g _19430_ (.A(count_cycle[49]), .B(_13333_), .Y(_13336_));
NOR_g _19431_ (.A(count_cycle[49]), .B(_13333_), .Y(_13337_));
NOR_g _19432_ (.A(_10963_), .B(_13337_), .Y(_13338_));
AND_g _19433_ (.A(_13336_), .B(_13338_), .Y(_00487_));
NOR_g _19434_ (.A(_11248_), .B(_13336_), .Y(_13339_));
NAND_g _19435_ (.A(_11248_), .B(_13336_), .Y(_13340_));
NAND_g _19436_ (.A(resetn), .B(_13340_), .Y(_13341_));
NOR_g _19437_ (.A(_13339_), .B(_13341_), .Y(_00488_));
NAND_g _19438_ (.A(count_cycle[51]), .B(_13339_), .Y(_13342_));
NOR_g _19439_ (.A(count_cycle[51]), .B(_13339_), .Y(_13343_));
NOR_g _19440_ (.A(_10963_), .B(_13343_), .Y(_13344_));
AND_g _19441_ (.A(_13342_), .B(_13344_), .Y(_00489_));
NOR_g _19442_ (.A(_11249_), .B(_13342_), .Y(_13345_));
NAND_g _19443_ (.A(_11249_), .B(_13342_), .Y(_13346_));
NAND_g _19444_ (.A(resetn), .B(_13346_), .Y(_13347_));
NOR_g _19445_ (.A(_13345_), .B(_13347_), .Y(_00490_));
NAND_g _19446_ (.A(count_cycle[53]), .B(_13345_), .Y(_13348_));
NOR_g _19447_ (.A(count_cycle[53]), .B(_13345_), .Y(_13349_));
NOR_g _19448_ (.A(_10963_), .B(_13349_), .Y(_13350_));
AND_g _19449_ (.A(_13348_), .B(_13350_), .Y(_00491_));
NOR_g _19450_ (.A(_11250_), .B(_13348_), .Y(_13351_));
NAND_g _19451_ (.A(_11250_), .B(_13348_), .Y(_13352_));
NAND_g _19452_ (.A(resetn), .B(_13352_), .Y(_13353_));
NOR_g _19453_ (.A(_13351_), .B(_13353_), .Y(_00492_));
NAND_g _19454_ (.A(count_cycle[55]), .B(_13351_), .Y(_13354_));
NOR_g _19455_ (.A(count_cycle[55]), .B(_13351_), .Y(_13355_));
NOR_g _19456_ (.A(_10963_), .B(_13355_), .Y(_13356_));
AND_g _19457_ (.A(_13354_), .B(_13356_), .Y(_00493_));
NOR_g _19458_ (.A(_11251_), .B(_13354_), .Y(_13357_));
NAND_g _19459_ (.A(_11251_), .B(_13354_), .Y(_13358_));
NAND_g _19460_ (.A(resetn), .B(_13358_), .Y(_13359_));
NOR_g _19461_ (.A(_13357_), .B(_13359_), .Y(_00494_));
NAND_g _19462_ (.A(count_cycle[57]), .B(_13357_), .Y(_13360_));
NOR_g _19463_ (.A(count_cycle[57]), .B(_13357_), .Y(_13361_));
NOR_g _19464_ (.A(_10963_), .B(_13361_), .Y(_13362_));
AND_g _19465_ (.A(_13360_), .B(_13362_), .Y(_00495_));
NOR_g _19466_ (.A(_11252_), .B(_13360_), .Y(_13363_));
NAND_g _19467_ (.A(_11252_), .B(_13360_), .Y(_13364_));
NAND_g _19468_ (.A(resetn), .B(_13364_), .Y(_13365_));
NOR_g _19469_ (.A(_13363_), .B(_13365_), .Y(_00496_));
NAND_g _19470_ (.A(count_cycle[59]), .B(_13363_), .Y(_13366_));
NOR_g _19471_ (.A(count_cycle[59]), .B(_13363_), .Y(_13367_));
NOR_g _19472_ (.A(_10963_), .B(_13367_), .Y(_13368_));
AND_g _19473_ (.A(_13366_), .B(_13368_), .Y(_00497_));
NOR_g _19474_ (.A(_11253_), .B(_13366_), .Y(_13369_));
NAND_g _19475_ (.A(_11253_), .B(_13366_), .Y(_13370_));
NAND_g _19476_ (.A(resetn), .B(_13370_), .Y(_13371_));
NOR_g _19477_ (.A(_13369_), .B(_13371_), .Y(_00498_));
NAND_g _19478_ (.A(count_cycle[61]), .B(_13369_), .Y(_13372_));
NOT_g _19479_ (.A(_13372_), .Y(_13373_));
NOR_g _19480_ (.A(count_cycle[61]), .B(_13369_), .Y(_13374_));
NOR_g _19481_ (.A(_10963_), .B(_13374_), .Y(_13375_));
AND_g _19482_ (.A(_13372_), .B(_13375_), .Y(_00499_));
NAND_g _19483_ (.A(count_cycle[62]), .B(_13373_), .Y(_13376_));
NAND_g _19484_ (.A(_11254_), .B(_13372_), .Y(_13377_));
AND_g _19485_ (.A(resetn), .B(_13377_), .Y(_13378_));
AND_g _19486_ (.A(_13376_), .B(_13378_), .Y(_00500_));
XNOR_g _19487_ (.A(count_cycle[63]), .B(_13376_), .Y(_13379_));
AND_g _19488_ (.A(resetn), .B(_13379_), .Y(_00501_));
NAND_g _19489_ (.A(_10905_), .B(_10971_), .Y(_13380_));
NOR_g _19490_ (.A(reg_sh[2]), .B(reg_sh[3]), .Y(_13381_));
AND_g _19491_ (.A(_11208_), .B(_13381_), .Y(_13382_));
NAND_g _19492_ (.A(_11208_), .B(_13381_), .Y(_13383_));
NAND_g _19493_ (.A(_11207_), .B(_13382_), .Y(_13384_));
NOR_g _19494_ (.A(reg_sh[1]), .B(_13384_), .Y(_13385_));
AND_g _19495_ (.A(cpu_state[2]), .B(_11257_), .Y(_13386_));
AND_g _19496_ (.A(_11268_), .B(_13386_), .Y(_13387_));
NAND_g _19497_ (.A(_11268_), .B(_13386_), .Y(_13388_));
NOR_g _19498_ (.A(_13385_), .B(_13388_), .Y(_13389_));
NOT_g _19499_ (.A(_13389_), .Y(_13390_));
NAND_g _19500_ (.A(_13380_), .B(_13389_), .Y(_13391_));
AND_g _19501_ (.A(_11206_), .B(_11256_), .Y(_13392_));
AND_g _19502_ (.A(cpu_state[1]), .B(_13392_), .Y(_13393_));
NAND_g _19503_ (.A(_11268_), .B(_13393_), .Y(_13394_));
NOT_g _19504_ (.A(_13394_), .Y(_13395_));
AND_g _19505_ (.A(mem_do_prefetch), .B(_11916_), .Y(_13396_));
NOR_g _19506_ (.A(mem_do_wdata), .B(_13396_), .Y(_13397_));
NOR_g _19507_ (.A(_13394_), .B(_13397_), .Y(_13398_));
NOT_g _19508_ (.A(_13398_), .Y(_13399_));
NAND_g _19509_ (.A(resetn), .B(_13399_), .Y(_13400_));
NAND_g _19510_ (.A(cpu_state[0]), .B(_11256_), .Y(_13401_));
NOR_g _19511_ (.A(cpu_state[1]), .B(_13401_), .Y(_13402_));
NAND_g _19512_ (.A(_11268_), .B(_13402_), .Y(_13403_));
NOT_g _19513_ (.A(_13403_), .Y(dbg_ascii_state[35]));
NOR_g _19514_ (.A(mem_do_rdata), .B(_13396_), .Y(_13404_));
NOR_g _19515_ (.A(_13403_), .B(_13404_), .Y(_13405_));
NOR_g _19516_ (.A(_13400_), .B(_13405_), .Y(_13406_));
AND_g _19517_ (.A(_11204_), .B(_11267_), .Y(_13407_));
AND_g _19518_ (.A(cpu_state[5]), .B(_13407_), .Y(_13408_));
AND_g _19519_ (.A(_11258_), .B(_13408_), .Y(_13409_));
NAND_g _19520_ (.A(_11258_), .B(_13408_), .Y(_13410_));
AND_g _19521_ (.A(_13388_), .B(_13394_), .Y(_13411_));
NOT_g _19522_ (.A(_13411_), .Y(dbg_ascii_state[36]));
AND_g _19523_ (.A(_13403_), .B(_13411_), .Y(_13412_));
NOT_g _19524_ (.A(_13412_), .Y(dbg_ascii_state[16]));
AND_g _19525_ (.A(_13394_), .B(_13403_), .Y(_13413_));
NAND_g _19526_ (.A(_13394_), .B(_13403_), .Y(_13414_));
NAND_g _19527_ (.A(_13410_), .B(_13412_), .Y(_13415_));
AND_g _19528_ (.A(_13385_), .B(_13387_), .Y(_13416_));
NOR_g _19529_ (.A(instr_srli), .B(instr_srai), .Y(_13417_));
NOR_g _19530_ (.A(instr_sra), .B(instr_srl), .Y(_13418_));
NAND_g _19531_ (.A(_13417_), .B(_13418_), .Y(_13419_));
NAND_g _19532_ (.A(_10909_), .B(_10969_), .Y(_13420_));
NOR_g _19533_ (.A(_13419_), .B(_13420_), .Y(_13421_));
AND_g _19534_ (.A(_13387_), .B(_13421_), .Y(_13422_));
NOR_g _19535_ (.A(_13416_), .B(_13422_), .Y(_13423_));
AND_g _19536_ (.A(_13415_), .B(_13423_), .Y(_13424_));
AND_g _19537_ (.A(_13406_), .B(_13424_), .Y(_13425_));
AND_g _19538_ (.A(_13391_), .B(_13425_), .Y(_13426_));
NOR_g _19539_ (.A(pcpi_rs1[31]), .B(_13426_), .Y(_13427_));
AND_g _19540_ (.A(dbg_ascii_state[35]), .B(_13404_), .Y(_13428_));
NAND_g _19541_ (.A(dbg_ascii_state[35]), .B(_13404_), .Y(_13429_));
AND_g _19542_ (.A(_13395_), .B(_13397_), .Y(_13430_));
NOT_g _19543_ (.A(_13430_), .Y(_13431_));
NAND_g _19544_ (.A(_13429_), .B(_13431_), .Y(_13432_));
NAND_g _19545_ (.A(decoded_imm[30]), .B(pcpi_rs1[30]), .Y(_13433_));
XOR_g _19546_ (.A(decoded_imm[30]), .B(pcpi_rs1[30]), .Y(_13434_));
NAND_g _19547_ (.A(decoded_imm[29]), .B(pcpi_rs1[29]), .Y(_13435_));
NOR_g _19548_ (.A(decoded_imm[29]), .B(pcpi_rs1[29]), .Y(_13436_));
NAND_g _19549_ (.A(decoded_imm[28]), .B(pcpi_rs1[28]), .Y(_13437_));
XOR_g _19550_ (.A(decoded_imm[28]), .B(pcpi_rs1[28]), .Y(_13438_));
NAND_g _19551_ (.A(decoded_imm[27]), .B(pcpi_rs1[27]), .Y(_13439_));
NOR_g _19552_ (.A(decoded_imm[27]), .B(pcpi_rs1[27]), .Y(_13440_));
NAND_g _19553_ (.A(decoded_imm[26]), .B(pcpi_rs1[26]), .Y(_13441_));
XOR_g _19554_ (.A(decoded_imm[26]), .B(pcpi_rs1[26]), .Y(_13442_));
NAND_g _19555_ (.A(decoded_imm[25]), .B(pcpi_rs1[25]), .Y(_13443_));
NAND_g _19556_ (.A(decoded_imm[24]), .B(pcpi_rs1[24]), .Y(_13444_));
XOR_g _19557_ (.A(decoded_imm[24]), .B(pcpi_rs1[24]), .Y(_13445_));
NOR_g _19558_ (.A(decoded_imm[23]), .B(pcpi_rs1[23]), .Y(_13446_));
NAND_g _19559_ (.A(decoded_imm[23]), .B(pcpi_rs1[23]), .Y(_13447_));
NAND_g _19560_ (.A(decoded_imm[22]), .B(pcpi_rs1[22]), .Y(_13448_));
XOR_g _19561_ (.A(decoded_imm[22]), .B(pcpi_rs1[22]), .Y(_13449_));
NAND_g _19562_ (.A(decoded_imm[21]), .B(pcpi_rs1[21]), .Y(_13450_));
NOR_g _19563_ (.A(decoded_imm[21]), .B(pcpi_rs1[21]), .Y(_13451_));
NAND_g _19564_ (.A(decoded_imm[20]), .B(pcpi_rs1[20]), .Y(_13452_));
XOR_g _19565_ (.A(decoded_imm[20]), .B(pcpi_rs1[20]), .Y(_13453_));
NOR_g _19566_ (.A(decoded_imm[19]), .B(pcpi_rs1[19]), .Y(_13454_));
NAND_g _19567_ (.A(decoded_imm[19]), .B(pcpi_rs1[19]), .Y(_13455_));
NAND_g _19568_ (.A(decoded_imm[18]), .B(pcpi_rs1[18]), .Y(_13456_));
XOR_g _19569_ (.A(decoded_imm[18]), .B(pcpi_rs1[18]), .Y(_13457_));
NAND_g _19570_ (.A(decoded_imm[17]), .B(pcpi_rs1[17]), .Y(_13458_));
NOR_g _19571_ (.A(decoded_imm[17]), .B(pcpi_rs1[17]), .Y(_13459_));
NAND_g _19572_ (.A(decoded_imm[16]), .B(pcpi_rs1[16]), .Y(_13460_));
XOR_g _19573_ (.A(decoded_imm[16]), .B(pcpi_rs1[16]), .Y(_13461_));
NOR_g _19574_ (.A(decoded_imm[15]), .B(pcpi_rs1[15]), .Y(_13462_));
NAND_g _19575_ (.A(decoded_imm[15]), .B(pcpi_rs1[15]), .Y(_13463_));
NAND_g _19576_ (.A(decoded_imm[14]), .B(pcpi_rs1[14]), .Y(_13464_));
XOR_g _19577_ (.A(decoded_imm[14]), .B(pcpi_rs1[14]), .Y(_13465_));
NAND_g _19578_ (.A(decoded_imm[13]), .B(pcpi_rs1[13]), .Y(_13466_));
NOR_g _19579_ (.A(decoded_imm[13]), .B(pcpi_rs1[13]), .Y(_13467_));
NAND_g _19580_ (.A(decoded_imm[12]), .B(pcpi_rs1[12]), .Y(_13468_));
XOR_g _19581_ (.A(decoded_imm[12]), .B(pcpi_rs1[12]), .Y(_13469_));
NAND_g _19582_ (.A(decoded_imm[11]), .B(pcpi_rs1[11]), .Y(_13470_));
NOR_g _19583_ (.A(decoded_imm[11]), .B(pcpi_rs1[11]), .Y(_13471_));
NAND_g _19584_ (.A(decoded_imm[10]), .B(pcpi_rs1[10]), .Y(_13472_));
XOR_g _19585_ (.A(decoded_imm[10]), .B(pcpi_rs1[10]), .Y(_13473_));
NAND_g _19586_ (.A(decoded_imm[9]), .B(pcpi_rs1[9]), .Y(_13474_));
NOR_g _19587_ (.A(decoded_imm[9]), .B(pcpi_rs1[9]), .Y(_13475_));
NAND_g _19588_ (.A(decoded_imm[8]), .B(pcpi_rs1[8]), .Y(_13476_));
XOR_g _19589_ (.A(decoded_imm[8]), .B(pcpi_rs1[8]), .Y(_13477_));
NAND_g _19590_ (.A(decoded_imm[7]), .B(pcpi_rs1[7]), .Y(_13478_));
NOR_g _19591_ (.A(decoded_imm[7]), .B(pcpi_rs1[7]), .Y(_13479_));
NAND_g _19592_ (.A(decoded_imm[6]), .B(pcpi_rs1[6]), .Y(_13480_));
XOR_g _19593_ (.A(decoded_imm[6]), .B(pcpi_rs1[6]), .Y(_13481_));
NAND_g _19594_ (.A(decoded_imm[5]), .B(pcpi_rs1[5]), .Y(_13482_));
NAND_g _19595_ (.A(decoded_imm[4]), .B(pcpi_rs1[4]), .Y(_13483_));
XOR_g _19596_ (.A(decoded_imm[4]), .B(pcpi_rs1[4]), .Y(_13484_));
NAND_g _19597_ (.A(decoded_imm[3]), .B(pcpi_rs1[3]), .Y(_13485_));
NOR_g _19598_ (.A(decoded_imm[3]), .B(pcpi_rs1[3]), .Y(_13486_));
NAND_g _19599_ (.A(decoded_imm[2]), .B(pcpi_rs1[2]), .Y(_13487_));
NAND_g _19600_ (.A(decoded_imm[1]), .B(pcpi_rs1[1]), .Y(_13488_));
AND_g _19601_ (.A(decoded_imm[0]), .B(pcpi_rs1[0]), .Y(_13489_));
XOR_g _19602_ (.A(decoded_imm[1]), .B(pcpi_rs1[1]), .Y(_13490_));
NAND_g _19603_ (.A(_13489_), .B(_13490_), .Y(_13491_));
NAND_g _19604_ (.A(_13488_), .B(_13491_), .Y(_13492_));
XOR_g _19605_ (.A(decoded_imm[2]), .B(pcpi_rs1[2]), .Y(_13493_));
NAND_g _19606_ (.A(_13492_), .B(_13493_), .Y(_13494_));
AND_g _19607_ (.A(_13487_), .B(_13494_), .Y(_13495_));
AND_g _19608_ (.A(_13485_), .B(_13495_), .Y(_13496_));
NOR_g _19609_ (.A(_13486_), .B(_13496_), .Y(_13497_));
NAND_g _19610_ (.A(_13484_), .B(_13497_), .Y(_13498_));
NAND_g _19611_ (.A(_13483_), .B(_13498_), .Y(_13499_));
XOR_g _19612_ (.A(decoded_imm[5]), .B(pcpi_rs1[5]), .Y(_13500_));
NAND_g _19613_ (.A(_13499_), .B(_13500_), .Y(_13501_));
NAND_g _19614_ (.A(_13482_), .B(_13501_), .Y(_13502_));
NAND_g _19615_ (.A(_13481_), .B(_13502_), .Y(_13503_));
AND_g _19616_ (.A(_13480_), .B(_13503_), .Y(_13504_));
AND_g _19617_ (.A(_13478_), .B(_13504_), .Y(_13505_));
NOR_g _19618_ (.A(_13479_), .B(_13505_), .Y(_13506_));
NAND_g _19619_ (.A(_13477_), .B(_13506_), .Y(_13507_));
AND_g _19620_ (.A(_13476_), .B(_13507_), .Y(_13508_));
AND_g _19621_ (.A(_13474_), .B(_13508_), .Y(_13509_));
NOR_g _19622_ (.A(_13475_), .B(_13509_), .Y(_13510_));
NAND_g _19623_ (.A(_13473_), .B(_13510_), .Y(_13511_));
AND_g _19624_ (.A(_13472_), .B(_13511_), .Y(_13512_));
AND_g _19625_ (.A(_13470_), .B(_13512_), .Y(_13513_));
NOR_g _19626_ (.A(_13471_), .B(_13513_), .Y(_13514_));
NAND_g _19627_ (.A(_13469_), .B(_13514_), .Y(_13515_));
AND_g _19628_ (.A(_13468_), .B(_13515_), .Y(_13516_));
AND_g _19629_ (.A(_13466_), .B(_13516_), .Y(_13517_));
NOR_g _19630_ (.A(_13467_), .B(_13517_), .Y(_13518_));
NAND_g _19631_ (.A(_13465_), .B(_13518_), .Y(_13519_));
AND_g _19632_ (.A(_13464_), .B(_13519_), .Y(_13520_));
AND_g _19633_ (.A(_13463_), .B(_13520_), .Y(_13521_));
NOR_g _19634_ (.A(_13462_), .B(_13521_), .Y(_13522_));
NAND_g _19635_ (.A(_13461_), .B(_13522_), .Y(_13523_));
AND_g _19636_ (.A(_13460_), .B(_13523_), .Y(_13524_));
AND_g _19637_ (.A(_13458_), .B(_13524_), .Y(_13525_));
NOR_g _19638_ (.A(_13459_), .B(_13525_), .Y(_13526_));
NAND_g _19639_ (.A(_13457_), .B(_13526_), .Y(_13527_));
AND_g _19640_ (.A(_13456_), .B(_13527_), .Y(_13528_));
AND_g _19641_ (.A(_13455_), .B(_13528_), .Y(_13529_));
NOR_g _19642_ (.A(_13454_), .B(_13529_), .Y(_13530_));
NAND_g _19643_ (.A(_13453_), .B(_13530_), .Y(_13531_));
AND_g _19644_ (.A(_13452_), .B(_13531_), .Y(_13532_));
AND_g _19645_ (.A(_13450_), .B(_13532_), .Y(_13533_));
NOR_g _19646_ (.A(_13451_), .B(_13533_), .Y(_13534_));
NAND_g _19647_ (.A(_13449_), .B(_13534_), .Y(_13535_));
AND_g _19648_ (.A(_13448_), .B(_13535_), .Y(_13536_));
AND_g _19649_ (.A(_13447_), .B(_13536_), .Y(_13537_));
NOR_g _19650_ (.A(_13446_), .B(_13537_), .Y(_13538_));
NAND_g _19651_ (.A(_13445_), .B(_13538_), .Y(_13539_));
NAND_g _19652_ (.A(_13444_), .B(_13539_), .Y(_13540_));
XOR_g _19653_ (.A(decoded_imm[25]), .B(pcpi_rs1[25]), .Y(_13541_));
NAND_g _19654_ (.A(_13540_), .B(_13541_), .Y(_13542_));
NAND_g _19655_ (.A(_13443_), .B(_13542_), .Y(_13543_));
NAND_g _19656_ (.A(_13442_), .B(_13543_), .Y(_13544_));
AND_g _19657_ (.A(_13441_), .B(_13544_), .Y(_13545_));
AND_g _19658_ (.A(_13439_), .B(_13545_), .Y(_13546_));
NOR_g _19659_ (.A(_13440_), .B(_13546_), .Y(_13547_));
NAND_g _19660_ (.A(_13438_), .B(_13547_), .Y(_13548_));
AND_g _19661_ (.A(_13437_), .B(_13548_), .Y(_13549_));
AND_g _19662_ (.A(_13435_), .B(_13549_), .Y(_13550_));
NOR_g _19663_ (.A(_13436_), .B(_13550_), .Y(_13551_));
NAND_g _19664_ (.A(_13434_), .B(_13551_), .Y(_13552_));
NAND_g _19665_ (.A(_13433_), .B(_13552_), .Y(_13553_));
XNOR_g _19666_ (.A(pcpi_rs1[31]), .B(decoded_imm[31]), .Y(_13554_));
XNOR_g _19667_ (.A(_13553_), .B(_13554_), .Y(_13555_));
NAND_g _19668_ (.A(_13432_), .B(_13555_), .Y(_13556_));
NOR_g _19669_ (.A(decoded_imm_j[15]), .B(decoded_imm_j[16]), .Y(_13557_));
NOR_g _19670_ (.A(decoded_imm_j[17]), .B(decoded_imm_j[18]), .Y(_13558_));
AND_g _19671_ (.A(_11048_), .B(_13558_), .Y(_13559_));
AND_g _19672_ (.A(_13557_), .B(_13559_), .Y(_13560_));
NAND_g _19673_ (.A(_13557_), .B(_13559_), .Y(_13561_));
NOR_g _19674_ (.A(instr_rdinstr), .B(instr_rdinstrh), .Y(_13562_));
NOR_g _19675_ (.A(instr_rdcycle), .B(instr_rdcycleh), .Y(_13563_));
AND_g _19676_ (.A(_10973_), .B(_13562_), .Y(_13564_));
AND_g _19677_ (.A(_13562_), .B(_13563_), .Y(_13565_));
NAND_g _19678_ (.A(_13562_), .B(_13563_), .Y(_13566_));
NOR_g _19679_ (.A(instr_beq), .B(instr_jalr), .Y(_13567_));
NOR_g _19680_ (.A(instr_bgeu), .B(instr_bltu), .Y(_13568_));
AND_g _19681_ (.A(_10920_), .B(_13568_), .Y(_13569_));
NOR_g _19682_ (.A(instr_blt), .B(instr_bne), .Y(_13570_));
AND_g _19683_ (.A(_13569_), .B(_13570_), .Y(_13571_));
NAND_g _19684_ (.A(_10921_), .B(_13567_), .Y(_13572_));
AND_g _19685_ (.A(_13567_), .B(_13571_), .Y(_13573_));
NAND_g _19686_ (.A(_12521_), .B(_13573_), .Y(_13574_));
NOR_g _19687_ (.A(instr_and), .B(instr_or), .Y(_13575_));
AND_g _19688_ (.A(_10913_), .B(_13418_), .Y(_13576_));
AND_g _19689_ (.A(_13575_), .B(_13576_), .Y(_13577_));
NOR_g _19690_ (.A(instr_lb), .B(instr_lbu), .Y(_13578_));
NOR_g _19691_ (.A(instr_lh), .B(instr_lhu), .Y(_13579_));
NOR_g _19692_ (.A(instr_andi), .B(instr_slli), .Y(_13580_));
NOR_g _19693_ (.A(instr_slli), .B(instr_srli), .Y(_13581_));
AND_g _19694_ (.A(_10969_), .B(_13417_), .Y(_13582_));
AND_g _19695_ (.A(_13417_), .B(_13580_), .Y(_13583_));
NOR_g _19696_ (.A(instr_sb), .B(instr_sw), .Y(_13584_));
AND_g _19697_ (.A(_10967_), .B(_13584_), .Y(_13585_));
AND_g _19698_ (.A(_10917_), .B(_13585_), .Y(_13586_));
NOR_g _19699_ (.A(instr_slti), .B(instr_addi), .Y(_13587_));
AND_g _19700_ (.A(_10915_), .B(_13587_), .Y(_13588_));
AND_g _19701_ (.A(_13585_), .B(_13588_), .Y(_13589_));
NOR_g _19702_ (.A(instr_slt), .B(instr_sll), .Y(_13590_));
AND_g _19703_ (.A(_10908_), .B(_13590_), .Y(_13591_));
NOR_g _19704_ (.A(instr_xor), .B(instr_sltu), .Y(_13592_));
AND_g _19705_ (.A(_10907_), .B(_12531_), .Y(_13593_));
AND_g _19706_ (.A(_13590_), .B(_13592_), .Y(_13594_));
AND_g _19707_ (.A(_10910_), .B(_13590_), .Y(_13595_));
AND_g _19708_ (.A(_12522_), .B(_13590_), .Y(_13596_));
AND_g _19709_ (.A(_13592_), .B(_13596_), .Y(_13597_));
NOR_g _19710_ (.A(instr_ori), .B(instr_xori), .Y(_13598_));
AND_g _19711_ (.A(_13575_), .B(_13598_), .Y(_13599_));
NOR_g _19712_ (.A(instr_lw), .B(instr_lbu), .Y(_13600_));
AND_g _19713_ (.A(_13579_), .B(_13600_), .Y(_13601_));
AND_g _19714_ (.A(_13599_), .B(_13601_), .Y(_13602_));
NOR_g _19715_ (.A(instr_lb), .B(_13566_), .Y(_13603_));
AND_g _19716_ (.A(_13589_), .B(_13603_), .Y(_13604_));
AND_g _19717_ (.A(_13418_), .B(_13583_), .Y(_13605_));
AND_g _19718_ (.A(_13602_), .B(_13605_), .Y(_13606_));
NAND_g _19719_ (.A(_13597_), .B(_13606_), .Y(_13607_));
NOR_g _19720_ (.A(_13574_), .B(_13607_), .Y(_13608_));
AND_g _19721_ (.A(_13604_), .B(_13608_), .Y(_13609_));
NAND_g _19722_ (.A(_13604_), .B(_13608_), .Y(_13610_));
AND_g _19723_ (.A(_13565_), .B(_13610_), .Y(_13611_));
AND_g _19724_ (.A(_11209_), .B(_13611_), .Y(_13612_));
AND_g _19725_ (.A(_13561_), .B(_13612_), .Y(_13613_));
NAND_g _19726_ (.A(cpuregs_4[31]), .B(_11213_), .Y(_13614_));
NAND_g _19727_ (.A(cpuregs_6[31]), .B(_00012_[1]), .Y(_13615_));
AND_g _19728_ (.A(_00012_[2]), .B(_13615_), .Y(_13616_));
NAND_g _19729_ (.A(_13614_), .B(_13616_), .Y(_13617_));
NAND_g _19730_ (.A(cpuregs_0[31]), .B(_11213_), .Y(_13618_));
NAND_g _19731_ (.A(cpuregs_2[31]), .B(_00012_[1]), .Y(_13619_));
AND_g _19732_ (.A(_11214_), .B(_13619_), .Y(_13620_));
NAND_g _19733_ (.A(_13618_), .B(_13620_), .Y(_13621_));
AND_g _19734_ (.A(_11212_), .B(_13621_), .Y(_13622_));
NAND_g _19735_ (.A(_13617_), .B(_13622_), .Y(_13623_));
NAND_g _19736_ (.A(cpuregs_5[31]), .B(_11213_), .Y(_13624_));
NAND_g _19737_ (.A(cpuregs_7[31]), .B(_00012_[1]), .Y(_13625_));
AND_g _19738_ (.A(_00012_[2]), .B(_13625_), .Y(_13626_));
NAND_g _19739_ (.A(_13624_), .B(_13626_), .Y(_13627_));
NAND_g _19740_ (.A(cpuregs_1[31]), .B(_11213_), .Y(_13628_));
NAND_g _19741_ (.A(cpuregs_3[31]), .B(_00012_[1]), .Y(_13629_));
AND_g _19742_ (.A(_11214_), .B(_13629_), .Y(_13630_));
NAND_g _19743_ (.A(_13628_), .B(_13630_), .Y(_13631_));
AND_g _19744_ (.A(_00012_[0]), .B(_13631_), .Y(_13632_));
NAND_g _19745_ (.A(_13627_), .B(_13632_), .Y(_13633_));
NAND_g _19746_ (.A(_13623_), .B(_13633_), .Y(_13634_));
NAND_g _19747_ (.A(_11215_), .B(_13634_), .Y(_13635_));
NAND_g _19748_ (.A(cpuregs_10[31]), .B(_11214_), .Y(_13636_));
NAND_g _19749_ (.A(cpuregs_14[31]), .B(_00012_[2]), .Y(_13637_));
AND_g _19750_ (.A(_00012_[1]), .B(_13637_), .Y(_13638_));
NAND_g _19751_ (.A(_13636_), .B(_13638_), .Y(_13639_));
NAND_g _19752_ (.A(cpuregs_8[31]), .B(_11214_), .Y(_13640_));
NAND_g _19753_ (.A(cpuregs_12[31]), .B(_00012_[2]), .Y(_13641_));
AND_g _19754_ (.A(_11213_), .B(_13641_), .Y(_13642_));
NAND_g _19755_ (.A(_13640_), .B(_13642_), .Y(_13643_));
AND_g _19756_ (.A(_11212_), .B(_13643_), .Y(_13644_));
NAND_g _19757_ (.A(_13639_), .B(_13644_), .Y(_13645_));
NAND_g _19758_ (.A(cpuregs_15[31]), .B(_00012_[2]), .Y(_13646_));
NAND_g _19759_ (.A(cpuregs_11[31]), .B(_11214_), .Y(_13647_));
AND_g _19760_ (.A(_00012_[1]), .B(_13647_), .Y(_13648_));
NAND_g _19761_ (.A(_13646_), .B(_13648_), .Y(_13649_));
NAND_g _19762_ (.A(cpuregs_9[31]), .B(_11214_), .Y(_13650_));
NAND_g _19763_ (.A(cpuregs_13[31]), .B(_00012_[2]), .Y(_13651_));
AND_g _19764_ (.A(_11213_), .B(_13651_), .Y(_13652_));
NAND_g _19765_ (.A(_13650_), .B(_13652_), .Y(_13653_));
AND_g _19766_ (.A(_00012_[0]), .B(_13653_), .Y(_13654_));
NAND_g _19767_ (.A(_13649_), .B(_13654_), .Y(_13655_));
NAND_g _19768_ (.A(_13645_), .B(_13655_), .Y(_13656_));
NAND_g _19769_ (.A(_00012_[3]), .B(_13656_), .Y(_13657_));
AND_g _19770_ (.A(_13635_), .B(_13657_), .Y(_13658_));
NAND_g _19771_ (.A(_11216_), .B(_13658_), .Y(_13659_));
AND_g _19772_ (.A(_13409_), .B(_13659_), .Y(_13660_));
NAND_g _19773_ (.A(cpuregs_20[31]), .B(_00012_[2]), .Y(_13661_));
NAND_g _19774_ (.A(cpuregs_16[31]), .B(_11214_), .Y(_13662_));
AND_g _19775_ (.A(_13661_), .B(_13662_), .Y(_13663_));
NOR_g _19776_ (.A(_00012_[0]), .B(_13663_), .Y(_13664_));
NAND_g _19777_ (.A(_11039_), .B(_00012_[2]), .Y(_13665_));
NOR_g _19778_ (.A(cpuregs_17[31]), .B(_00012_[2]), .Y(_13666_));
NOR_g _19779_ (.A(_11212_), .B(_13666_), .Y(_13667_));
AND_g _19780_ (.A(_13665_), .B(_13667_), .Y(_13668_));
NOR_g _19781_ (.A(_13664_), .B(_13668_), .Y(_13669_));
NAND_g _19782_ (.A(_11213_), .B(_13669_), .Y(_13670_));
NAND_g _19783_ (.A(cpuregs_22[31]), .B(_00012_[2]), .Y(_13671_));
NAND_g _19784_ (.A(cpuregs_18[31]), .B(_11214_), .Y(_13672_));
AND_g _19785_ (.A(_13671_), .B(_13672_), .Y(_13673_));
NOR_g _19786_ (.A(_00012_[0]), .B(_13673_), .Y(_13674_));
NAND_g _19787_ (.A(_11192_), .B(_00012_[2]), .Y(_13675_));
NOR_g _19788_ (.A(cpuregs_19[31]), .B(_00012_[2]), .Y(_13676_));
NOR_g _19789_ (.A(_11212_), .B(_13676_), .Y(_13677_));
AND_g _19790_ (.A(_13675_), .B(_13677_), .Y(_13678_));
NOR_g _19791_ (.A(_13674_), .B(_13678_), .Y(_13679_));
NAND_g _19792_ (.A(_00012_[1]), .B(_13679_), .Y(_13680_));
AND_g _19793_ (.A(_13670_), .B(_13680_), .Y(_13681_));
NAND_g _19794_ (.A(cpuregs_27[31]), .B(_00012_[0]), .Y(_13682_));
NAND_g _19795_ (.A(cpuregs_26[31]), .B(_11212_), .Y(_13683_));
AND_g _19796_ (.A(_11214_), .B(_13683_), .Y(_13684_));
NAND_g _19797_ (.A(_13682_), .B(_13684_), .Y(_13685_));
NAND_g _19798_ (.A(cpuregs_31[31]), .B(_00012_[0]), .Y(_13686_));
NAND_g _19799_ (.A(cpuregs_30[31]), .B(_11212_), .Y(_13687_));
AND_g _19800_ (.A(_00012_[2]), .B(_13687_), .Y(_13688_));
NAND_g _19801_ (.A(_13686_), .B(_13688_), .Y(_13689_));
NAND_g _19802_ (.A(_13685_), .B(_13689_), .Y(_13690_));
NAND_g _19803_ (.A(_00012_[1]), .B(_13690_), .Y(_13691_));
NAND_g _19804_ (.A(cpuregs_25[31]), .B(_00012_[0]), .Y(_13692_));
NAND_g _19805_ (.A(cpuregs_24[31]), .B(_11212_), .Y(_13693_));
AND_g _19806_ (.A(_11214_), .B(_13693_), .Y(_13694_));
NAND_g _19807_ (.A(_13692_), .B(_13694_), .Y(_13695_));
NAND_g _19808_ (.A(cpuregs_29[31]), .B(_00012_[0]), .Y(_13696_));
NAND_g _19809_ (.A(cpuregs_28[31]), .B(_11212_), .Y(_13697_));
AND_g _19810_ (.A(_00012_[2]), .B(_13697_), .Y(_13698_));
NAND_g _19811_ (.A(_13696_), .B(_13698_), .Y(_13699_));
NAND_g _19812_ (.A(_13695_), .B(_13699_), .Y(_13700_));
NAND_g _19813_ (.A(_11213_), .B(_13700_), .Y(_13701_));
AND_g _19814_ (.A(_00012_[3]), .B(_13691_), .Y(_13702_));
NAND_g _19815_ (.A(_13701_), .B(_13702_), .Y(_13703_));
NAND_g _19816_ (.A(_11215_), .B(_13681_), .Y(_13704_));
AND_g _19817_ (.A(_13703_), .B(_13704_), .Y(_13705_));
NAND_g _19818_ (.A(_00012_[4]), .B(_13705_), .Y(_13706_));
NAND_g _19819_ (.A(pcpi_rs1[27]), .B(_13420_), .Y(_13707_));
NAND_g _19820_ (.A(pcpi_rs1[30]), .B(_13420_), .Y(_13708_));
NAND_g _19821_ (.A(_13382_), .B(_13708_), .Y(_13709_));
NAND_g _19822_ (.A(_13383_), .B(_13707_), .Y(_13710_));
AND_g _19823_ (.A(_13709_), .B(_13710_), .Y(_13711_));
NAND_g _19824_ (.A(_13389_), .B(_13711_), .Y(_13712_));
AND_g _19825_ (.A(_10979_), .B(is_lui_auipc_jal), .Y(_13713_));
AND_g _19826_ (.A(_13409_), .B(_13713_), .Y(_13714_));
NAND_g _19827_ (.A(reg_pc[31]), .B(_13714_), .Y(_13715_));
NAND_g _19828_ (.A(_13712_), .B(_13715_), .Y(_13716_));
AND_g _19829_ (.A(_13613_), .B(_13706_), .Y(_13717_));
AND_g _19830_ (.A(_13660_), .B(_13717_), .Y(_13718_));
NOR_g _19831_ (.A(_13716_), .B(_13718_), .Y(_13719_));
AND_g _19832_ (.A(_13556_), .B(_13719_), .Y(_13720_));
AND_g _19833_ (.A(_13426_), .B(_13720_), .Y(_13721_));
NOR_g _19834_ (.A(_13427_), .B(_13721_), .Y(_00502_));
NAND_g _19835_ (.A(cpu_state[4]), .B(_11267_), .Y(_13722_));
NOR_g _19836_ (.A(cpu_state[5]), .B(_13722_), .Y(_13723_));
AND_g _19837_ (.A(_11258_), .B(_13723_), .Y(_13724_));
NAND_g _19838_ (.A(_11258_), .B(_13723_), .Y(_13725_));
AND_g _19839_ (.A(_13410_), .B(_13725_), .Y(_13726_));
NOT_g _19840_ (.A(_13726_), .Y(dbg_ascii_state[46]));
AND_g _19841_ (.A(resetn), .B(dbg_ascii_state[46]), .Y(_13727_));
NAND_g _19842_ (.A(resetn), .B(dbg_ascii_state[46]), .Y(_13728_));
NOR_g _19843_ (.A(pcpi_rs2[0]), .B(_13727_), .Y(_13729_));
NOR_g _19844_ (.A(decoded_imm_j[11]), .B(decoded_imm_j[3]), .Y(_13730_));
NOR_g _19845_ (.A(decoded_imm_j[1]), .B(decoded_imm_j[2]), .Y(_13731_));
AND_g _19846_ (.A(_11049_), .B(_13731_), .Y(_13732_));
AND_g _19847_ (.A(_13730_), .B(_13732_), .Y(_13733_));
NAND_g _19848_ (.A(_13730_), .B(_13732_), .Y(_13734_));
NAND_g _19849_ (.A(_11171_), .B(_00011_[2]), .Y(_13735_));
NOR_g _19850_ (.A(cpuregs_26[0]), .B(_00011_[2]), .Y(_13736_));
NOR_g _19851_ (.A(_00011_[0]), .B(_13736_), .Y(_13737_));
NAND_g _19852_ (.A(_13735_), .B(_13737_), .Y(_13738_));
NAND_g _19853_ (.A(_11087_), .B(_00011_[2]), .Y(_13739_));
NOR_g _19854_ (.A(cpuregs_27[0]), .B(_00011_[2]), .Y(_13740_));
NOR_g _19855_ (.A(_11217_), .B(_13740_), .Y(_13741_));
NAND_g _19856_ (.A(_13739_), .B(_13741_), .Y(_13742_));
NAND_g _19857_ (.A(_13738_), .B(_13742_), .Y(_13743_));
NAND_g _19858_ (.A(_00011_[3]), .B(_13743_), .Y(_13744_));
NAND_g _19859_ (.A(cpuregs_22[0]), .B(_00011_[2]), .Y(_13745_));
NAND_g _19860_ (.A(cpuregs_18[0]), .B(_11219_), .Y(_13746_));
AND_g _19861_ (.A(_13745_), .B(_13746_), .Y(_13747_));
NAND_g _19862_ (.A(_11217_), .B(_13747_), .Y(_13748_));
NAND_g _19863_ (.A(cpuregs_23[0]), .B(_00011_[2]), .Y(_13749_));
NAND_g _19864_ (.A(cpuregs_19[0]), .B(_11219_), .Y(_13750_));
AND_g _19865_ (.A(_00011_[0]), .B(_13750_), .Y(_13751_));
NAND_g _19866_ (.A(_13749_), .B(_13751_), .Y(_13752_));
AND_g _19867_ (.A(_11220_), .B(_13752_), .Y(_13753_));
NAND_g _19868_ (.A(_13748_), .B(_13753_), .Y(_13754_));
AND_g _19869_ (.A(_13744_), .B(_13754_), .Y(_13755_));
NAND_g _19870_ (.A(cpuregs_6[0]), .B(_00011_[2]), .Y(_13756_));
NAND_g _19871_ (.A(cpuregs_2[0]), .B(_11219_), .Y(_13757_));
AND_g _19872_ (.A(_11217_), .B(_13757_), .Y(_13758_));
NAND_g _19873_ (.A(_13756_), .B(_13758_), .Y(_13759_));
NAND_g _19874_ (.A(cpuregs_3[0]), .B(_11219_), .Y(_13760_));
NAND_g _19875_ (.A(cpuregs_7[0]), .B(_00011_[2]), .Y(_13761_));
AND_g _19876_ (.A(_00011_[0]), .B(_13761_), .Y(_13762_));
NAND_g _19877_ (.A(_13760_), .B(_13762_), .Y(_13763_));
NOR_g _19878_ (.A(cpuregs_11[0]), .B(_00011_[2]), .Y(_13764_));
NAND_g _19879_ (.A(_11156_), .B(_00011_[2]), .Y(_13765_));
NOR_g _19880_ (.A(cpuregs_10[0]), .B(_00011_[2]), .Y(_13766_));
NOR_g _19881_ (.A(cpuregs_14[0]), .B(_11219_), .Y(_13767_));
NOR_g _19882_ (.A(_13766_), .B(_13767_), .Y(_13768_));
NAND_g _19883_ (.A(_13759_), .B(_13763_), .Y(_13769_));
NAND_g _19884_ (.A(_11220_), .B(_13769_), .Y(_13770_));
NAND_g _19885_ (.A(_11217_), .B(_13768_), .Y(_13771_));
NOR_g _19886_ (.A(_11217_), .B(_13764_), .Y(_13772_));
NAND_g _19887_ (.A(_13765_), .B(_13772_), .Y(_13773_));
AND_g _19888_ (.A(_00011_[3]), .B(_13773_), .Y(_13774_));
NAND_g _19889_ (.A(_13771_), .B(_13774_), .Y(_13775_));
NAND_g _19890_ (.A(_13770_), .B(_13775_), .Y(_13776_));
NAND_g _19891_ (.A(_11093_), .B(_00011_[2]), .Y(_13777_));
NOR_g _19892_ (.A(cpuregs_24[0]), .B(_00011_[2]), .Y(_13778_));
NOR_g _19893_ (.A(_00011_[0]), .B(_13778_), .Y(_13779_));
NAND_g _19894_ (.A(_13777_), .B(_13779_), .Y(_13780_));
NAND_g _19895_ (.A(_10922_), .B(_00011_[2]), .Y(_13781_));
NOR_g _19896_ (.A(cpuregs_25[0]), .B(_00011_[2]), .Y(_13782_));
NOR_g _19897_ (.A(_11217_), .B(_13782_), .Y(_13783_));
NAND_g _19898_ (.A(_13781_), .B(_13783_), .Y(_13784_));
NAND_g _19899_ (.A(_13780_), .B(_13784_), .Y(_13785_));
NAND_g _19900_ (.A(_00011_[3]), .B(_13785_), .Y(_13786_));
NAND_g _19901_ (.A(cpuregs_20[0]), .B(_00011_[2]), .Y(_13787_));
NAND_g _19902_ (.A(cpuregs_16[0]), .B(_11219_), .Y(_13788_));
AND_g _19903_ (.A(_13787_), .B(_13788_), .Y(_13789_));
NAND_g _19904_ (.A(_11217_), .B(_13789_), .Y(_13790_));
NAND_g _19905_ (.A(cpuregs_21[0]), .B(_00011_[2]), .Y(_13791_));
NAND_g _19906_ (.A(cpuregs_17[0]), .B(_11219_), .Y(_13792_));
AND_g _19907_ (.A(_00011_[0]), .B(_13792_), .Y(_13793_));
NAND_g _19908_ (.A(_13791_), .B(_13793_), .Y(_13794_));
AND_g _19909_ (.A(_11220_), .B(_13794_), .Y(_13795_));
NAND_g _19910_ (.A(_13790_), .B(_13795_), .Y(_13796_));
AND_g _19911_ (.A(_13786_), .B(_13796_), .Y(_13797_));
NAND_g _19912_ (.A(cpuregs_4[0]), .B(_00011_[2]), .Y(_13798_));
NAND_g _19913_ (.A(cpuregs_0[0]), .B(_11219_), .Y(_13799_));
AND_g _19914_ (.A(_11217_), .B(_13799_), .Y(_13800_));
NAND_g _19915_ (.A(_13798_), .B(_13800_), .Y(_13801_));
NAND_g _19916_ (.A(cpuregs_1[0]), .B(_11219_), .Y(_13802_));
NAND_g _19917_ (.A(cpuregs_5[0]), .B(_00011_[2]), .Y(_13803_));
AND_g _19918_ (.A(_00011_[0]), .B(_13803_), .Y(_13804_));
NAND_g _19919_ (.A(_13802_), .B(_13804_), .Y(_13805_));
NOR_g _19920_ (.A(cpuregs_8[0]), .B(_00011_[2]), .Y(_13806_));
NOR_g _19921_ (.A(cpuregs_12[0]), .B(_11219_), .Y(_13807_));
NOR_g _19922_ (.A(_13806_), .B(_13807_), .Y(_13808_));
NOR_g _19923_ (.A(cpuregs_9[0]), .B(_00011_[2]), .Y(_13809_));
NAND_g _19924_ (.A(_11139_), .B(_00011_[2]), .Y(_13810_));
NAND_g _19925_ (.A(_13801_), .B(_13805_), .Y(_13811_));
NAND_g _19926_ (.A(_11220_), .B(_13811_), .Y(_13812_));
NAND_g _19927_ (.A(_11217_), .B(_13808_), .Y(_13813_));
NOR_g _19928_ (.A(_11217_), .B(_13809_), .Y(_13814_));
NAND_g _19929_ (.A(_13810_), .B(_13814_), .Y(_13815_));
AND_g _19930_ (.A(_00011_[3]), .B(_13815_), .Y(_13816_));
NAND_g _19931_ (.A(_13813_), .B(_13816_), .Y(_13817_));
NAND_g _19932_ (.A(_13812_), .B(_13817_), .Y(_13818_));
NAND_g _19933_ (.A(_00011_[1]), .B(_13755_), .Y(_13819_));
NAND_g _19934_ (.A(_11218_), .B(_13797_), .Y(_13820_));
AND_g _19935_ (.A(_00011_[4]), .B(_13820_), .Y(_13821_));
NAND_g _19936_ (.A(_13819_), .B(_13821_), .Y(_13822_));
NAND_g _19937_ (.A(_00011_[1]), .B(_13776_), .Y(_13823_));
NAND_g _19938_ (.A(_11218_), .B(_13818_), .Y(_13824_));
AND_g _19939_ (.A(_13823_), .B(_13824_), .Y(_13825_));
NAND_g _19940_ (.A(_11221_), .B(_13825_), .Y(_13826_));
NAND_g _19941_ (.A(_13822_), .B(_13826_), .Y(_13827_));
AND_g _19942_ (.A(_13734_), .B(_13827_), .Y(_13828_));
NOR_g _19943_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi), .B(is_lui_auipc_jal), .Y(_13829_));
NAND_g _19944_ (.A(_10978_), .B(_11209_), .Y(_13830_));
NAND_g _19945_ (.A(_10977_), .B(_13611_), .Y(_13831_));
NOR_g _19946_ (.A(is_lb_lh_lw_lbu_lhu), .B(_13831_), .Y(_13832_));
AND_g _19947_ (.A(_13829_), .B(_13832_), .Y(_13833_));
NAND_g _19948_ (.A(_13829_), .B(_13832_), .Y(_13834_));
AND_g _19949_ (.A(_13828_), .B(_13833_), .Y(_13835_));
NAND_g _19950_ (.A(_13828_), .B(_13833_), .Y(_13836_));
NAND_g _19951_ (.A(decoded_imm[0]), .B(_13830_), .Y(_13837_));
NAND_g _19952_ (.A(_13836_), .B(_13837_), .Y(_13838_));
NAND_g _19953_ (.A(_13409_), .B(_13838_), .Y(_13839_));
AND_g _19954_ (.A(_13724_), .B(_13828_), .Y(_13840_));
NOR_g _19955_ (.A(_13728_), .B(_13840_), .Y(_13841_));
AND_g _19956_ (.A(_13839_), .B(_13841_), .Y(_13842_));
NOR_g _19957_ (.A(_13729_), .B(_13842_), .Y(_00503_));
NAND_g _19958_ (.A(_10982_), .B(_13728_), .Y(_13843_));
NAND_g _19959_ (.A(cpuregs_19[1]), .B(_11219_), .Y(_13844_));
NAND_g _19960_ (.A(cpuregs_23[1]), .B(_00011_[2]), .Y(_13845_));
AND_g _19961_ (.A(_00011_[0]), .B(_13845_), .Y(_13846_));
NAND_g _19962_ (.A(_13844_), .B(_13846_), .Y(_13847_));
NAND_g _19963_ (.A(cpuregs_18[1]), .B(_11219_), .Y(_13848_));
NAND_g _19964_ (.A(cpuregs_22[1]), .B(_00011_[2]), .Y(_13849_));
AND_g _19965_ (.A(_11217_), .B(_13849_), .Y(_13850_));
NAND_g _19966_ (.A(_13848_), .B(_13850_), .Y(_13851_));
AND_g _19967_ (.A(_11220_), .B(_13851_), .Y(_13852_));
NAND_g _19968_ (.A(_13847_), .B(_13852_), .Y(_13853_));
NAND_g _19969_ (.A(cpuregs_27[1]), .B(_11219_), .Y(_13854_));
NAND_g _19970_ (.A(cpuregs_31[1]), .B(_00011_[2]), .Y(_13855_));
AND_g _19971_ (.A(_00011_[0]), .B(_13855_), .Y(_13856_));
NAND_g _19972_ (.A(_13854_), .B(_13856_), .Y(_13857_));
NAND_g _19973_ (.A(cpuregs_26[1]), .B(_11219_), .Y(_13858_));
NAND_g _19974_ (.A(cpuregs_30[1]), .B(_00011_[2]), .Y(_13859_));
AND_g _19975_ (.A(_11217_), .B(_13859_), .Y(_13860_));
NAND_g _19976_ (.A(_13858_), .B(_13860_), .Y(_13861_));
AND_g _19977_ (.A(_00011_[3]), .B(_13861_), .Y(_13862_));
NAND_g _19978_ (.A(_13857_), .B(_13862_), .Y(_13863_));
NAND_g _19979_ (.A(_13853_), .B(_13863_), .Y(_13864_));
NAND_g _19980_ (.A(_00011_[1]), .B(_13864_), .Y(_13865_));
NAND_g _19981_ (.A(cpuregs_21[1]), .B(_00011_[2]), .Y(_13866_));
NAND_g _19982_ (.A(cpuregs_17[1]), .B(_11219_), .Y(_13867_));
AND_g _19983_ (.A(_00011_[0]), .B(_13867_), .Y(_13868_));
NAND_g _19984_ (.A(_13866_), .B(_13868_), .Y(_13869_));
NAND_g _19985_ (.A(cpuregs_20[1]), .B(_00011_[2]), .Y(_13870_));
NAND_g _19986_ (.A(cpuregs_16[1]), .B(_11219_), .Y(_13871_));
AND_g _19987_ (.A(_11217_), .B(_13871_), .Y(_13872_));
NAND_g _19988_ (.A(_13870_), .B(_13872_), .Y(_13873_));
AND_g _19989_ (.A(_11220_), .B(_13873_), .Y(_13874_));
NAND_g _19990_ (.A(_13869_), .B(_13874_), .Y(_13875_));
NAND_g _19991_ (.A(cpuregs_25[1]), .B(_11219_), .Y(_13876_));
NAND_g _19992_ (.A(cpuregs_29[1]), .B(_00011_[2]), .Y(_13877_));
AND_g _19993_ (.A(_00011_[0]), .B(_13877_), .Y(_13878_));
NAND_g _19994_ (.A(_13876_), .B(_13878_), .Y(_13879_));
NAND_g _19995_ (.A(cpuregs_24[1]), .B(_11219_), .Y(_13880_));
NAND_g _19996_ (.A(cpuregs_28[1]), .B(_00011_[2]), .Y(_13881_));
AND_g _19997_ (.A(_11217_), .B(_13881_), .Y(_13882_));
NAND_g _19998_ (.A(_13880_), .B(_13882_), .Y(_13883_));
AND_g _19999_ (.A(_00011_[3]), .B(_13883_), .Y(_13884_));
NAND_g _20000_ (.A(_13879_), .B(_13884_), .Y(_13885_));
NAND_g _20001_ (.A(_13875_), .B(_13885_), .Y(_13886_));
NAND_g _20002_ (.A(_11218_), .B(_13886_), .Y(_13887_));
NAND_g _20003_ (.A(_13865_), .B(_13887_), .Y(_13888_));
NAND_g _20004_ (.A(_00011_[4]), .B(_13888_), .Y(_13889_));
NAND_g _20005_ (.A(cpuregs_6[1]), .B(_00011_[2]), .Y(_13890_));
NAND_g _20006_ (.A(cpuregs_2[1]), .B(_11219_), .Y(_13891_));
AND_g _20007_ (.A(_13890_), .B(_13891_), .Y(_13892_));
NAND_g _20008_ (.A(_11217_), .B(_13892_), .Y(_13893_));
NAND_g _20009_ (.A(cpuregs_7[1]), .B(_00011_[2]), .Y(_13894_));
NAND_g _20010_ (.A(cpuregs_3[1]), .B(_11219_), .Y(_13895_));
AND_g _20011_ (.A(_00011_[0]), .B(_13895_), .Y(_13896_));
NAND_g _20012_ (.A(_13894_), .B(_13896_), .Y(_13897_));
AND_g _20013_ (.A(_11220_), .B(_13897_), .Y(_13898_));
NAND_g _20014_ (.A(_13893_), .B(_13898_), .Y(_13899_));
NOR_g _20015_ (.A(cpuregs_10[1]), .B(_00011_[2]), .Y(_13900_));
NOR_g _20016_ (.A(cpuregs_14[1]), .B(_11219_), .Y(_13901_));
NOR_g _20017_ (.A(_13900_), .B(_13901_), .Y(_13902_));
NOR_g _20018_ (.A(cpuregs_11[1]), .B(_00011_[2]), .Y(_13903_));
NOT_g _20019_ (.A(_13903_), .Y(_13904_));
NAND_g _20020_ (.A(_11157_), .B(_00011_[2]), .Y(_13905_));
AND_g _20021_ (.A(_00011_[0]), .B(_13905_), .Y(_13906_));
NAND_g _20022_ (.A(_13904_), .B(_13906_), .Y(_13907_));
NAND_g _20023_ (.A(_11217_), .B(_13902_), .Y(_13908_));
NAND_g _20024_ (.A(_13907_), .B(_13908_), .Y(_13909_));
NAND_g _20025_ (.A(_00011_[3]), .B(_13909_), .Y(_13910_));
AND_g _20026_ (.A(_13899_), .B(_13910_), .Y(_13911_));
NAND_g _20027_ (.A(cpuregs_4[1]), .B(_00011_[2]), .Y(_13912_));
NAND_g _20028_ (.A(cpuregs_0[1]), .B(_11219_), .Y(_13913_));
AND_g _20029_ (.A(_11217_), .B(_13913_), .Y(_13914_));
NAND_g _20030_ (.A(_13912_), .B(_13914_), .Y(_13915_));
NAND_g _20031_ (.A(cpuregs_1[1]), .B(_11219_), .Y(_13916_));
NAND_g _20032_ (.A(cpuregs_5[1]), .B(_00011_[2]), .Y(_13917_));
AND_g _20033_ (.A(_00011_[0]), .B(_13917_), .Y(_13918_));
NAND_g _20034_ (.A(_13916_), .B(_13918_), .Y(_13919_));
NOR_g _20035_ (.A(cpuregs_9[1]), .B(_00011_[2]), .Y(_13920_));
NAND_g _20036_ (.A(_11140_), .B(_00011_[2]), .Y(_13921_));
NOR_g _20037_ (.A(cpuregs_8[1]), .B(_00011_[2]), .Y(_13922_));
NOR_g _20038_ (.A(cpuregs_12[1]), .B(_11219_), .Y(_13923_));
NOR_g _20039_ (.A(_13922_), .B(_13923_), .Y(_13924_));
NAND_g _20040_ (.A(_13915_), .B(_13919_), .Y(_13925_));
NAND_g _20041_ (.A(_11220_), .B(_13925_), .Y(_13926_));
NAND_g _20042_ (.A(_11217_), .B(_13924_), .Y(_13927_));
NOR_g _20043_ (.A(_11217_), .B(_13920_), .Y(_13928_));
NAND_g _20044_ (.A(_13921_), .B(_13928_), .Y(_13929_));
AND_g _20045_ (.A(_00011_[3]), .B(_13929_), .Y(_13930_));
NAND_g _20046_ (.A(_13927_), .B(_13930_), .Y(_13931_));
NAND_g _20047_ (.A(_13926_), .B(_13931_), .Y(_13932_));
NAND_g _20048_ (.A(_11218_), .B(_13932_), .Y(_13933_));
NAND_g _20049_ (.A(_00011_[1]), .B(_13911_), .Y(_13934_));
AND_g _20050_ (.A(_13933_), .B(_13934_), .Y(_13935_));
NAND_g _20051_ (.A(_11221_), .B(_13935_), .Y(_13936_));
NAND_g _20052_ (.A(_13889_), .B(_13936_), .Y(_13937_));
AND_g _20053_ (.A(_13734_), .B(_13937_), .Y(_13938_));
AND_g _20054_ (.A(_13409_), .B(_13833_), .Y(_13939_));
NAND_g _20055_ (.A(_13409_), .B(_13833_), .Y(_13940_));
NAND_g _20056_ (.A(_13938_), .B(_13939_), .Y(_13941_));
NAND_g _20057_ (.A(_13724_), .B(_13938_), .Y(_13942_));
NOT_g _20058_ (.A(_13942_), .Y(_13943_));
AND_g _20059_ (.A(decoded_imm[1]), .B(_13830_), .Y(_13944_));
NAND_g _20060_ (.A(_13409_), .B(_13944_), .Y(_13945_));
AND_g _20061_ (.A(_13727_), .B(_13945_), .Y(_13946_));
AND_g _20062_ (.A(_13942_), .B(_13946_), .Y(_13947_));
NAND_g _20063_ (.A(_13833_), .B(_13938_), .Y(_13948_));
NAND_g _20064_ (.A(_13941_), .B(_13947_), .Y(_13949_));
AND_g _20065_ (.A(_13843_), .B(_13949_), .Y(_00504_));
NAND_g _20066_ (.A(_10983_), .B(_13728_), .Y(_13950_));
NAND_g _20067_ (.A(cpuregs_31[2]), .B(_00011_[1]), .Y(_13951_));
NAND_g _20068_ (.A(cpuregs_29[2]), .B(_11218_), .Y(_13952_));
NAND_g _20069_ (.A(_13951_), .B(_13952_), .Y(_13953_));
NAND_g _20070_ (.A(_00011_[2]), .B(_13953_), .Y(_13954_));
NAND_g _20071_ (.A(cpuregs_27[2]), .B(_00011_[1]), .Y(_13955_));
NAND_g _20072_ (.A(cpuregs_25[2]), .B(_11218_), .Y(_13956_));
NAND_g _20073_ (.A(_13955_), .B(_13956_), .Y(_13957_));
NAND_g _20074_ (.A(_11219_), .B(_13957_), .Y(_13958_));
NAND_g _20075_ (.A(_13954_), .B(_13958_), .Y(_13959_));
NAND_g _20076_ (.A(_00011_[0]), .B(_13959_), .Y(_13960_));
NAND_g _20077_ (.A(cpuregs_30[2]), .B(_00011_[1]), .Y(_13961_));
NAND_g _20078_ (.A(cpuregs_28[2]), .B(_11218_), .Y(_13962_));
NAND_g _20079_ (.A(_13961_), .B(_13962_), .Y(_13963_));
NAND_g _20080_ (.A(_00011_[2]), .B(_13963_), .Y(_13964_));
NAND_g _20081_ (.A(cpuregs_26[2]), .B(_00011_[1]), .Y(_13965_));
NAND_g _20082_ (.A(cpuregs_24[2]), .B(_11218_), .Y(_13966_));
NAND_g _20083_ (.A(_13965_), .B(_13966_), .Y(_13967_));
NAND_g _20084_ (.A(_11219_), .B(_13967_), .Y(_13968_));
NAND_g _20085_ (.A(_13964_), .B(_13968_), .Y(_13969_));
AND_g _20086_ (.A(_11217_), .B(_13969_), .Y(_13970_));
NOT_g _20087_ (.A(_13970_), .Y(_13971_));
NAND_g _20088_ (.A(_13960_), .B(_13971_), .Y(_13972_));
NAND_g _20089_ (.A(_00011_[3]), .B(_13972_), .Y(_13973_));
NOR_g _20090_ (.A(cpuregs_18[2]), .B(_00011_[2]), .Y(_13974_));
NOR_g _20091_ (.A(cpuregs_22[2]), .B(_11219_), .Y(_13975_));
NOR_g _20092_ (.A(_13974_), .B(_13975_), .Y(_13976_));
NOR_g _20093_ (.A(cpuregs_16[2]), .B(_00011_[2]), .Y(_13977_));
NOR_g _20094_ (.A(cpuregs_20[2]), .B(_11219_), .Y(_13978_));
NOR_g _20095_ (.A(_13977_), .B(_13978_), .Y(_13979_));
NAND_g _20096_ (.A(_11178_), .B(_00011_[2]), .Y(_13980_));
NOR_g _20097_ (.A(cpuregs_19[2]), .B(_00011_[2]), .Y(_13981_));
NOR_g _20098_ (.A(cpuregs_17[2]), .B(_00011_[2]), .Y(_13982_));
NAND_g _20099_ (.A(_11023_), .B(_00011_[2]), .Y(_13983_));
NOR_g _20100_ (.A(_11217_), .B(_13981_), .Y(_13984_));
NAND_g _20101_ (.A(_13980_), .B(_13984_), .Y(_13985_));
NAND_g _20102_ (.A(_11217_), .B(_13976_), .Y(_13986_));
AND_g _20103_ (.A(_13985_), .B(_13986_), .Y(_13987_));
NAND_g _20104_ (.A(_00011_[1]), .B(_13987_), .Y(_13988_));
NOR_g _20105_ (.A(_11217_), .B(_13982_), .Y(_13989_));
NAND_g _20106_ (.A(_13983_), .B(_13989_), .Y(_13990_));
NAND_g _20107_ (.A(_11217_), .B(_13979_), .Y(_13991_));
AND_g _20108_ (.A(_13990_), .B(_13991_), .Y(_13992_));
NAND_g _20109_ (.A(_11218_), .B(_13992_), .Y(_13993_));
AND_g _20110_ (.A(_13988_), .B(_13993_), .Y(_13994_));
NAND_g _20111_ (.A(_11220_), .B(_13994_), .Y(_13995_));
AND_g _20112_ (.A(_13973_), .B(_13995_), .Y(_13996_));
NAND_g _20113_ (.A(cpuregs_13[2]), .B(_11218_), .Y(_13997_));
NAND_g _20114_ (.A(cpuregs_15[2]), .B(_00011_[1]), .Y(_13998_));
AND_g _20115_ (.A(_00011_[2]), .B(_13998_), .Y(_13999_));
NAND_g _20116_ (.A(_13997_), .B(_13999_), .Y(_14000_));
NAND_g _20117_ (.A(cpuregs_9[2]), .B(_11218_), .Y(_14001_));
NAND_g _20118_ (.A(cpuregs_11[2]), .B(_00011_[1]), .Y(_14002_));
AND_g _20119_ (.A(_11219_), .B(_14002_), .Y(_14003_));
NAND_g _20120_ (.A(_14001_), .B(_14003_), .Y(_14004_));
AND_g _20121_ (.A(_00011_[0]), .B(_14004_), .Y(_14005_));
NAND_g _20122_ (.A(_14000_), .B(_14005_), .Y(_14006_));
NAND_g _20123_ (.A(cpuregs_12[2]), .B(_11218_), .Y(_14007_));
NAND_g _20124_ (.A(cpuregs_14[2]), .B(_00011_[1]), .Y(_14008_));
AND_g _20125_ (.A(_00011_[2]), .B(_14008_), .Y(_14009_));
NAND_g _20126_ (.A(_14007_), .B(_14009_), .Y(_14010_));
NAND_g _20127_ (.A(cpuregs_8[2]), .B(_11218_), .Y(_14011_));
NAND_g _20128_ (.A(cpuregs_10[2]), .B(_00011_[1]), .Y(_14012_));
AND_g _20129_ (.A(_11219_), .B(_14012_), .Y(_14013_));
NAND_g _20130_ (.A(_14011_), .B(_14013_), .Y(_14014_));
AND_g _20131_ (.A(_11217_), .B(_14014_), .Y(_14015_));
NAND_g _20132_ (.A(_14010_), .B(_14015_), .Y(_14016_));
NAND_g _20133_ (.A(_14006_), .B(_14016_), .Y(_14017_));
NAND_g _20134_ (.A(_00011_[3]), .B(_14017_), .Y(_14018_));
NAND_g _20135_ (.A(_10937_), .B(_00011_[2]), .Y(_14019_));
NOR_g _20136_ (.A(cpuregs_2[2]), .B(_00011_[2]), .Y(_14020_));
NOR_g _20137_ (.A(_00011_[0]), .B(_14020_), .Y(_14021_));
NAND_g _20138_ (.A(_14019_), .B(_14021_), .Y(_14022_));
NAND_g _20139_ (.A(_11123_), .B(_00011_[2]), .Y(_14023_));
NOR_g _20140_ (.A(cpuregs_3[2]), .B(_00011_[2]), .Y(_14024_));
NOR_g _20141_ (.A(_11217_), .B(_14024_), .Y(_14025_));
NAND_g _20142_ (.A(_14023_), .B(_14025_), .Y(_14026_));
AND_g _20143_ (.A(_14022_), .B(_14026_), .Y(_14027_));
NAND_g _20144_ (.A(_10949_), .B(_00011_[2]), .Y(_14028_));
NOR_g _20145_ (.A(cpuregs_0[2]), .B(_00011_[2]), .Y(_14029_));
NOR_g _20146_ (.A(_00011_[0]), .B(_14029_), .Y(_14030_));
NAND_g _20147_ (.A(_14028_), .B(_14030_), .Y(_14031_));
NAND_g _20148_ (.A(_11107_), .B(_00011_[2]), .Y(_14032_));
NOR_g _20149_ (.A(cpuregs_1[2]), .B(_00011_[2]), .Y(_14033_));
NOR_g _20150_ (.A(_11217_), .B(_14033_), .Y(_14034_));
NAND_g _20151_ (.A(_14032_), .B(_14034_), .Y(_14035_));
AND_g _20152_ (.A(_14031_), .B(_14035_), .Y(_14036_));
NAND_g _20153_ (.A(_00011_[1]), .B(_14027_), .Y(_14037_));
NAND_g _20154_ (.A(_11218_), .B(_14036_), .Y(_14038_));
AND_g _20155_ (.A(_14037_), .B(_14038_), .Y(_14039_));
NAND_g _20156_ (.A(_11220_), .B(_14039_), .Y(_14040_));
AND_g _20157_ (.A(_14018_), .B(_14040_), .Y(_14041_));
NAND_g _20158_ (.A(_00011_[4]), .B(_13996_), .Y(_14042_));
NAND_g _20159_ (.A(_11221_), .B(_14041_), .Y(_14043_));
AND_g _20160_ (.A(_13734_), .B(_14043_), .Y(_14044_));
AND_g _20161_ (.A(_14042_), .B(_14044_), .Y(_14045_));
NAND_g _20162_ (.A(_13939_), .B(_14045_), .Y(_14046_));
NAND_g _20163_ (.A(_13724_), .B(_14045_), .Y(_14047_));
AND_g _20164_ (.A(decoded_imm[2]), .B(_13830_), .Y(_14048_));
NAND_g _20165_ (.A(_13409_), .B(_14048_), .Y(_14049_));
AND_g _20166_ (.A(_13727_), .B(_14049_), .Y(_14050_));
AND_g _20167_ (.A(_14047_), .B(_14050_), .Y(_14051_));
NAND_g _20168_ (.A(_14046_), .B(_14051_), .Y(_14052_));
AND_g _20169_ (.A(_13950_), .B(_14052_), .Y(_00505_));
NOR_g _20170_ (.A(pcpi_rs2[3]), .B(_13727_), .Y(_14053_));
NAND_g _20171_ (.A(cpuregs_29[3]), .B(_00011_[2]), .Y(_14054_));
NAND_g _20172_ (.A(cpuregs_25[3]), .B(_11219_), .Y(_14055_));
AND_g _20173_ (.A(_00011_[0]), .B(_14055_), .Y(_14056_));
NAND_g _20174_ (.A(_14054_), .B(_14056_), .Y(_14057_));
NAND_g _20175_ (.A(cpuregs_24[3]), .B(_11219_), .Y(_14058_));
NAND_g _20176_ (.A(cpuregs_28[3]), .B(_00011_[2]), .Y(_14059_));
AND_g _20177_ (.A(_11217_), .B(_14059_), .Y(_14060_));
NAND_g _20178_ (.A(_14058_), .B(_14060_), .Y(_14061_));
AND_g _20179_ (.A(_11218_), .B(_14061_), .Y(_14062_));
NAND_g _20180_ (.A(_14057_), .B(_14062_), .Y(_14063_));
NAND_g _20181_ (.A(cpuregs_27[3]), .B(_11219_), .Y(_14064_));
NAND_g _20182_ (.A(cpuregs_31[3]), .B(_00011_[2]), .Y(_14065_));
AND_g _20183_ (.A(_00011_[0]), .B(_14065_), .Y(_14066_));
NAND_g _20184_ (.A(_14064_), .B(_14066_), .Y(_14067_));
NAND_g _20185_ (.A(cpuregs_26[3]), .B(_11219_), .Y(_14068_));
NAND_g _20186_ (.A(cpuregs_30[3]), .B(_00011_[2]), .Y(_14069_));
AND_g _20187_ (.A(_11217_), .B(_14069_), .Y(_14070_));
NAND_g _20188_ (.A(_14068_), .B(_14070_), .Y(_14071_));
AND_g _20189_ (.A(_00011_[1]), .B(_14071_), .Y(_14072_));
NAND_g _20190_ (.A(_14067_), .B(_14072_), .Y(_14073_));
NAND_g _20191_ (.A(_14063_), .B(_14073_), .Y(_14074_));
NAND_g _20192_ (.A(_00011_[4]), .B(_14074_), .Y(_14075_));
NAND_g _20193_ (.A(cpuregs_14[3]), .B(_11217_), .Y(_14076_));
NAND_g _20194_ (.A(cpuregs_15[3]), .B(_00011_[0]), .Y(_14077_));
NAND_g _20195_ (.A(_14076_), .B(_14077_), .Y(_14078_));
NAND_g _20196_ (.A(_00011_[2]), .B(_14078_), .Y(_14079_));
NAND_g _20197_ (.A(cpuregs_10[3]), .B(_11217_), .Y(_14080_));
NAND_g _20198_ (.A(cpuregs_11[3]), .B(_00011_[0]), .Y(_14081_));
NAND_g _20199_ (.A(_14080_), .B(_14081_), .Y(_14082_));
NAND_g _20200_ (.A(_11219_), .B(_14082_), .Y(_14083_));
NAND_g _20201_ (.A(_14079_), .B(_14083_), .Y(_14084_));
NAND_g _20202_ (.A(_00011_[1]), .B(_14084_), .Y(_14085_));
NAND_g _20203_ (.A(cpuregs_12[3]), .B(_11217_), .Y(_14086_));
NAND_g _20204_ (.A(cpuregs_13[3]), .B(_00011_[0]), .Y(_14087_));
NAND_g _20205_ (.A(_14086_), .B(_14087_), .Y(_14088_));
NAND_g _20206_ (.A(_00011_[2]), .B(_14088_), .Y(_14089_));
NAND_g _20207_ (.A(cpuregs_8[3]), .B(_11217_), .Y(_14090_));
NAND_g _20208_ (.A(cpuregs_9[3]), .B(_00011_[0]), .Y(_14091_));
NAND_g _20209_ (.A(_14090_), .B(_14091_), .Y(_14092_));
NAND_g _20210_ (.A(_11219_), .B(_14092_), .Y(_14093_));
NAND_g _20211_ (.A(_14089_), .B(_14093_), .Y(_14094_));
NAND_g _20212_ (.A(_11218_), .B(_14094_), .Y(_14095_));
NAND_g _20213_ (.A(_14085_), .B(_14095_), .Y(_14096_));
AND_g _20214_ (.A(_11221_), .B(_14096_), .Y(_14097_));
NOT_g _20215_ (.A(_14097_), .Y(_14098_));
NAND_g _20216_ (.A(_14075_), .B(_14098_), .Y(_14099_));
NAND_g _20217_ (.A(_00011_[3]), .B(_14099_), .Y(_14100_));
NAND_g _20218_ (.A(cpuregs_1[3]), .B(_11219_), .Y(_14101_));
NAND_g _20219_ (.A(cpuregs_5[3]), .B(_00011_[2]), .Y(_14102_));
AND_g _20220_ (.A(_00011_[0]), .B(_14102_), .Y(_14103_));
NAND_g _20221_ (.A(_14101_), .B(_14103_), .Y(_14104_));
NAND_g _20222_ (.A(cpuregs_0[3]), .B(_11219_), .Y(_14105_));
NAND_g _20223_ (.A(cpuregs_4[3]), .B(_00011_[2]), .Y(_14106_));
AND_g _20224_ (.A(_11217_), .B(_14106_), .Y(_14107_));
NAND_g _20225_ (.A(_14105_), .B(_14107_), .Y(_14108_));
AND_g _20226_ (.A(_11218_), .B(_14108_), .Y(_14109_));
NAND_g _20227_ (.A(_14104_), .B(_14109_), .Y(_14110_));
NAND_g _20228_ (.A(cpuregs_3[3]), .B(_11219_), .Y(_14111_));
NAND_g _20229_ (.A(cpuregs_7[3]), .B(_00011_[2]), .Y(_14112_));
AND_g _20230_ (.A(_00011_[0]), .B(_14112_), .Y(_14113_));
NAND_g _20231_ (.A(_14111_), .B(_14113_), .Y(_14114_));
NAND_g _20232_ (.A(cpuregs_2[3]), .B(_11219_), .Y(_14115_));
NAND_g _20233_ (.A(cpuregs_6[3]), .B(_00011_[2]), .Y(_14116_));
AND_g _20234_ (.A(_11217_), .B(_14116_), .Y(_14117_));
NAND_g _20235_ (.A(_14115_), .B(_14117_), .Y(_14118_));
AND_g _20236_ (.A(_00011_[1]), .B(_14118_), .Y(_14119_));
NAND_g _20237_ (.A(_14114_), .B(_14119_), .Y(_14120_));
NAND_g _20238_ (.A(_14110_), .B(_14120_), .Y(_14121_));
NAND_g _20239_ (.A(_11221_), .B(_14121_), .Y(_14122_));
NAND_g _20240_ (.A(cpuregs_19[3]), .B(_00011_[1]), .Y(_14123_));
NAND_g _20241_ (.A(cpuregs_17[3]), .B(_11218_), .Y(_14124_));
NAND_g _20242_ (.A(_14123_), .B(_14124_), .Y(_14125_));
NAND_g _20243_ (.A(_11219_), .B(_14125_), .Y(_14126_));
NAND_g _20244_ (.A(cpuregs_23[3]), .B(_00011_[1]), .Y(_14127_));
NAND_g _20245_ (.A(cpuregs_21[3]), .B(_11218_), .Y(_14128_));
NAND_g _20246_ (.A(_14127_), .B(_14128_), .Y(_14129_));
NAND_g _20247_ (.A(_00011_[2]), .B(_14129_), .Y(_14130_));
AND_g _20248_ (.A(_00011_[0]), .B(_14130_), .Y(_14131_));
NAND_g _20249_ (.A(_14126_), .B(_14131_), .Y(_14132_));
NAND_g _20250_ (.A(cpuregs_18[3]), .B(_00011_[1]), .Y(_14133_));
NAND_g _20251_ (.A(cpuregs_16[3]), .B(_11218_), .Y(_14134_));
NAND_g _20252_ (.A(_14133_), .B(_14134_), .Y(_14135_));
NAND_g _20253_ (.A(_11219_), .B(_14135_), .Y(_14136_));
NAND_g _20254_ (.A(cpuregs_22[3]), .B(_00011_[1]), .Y(_14137_));
NAND_g _20255_ (.A(cpuregs_20[3]), .B(_11218_), .Y(_14138_));
NAND_g _20256_ (.A(_14137_), .B(_14138_), .Y(_14139_));
NAND_g _20257_ (.A(_00011_[2]), .B(_14139_), .Y(_14140_));
AND_g _20258_ (.A(_11217_), .B(_14140_), .Y(_14141_));
NAND_g _20259_ (.A(_14136_), .B(_14141_), .Y(_14142_));
AND_g _20260_ (.A(_00011_[4]), .B(_14142_), .Y(_14143_));
NAND_g _20261_ (.A(_14132_), .B(_14143_), .Y(_14144_));
NAND_g _20262_ (.A(_14122_), .B(_14144_), .Y(_14145_));
NAND_g _20263_ (.A(_11220_), .B(_14145_), .Y(_14146_));
NAND_g _20264_ (.A(_14100_), .B(_14146_), .Y(_14147_));
AND_g _20265_ (.A(_13734_), .B(_14147_), .Y(_14148_));
AND_g _20266_ (.A(_13833_), .B(_14148_), .Y(_14149_));
NAND_g _20267_ (.A(_13833_), .B(_14148_), .Y(_14150_));
NAND_g _20268_ (.A(decoded_imm[3]), .B(_13830_), .Y(_14151_));
NAND_g _20269_ (.A(_14150_), .B(_14151_), .Y(_14152_));
NAND_g _20270_ (.A(_13409_), .B(_14152_), .Y(_14153_));
AND_g _20271_ (.A(_13724_), .B(_14148_), .Y(_14154_));
NOR_g _20272_ (.A(_13728_), .B(_14154_), .Y(_14155_));
AND_g _20273_ (.A(_14153_), .B(_14155_), .Y(_14156_));
NOR_g _20274_ (.A(_14053_), .B(_14156_), .Y(_00506_));
NAND_g _20275_ (.A(_10984_), .B(_13728_), .Y(_14157_));
NAND_g _20276_ (.A(_11094_), .B(_00011_[2]), .Y(_14158_));
NOR_g _20277_ (.A(cpuregs_24[4]), .B(_00011_[2]), .Y(_14159_));
NOR_g _20278_ (.A(_00011_[0]), .B(_14159_), .Y(_14160_));
NAND_g _20279_ (.A(_14158_), .B(_14160_), .Y(_14161_));
NAND_g _20280_ (.A(_10923_), .B(_00011_[2]), .Y(_14162_));
NOR_g _20281_ (.A(cpuregs_25[4]), .B(_00011_[2]), .Y(_14163_));
NOR_g _20282_ (.A(_11217_), .B(_14163_), .Y(_14164_));
NAND_g _20283_ (.A(_14162_), .B(_14164_), .Y(_14165_));
NAND_g _20284_ (.A(_14161_), .B(_14165_), .Y(_14166_));
NAND_g _20285_ (.A(_00011_[3]), .B(_14166_), .Y(_14167_));
NAND_g _20286_ (.A(cpuregs_20[4]), .B(_00011_[2]), .Y(_14168_));
NAND_g _20287_ (.A(cpuregs_16[4]), .B(_11219_), .Y(_14169_));
AND_g _20288_ (.A(_14168_), .B(_14169_), .Y(_14170_));
NAND_g _20289_ (.A(_11217_), .B(_14170_), .Y(_14171_));
NAND_g _20290_ (.A(cpuregs_21[4]), .B(_00011_[2]), .Y(_14172_));
NAND_g _20291_ (.A(cpuregs_17[4]), .B(_11219_), .Y(_14173_));
AND_g _20292_ (.A(_00011_[0]), .B(_14173_), .Y(_14174_));
NAND_g _20293_ (.A(_14172_), .B(_14174_), .Y(_14175_));
AND_g _20294_ (.A(_11220_), .B(_14175_), .Y(_14176_));
NAND_g _20295_ (.A(_14171_), .B(_14176_), .Y(_14177_));
AND_g _20296_ (.A(_14167_), .B(_14177_), .Y(_14178_));
NAND_g _20297_ (.A(cpuregs_4[4]), .B(_00011_[2]), .Y(_14179_));
NAND_g _20298_ (.A(cpuregs_0[4]), .B(_11219_), .Y(_14180_));
AND_g _20299_ (.A(_11217_), .B(_14180_), .Y(_14181_));
NAND_g _20300_ (.A(_14179_), .B(_14181_), .Y(_14182_));
NAND_g _20301_ (.A(cpuregs_1[4]), .B(_11219_), .Y(_14183_));
NAND_g _20302_ (.A(cpuregs_5[4]), .B(_00011_[2]), .Y(_14184_));
AND_g _20303_ (.A(_00011_[0]), .B(_14184_), .Y(_14185_));
NAND_g _20304_ (.A(_14183_), .B(_14185_), .Y(_14186_));
NOR_g _20305_ (.A(cpuregs_8[4]), .B(_00011_[2]), .Y(_14187_));
NOR_g _20306_ (.A(cpuregs_12[4]), .B(_11219_), .Y(_14188_));
NOR_g _20307_ (.A(_14187_), .B(_14188_), .Y(_14189_));
NOR_g _20308_ (.A(cpuregs_9[4]), .B(_00011_[2]), .Y(_14190_));
NAND_g _20309_ (.A(_11141_), .B(_00011_[2]), .Y(_14191_));
NAND_g _20310_ (.A(_14182_), .B(_14186_), .Y(_14192_));
NAND_g _20311_ (.A(_11220_), .B(_14192_), .Y(_14193_));
NAND_g _20312_ (.A(_11217_), .B(_14189_), .Y(_14194_));
NOR_g _20313_ (.A(_11217_), .B(_14190_), .Y(_14195_));
NAND_g _20314_ (.A(_14191_), .B(_14195_), .Y(_14196_));
AND_g _20315_ (.A(_00011_[3]), .B(_14196_), .Y(_14197_));
NAND_g _20316_ (.A(_14194_), .B(_14197_), .Y(_14198_));
NAND_g _20317_ (.A(_14193_), .B(_14198_), .Y(_14199_));
NAND_g _20318_ (.A(_11172_), .B(_00011_[2]), .Y(_14200_));
NOR_g _20319_ (.A(cpuregs_26[4]), .B(_00011_[2]), .Y(_14201_));
NOR_g _20320_ (.A(_00011_[0]), .B(_14201_), .Y(_14202_));
NAND_g _20321_ (.A(_14200_), .B(_14202_), .Y(_14203_));
NOR_g _20322_ (.A(cpuregs_27[4]), .B(_00011_[2]), .Y(_14204_));
NAND_g _20323_ (.A(_11088_), .B(_00011_[2]), .Y(_14205_));
NOR_g _20324_ (.A(_11217_), .B(_14204_), .Y(_14206_));
NAND_g _20325_ (.A(_14205_), .B(_14206_), .Y(_14207_));
NAND_g _20326_ (.A(_14203_), .B(_14207_), .Y(_14208_));
NAND_g _20327_ (.A(_00011_[3]), .B(_14208_), .Y(_14209_));
NAND_g _20328_ (.A(cpuregs_22[4]), .B(_00011_[2]), .Y(_14210_));
NAND_g _20329_ (.A(cpuregs_18[4]), .B(_11219_), .Y(_14211_));
AND_g _20330_ (.A(_11217_), .B(_14211_), .Y(_14212_));
NAND_g _20331_ (.A(_14210_), .B(_14212_), .Y(_14213_));
NAND_g _20332_ (.A(cpuregs_19[4]), .B(_11219_), .Y(_14214_));
NAND_g _20333_ (.A(cpuregs_23[4]), .B(_00011_[2]), .Y(_14215_));
AND_g _20334_ (.A(_00011_[0]), .B(_14215_), .Y(_14216_));
NAND_g _20335_ (.A(_14214_), .B(_14216_), .Y(_14217_));
AND_g _20336_ (.A(_14213_), .B(_14217_), .Y(_14218_));
NAND_g _20337_ (.A(_11220_), .B(_14218_), .Y(_14219_));
AND_g _20338_ (.A(_14209_), .B(_14219_), .Y(_14220_));
NAND_g _20339_ (.A(_00011_[1]), .B(_14220_), .Y(_14221_));
NAND_g _20340_ (.A(_11218_), .B(_14178_), .Y(_14222_));
AND_g _20341_ (.A(_00011_[4]), .B(_14222_), .Y(_14223_));
NAND_g _20342_ (.A(_14221_), .B(_14223_), .Y(_14224_));
NAND_g _20343_ (.A(cpuregs_6[4]), .B(_00011_[2]), .Y(_14225_));
NAND_g _20344_ (.A(cpuregs_2[4]), .B(_11219_), .Y(_14226_));
AND_g _20345_ (.A(_14225_), .B(_14226_), .Y(_14227_));
NAND_g _20346_ (.A(_11217_), .B(_14227_), .Y(_14228_));
NAND_g _20347_ (.A(cpuregs_7[4]), .B(_00011_[2]), .Y(_14229_));
NAND_g _20348_ (.A(cpuregs_3[4]), .B(_11219_), .Y(_14230_));
AND_g _20349_ (.A(_00011_[0]), .B(_14230_), .Y(_14231_));
NAND_g _20350_ (.A(_14229_), .B(_14231_), .Y(_14232_));
AND_g _20351_ (.A(_11220_), .B(_14232_), .Y(_14233_));
NAND_g _20352_ (.A(_14228_), .B(_14233_), .Y(_14234_));
NOR_g _20353_ (.A(cpuregs_11[4]), .B(_00011_[2]), .Y(_14235_));
NOT_g _20354_ (.A(_14235_), .Y(_14236_));
NAND_g _20355_ (.A(_11158_), .B(_00011_[2]), .Y(_14237_));
AND_g _20356_ (.A(_00011_[0]), .B(_14237_), .Y(_14238_));
NAND_g _20357_ (.A(_14236_), .B(_14238_), .Y(_14239_));
NOR_g _20358_ (.A(cpuregs_10[4]), .B(_00011_[2]), .Y(_14240_));
NOR_g _20359_ (.A(cpuregs_14[4]), .B(_11219_), .Y(_14241_));
NOR_g _20360_ (.A(_14240_), .B(_14241_), .Y(_14242_));
NAND_g _20361_ (.A(_11217_), .B(_14242_), .Y(_14243_));
NAND_g _20362_ (.A(_14239_), .B(_14243_), .Y(_14244_));
NAND_g _20363_ (.A(_00011_[3]), .B(_14244_), .Y(_14245_));
AND_g _20364_ (.A(_14234_), .B(_14245_), .Y(_14246_));
NAND_g _20365_ (.A(_00011_[1]), .B(_14246_), .Y(_14247_));
NAND_g _20366_ (.A(_11218_), .B(_14199_), .Y(_14248_));
AND_g _20367_ (.A(_14247_), .B(_14248_), .Y(_14249_));
NAND_g _20368_ (.A(_11221_), .B(_14249_), .Y(_14250_));
NAND_g _20369_ (.A(_14224_), .B(_14250_), .Y(_14251_));
AND_g _20370_ (.A(_13734_), .B(_14251_), .Y(_14252_));
AND_g _20371_ (.A(_13833_), .B(_14252_), .Y(_14253_));
NAND_g _20372_ (.A(_13833_), .B(_14252_), .Y(_14254_));
NAND_g _20373_ (.A(decoded_imm[4]), .B(_13830_), .Y(_14255_));
NAND_g _20374_ (.A(_14254_), .B(_14255_), .Y(_14256_));
NAND_g _20375_ (.A(_13409_), .B(_14256_), .Y(_14257_));
NAND_g _20376_ (.A(_13724_), .B(_14252_), .Y(_14258_));
NOT_g _20377_ (.A(_14258_), .Y(_14259_));
AND_g _20378_ (.A(_13727_), .B(_14258_), .Y(_14260_));
NAND_g _20379_ (.A(_14257_), .B(_14260_), .Y(_14261_));
AND_g _20380_ (.A(_14157_), .B(_14261_), .Y(_00507_));
NAND_g _20381_ (.A(_10985_), .B(_13728_), .Y(_14262_));
NAND_g _20382_ (.A(cpuregs_19[5]), .B(_11219_), .Y(_14263_));
NAND_g _20383_ (.A(cpuregs_23[5]), .B(_00011_[2]), .Y(_14264_));
AND_g _20384_ (.A(_00011_[0]), .B(_14264_), .Y(_14265_));
NAND_g _20385_ (.A(_14263_), .B(_14265_), .Y(_14266_));
NAND_g _20386_ (.A(cpuregs_18[5]), .B(_11219_), .Y(_14267_));
NAND_g _20387_ (.A(cpuregs_22[5]), .B(_00011_[2]), .Y(_14268_));
AND_g _20388_ (.A(_11217_), .B(_14268_), .Y(_14269_));
NAND_g _20389_ (.A(_14267_), .B(_14269_), .Y(_14270_));
AND_g _20390_ (.A(_11220_), .B(_14270_), .Y(_14271_));
NAND_g _20391_ (.A(_14266_), .B(_14271_), .Y(_14272_));
NAND_g _20392_ (.A(cpuregs_27[5]), .B(_11219_), .Y(_14273_));
NAND_g _20393_ (.A(cpuregs_31[5]), .B(_00011_[2]), .Y(_14274_));
AND_g _20394_ (.A(_00011_[0]), .B(_14274_), .Y(_14275_));
NAND_g _20395_ (.A(_14273_), .B(_14275_), .Y(_14276_));
NAND_g _20396_ (.A(cpuregs_26[5]), .B(_11219_), .Y(_14277_));
NAND_g _20397_ (.A(cpuregs_30[5]), .B(_00011_[2]), .Y(_14278_));
AND_g _20398_ (.A(_11217_), .B(_14278_), .Y(_14279_));
NAND_g _20399_ (.A(_14277_), .B(_14279_), .Y(_14280_));
AND_g _20400_ (.A(_00011_[3]), .B(_14280_), .Y(_14281_));
NAND_g _20401_ (.A(_14276_), .B(_14281_), .Y(_14282_));
NAND_g _20402_ (.A(_14272_), .B(_14282_), .Y(_14283_));
NAND_g _20403_ (.A(_00011_[1]), .B(_14283_), .Y(_14284_));
NOR_g _20404_ (.A(cpuregs_16[5]), .B(_00011_[2]), .Y(_14285_));
NOR_g _20405_ (.A(cpuregs_20[5]), .B(_11219_), .Y(_14286_));
NOR_g _20406_ (.A(_14285_), .B(_14286_), .Y(_14287_));
NOR_g _20407_ (.A(cpuregs_17[5]), .B(_00011_[2]), .Y(_14288_));
NAND_g _20408_ (.A(_11024_), .B(_00011_[2]), .Y(_14289_));
NOR_g _20409_ (.A(cpuregs_24[5]), .B(_00011_[2]), .Y(_14290_));
NOR_g _20410_ (.A(cpuregs_28[5]), .B(_11219_), .Y(_14291_));
NOR_g _20411_ (.A(_14290_), .B(_14291_), .Y(_14292_));
NOR_g _20412_ (.A(cpuregs_25[5]), .B(_00011_[2]), .Y(_14293_));
NAND_g _20413_ (.A(_10924_), .B(_00011_[2]), .Y(_14294_));
NAND_g _20414_ (.A(_11217_), .B(_14287_), .Y(_14295_));
NOR_g _20415_ (.A(_11217_), .B(_14288_), .Y(_14296_));
NAND_g _20416_ (.A(_14289_), .B(_14296_), .Y(_14297_));
AND_g _20417_ (.A(_14295_), .B(_14297_), .Y(_14298_));
NAND_g _20418_ (.A(_11220_), .B(_14298_), .Y(_14299_));
NOR_g _20419_ (.A(_11217_), .B(_14293_), .Y(_14300_));
NAND_g _20420_ (.A(_14294_), .B(_14300_), .Y(_14301_));
NAND_g _20421_ (.A(_11217_), .B(_14292_), .Y(_14302_));
AND_g _20422_ (.A(_14301_), .B(_14302_), .Y(_14303_));
NAND_g _20423_ (.A(_00011_[3]), .B(_14303_), .Y(_14304_));
AND_g _20424_ (.A(_14299_), .B(_14304_), .Y(_14305_));
NAND_g _20425_ (.A(_11218_), .B(_14305_), .Y(_14306_));
NAND_g _20426_ (.A(cpuregs_14[5]), .B(_11217_), .Y(_14307_));
NAND_g _20427_ (.A(cpuregs_15[5]), .B(_00011_[0]), .Y(_14308_));
NAND_g _20428_ (.A(_14307_), .B(_14308_), .Y(_14309_));
NAND_g _20429_ (.A(_00011_[2]), .B(_14309_), .Y(_14310_));
NAND_g _20430_ (.A(cpuregs_10[5]), .B(_11217_), .Y(_14311_));
NAND_g _20431_ (.A(cpuregs_11[5]), .B(_00011_[0]), .Y(_14312_));
NAND_g _20432_ (.A(_14311_), .B(_14312_), .Y(_14313_));
NAND_g _20433_ (.A(_11219_), .B(_14313_), .Y(_14314_));
NAND_g _20434_ (.A(_14310_), .B(_14314_), .Y(_14315_));
NAND_g _20435_ (.A(_00011_[3]), .B(_14315_), .Y(_14316_));
NAND_g _20436_ (.A(cpuregs_6[5]), .B(_11217_), .Y(_14317_));
NAND_g _20437_ (.A(cpuregs_7[5]), .B(_00011_[0]), .Y(_14318_));
NAND_g _20438_ (.A(_14317_), .B(_14318_), .Y(_14319_));
NAND_g _20439_ (.A(_00011_[2]), .B(_14319_), .Y(_14320_));
NAND_g _20440_ (.A(cpuregs_2[5]), .B(_11217_), .Y(_14321_));
NAND_g _20441_ (.A(cpuregs_3[5]), .B(_00011_[0]), .Y(_14322_));
NAND_g _20442_ (.A(_14321_), .B(_14322_), .Y(_14323_));
NAND_g _20443_ (.A(_11219_), .B(_14323_), .Y(_14324_));
NAND_g _20444_ (.A(_14320_), .B(_14324_), .Y(_14325_));
NAND_g _20445_ (.A(_11220_), .B(_14325_), .Y(_14326_));
NAND_g _20446_ (.A(_14316_), .B(_14326_), .Y(_14327_));
NAND_g _20447_ (.A(_00011_[1]), .B(_14327_), .Y(_14328_));
NOR_g _20448_ (.A(cpuregs_9[5]), .B(_00011_[2]), .Y(_14329_));
NOT_g _20449_ (.A(_14329_), .Y(_14330_));
NAND_g _20450_ (.A(_11142_), .B(_00011_[2]), .Y(_14331_));
AND_g _20451_ (.A(_00011_[0]), .B(_14331_), .Y(_14332_));
NAND_g _20452_ (.A(_14330_), .B(_14332_), .Y(_14333_));
NOR_g _20453_ (.A(cpuregs_8[5]), .B(_00011_[2]), .Y(_14334_));
NOR_g _20454_ (.A(cpuregs_12[5]), .B(_11219_), .Y(_14335_));
NOR_g _20455_ (.A(_14334_), .B(_14335_), .Y(_14336_));
NAND_g _20456_ (.A(_11217_), .B(_14336_), .Y(_14337_));
NAND_g _20457_ (.A(_14333_), .B(_14337_), .Y(_14338_));
NAND_g _20458_ (.A(_00011_[3]), .B(_14338_), .Y(_14339_));
NAND_g _20459_ (.A(cpuregs_4[5]), .B(_00011_[2]), .Y(_14340_));
NAND_g _20460_ (.A(cpuregs_0[5]), .B(_11219_), .Y(_14341_));
AND_g _20461_ (.A(_14340_), .B(_14341_), .Y(_14342_));
NAND_g _20462_ (.A(_11217_), .B(_14342_), .Y(_14343_));
NAND_g _20463_ (.A(cpuregs_5[5]), .B(_00011_[2]), .Y(_14344_));
NAND_g _20464_ (.A(cpuregs_1[5]), .B(_11219_), .Y(_14345_));
AND_g _20465_ (.A(_00011_[0]), .B(_14345_), .Y(_14346_));
NAND_g _20466_ (.A(_14344_), .B(_14346_), .Y(_14347_));
AND_g _20467_ (.A(_11220_), .B(_14347_), .Y(_14348_));
NAND_g _20468_ (.A(_14343_), .B(_14348_), .Y(_14349_));
NAND_g _20469_ (.A(_14339_), .B(_14349_), .Y(_14350_));
NAND_g _20470_ (.A(_11218_), .B(_14350_), .Y(_14351_));
AND_g _20471_ (.A(_14328_), .B(_14351_), .Y(_14352_));
AND_g _20472_ (.A(_00011_[4]), .B(_14284_), .Y(_14353_));
NAND_g _20473_ (.A(_14306_), .B(_14353_), .Y(_14354_));
NAND_g _20474_ (.A(_11221_), .B(_14352_), .Y(_14355_));
AND_g _20475_ (.A(_14354_), .B(_14355_), .Y(_14356_));
AND_g _20476_ (.A(_13734_), .B(_14356_), .Y(_14357_));
NAND_g _20477_ (.A(_13725_), .B(_13940_), .Y(_14358_));
NAND_g _20478_ (.A(_14357_), .B(_14358_), .Y(_14359_));
AND_g _20479_ (.A(decoded_imm[5]), .B(_13830_), .Y(_14360_));
NAND_g _20480_ (.A(_13409_), .B(_14360_), .Y(_14361_));
AND_g _20481_ (.A(_13727_), .B(_14361_), .Y(_14362_));
NAND_g _20482_ (.A(_14359_), .B(_14362_), .Y(_14363_));
AND_g _20483_ (.A(_14262_), .B(_14363_), .Y(_00508_));
NAND_g _20484_ (.A(_10986_), .B(_13728_), .Y(_14364_));
NAND_g _20485_ (.A(cpuregs_31[6]), .B(_00011_[1]), .Y(_14365_));
NAND_g _20486_ (.A(cpuregs_29[6]), .B(_11218_), .Y(_14366_));
NAND_g _20487_ (.A(_14365_), .B(_14366_), .Y(_14367_));
NAND_g _20488_ (.A(_00011_[2]), .B(_14367_), .Y(_14368_));
NAND_g _20489_ (.A(cpuregs_27[6]), .B(_00011_[1]), .Y(_14369_));
NAND_g _20490_ (.A(cpuregs_25[6]), .B(_11218_), .Y(_14370_));
NAND_g _20491_ (.A(_14369_), .B(_14370_), .Y(_14371_));
NAND_g _20492_ (.A(_11219_), .B(_14371_), .Y(_14372_));
NAND_g _20493_ (.A(_14368_), .B(_14372_), .Y(_14373_));
NAND_g _20494_ (.A(_00011_[0]), .B(_14373_), .Y(_14374_));
NAND_g _20495_ (.A(cpuregs_30[6]), .B(_00011_[1]), .Y(_14375_));
NAND_g _20496_ (.A(cpuregs_28[6]), .B(_11218_), .Y(_14376_));
NAND_g _20497_ (.A(_14375_), .B(_14376_), .Y(_14377_));
NAND_g _20498_ (.A(_00011_[2]), .B(_14377_), .Y(_14378_));
NAND_g _20499_ (.A(cpuregs_26[6]), .B(_00011_[1]), .Y(_14379_));
NAND_g _20500_ (.A(cpuregs_24[6]), .B(_11218_), .Y(_14380_));
NAND_g _20501_ (.A(_14379_), .B(_14380_), .Y(_14381_));
NAND_g _20502_ (.A(_11219_), .B(_14381_), .Y(_14382_));
NAND_g _20503_ (.A(_14378_), .B(_14382_), .Y(_14383_));
AND_g _20504_ (.A(_11217_), .B(_14383_), .Y(_14384_));
NOT_g _20505_ (.A(_14384_), .Y(_14385_));
NAND_g _20506_ (.A(_14374_), .B(_14385_), .Y(_14386_));
NAND_g _20507_ (.A(_00011_[3]), .B(_14386_), .Y(_14387_));
NOR_g _20508_ (.A(cpuregs_18[6]), .B(_00011_[2]), .Y(_14388_));
NOR_g _20509_ (.A(cpuregs_22[6]), .B(_11219_), .Y(_14389_));
NOR_g _20510_ (.A(_14388_), .B(_14389_), .Y(_14390_));
NOR_g _20511_ (.A(cpuregs_16[6]), .B(_00011_[2]), .Y(_14391_));
AND_g _20512_ (.A(_11194_), .B(_00011_[2]), .Y(_14392_));
NOR_g _20513_ (.A(_14391_), .B(_14392_), .Y(_14393_));
NAND_g _20514_ (.A(_11179_), .B(_00011_[2]), .Y(_14394_));
NOR_g _20515_ (.A(cpuregs_19[6]), .B(_00011_[2]), .Y(_14395_));
NOR_g _20516_ (.A(cpuregs_17[6]), .B(_00011_[2]), .Y(_14396_));
NAND_g _20517_ (.A(_11025_), .B(_00011_[2]), .Y(_14397_));
NOR_g _20518_ (.A(_11217_), .B(_14395_), .Y(_14398_));
NAND_g _20519_ (.A(_14394_), .B(_14398_), .Y(_14399_));
NAND_g _20520_ (.A(_11217_), .B(_14390_), .Y(_14400_));
AND_g _20521_ (.A(_14399_), .B(_14400_), .Y(_14401_));
NAND_g _20522_ (.A(_00011_[1]), .B(_14401_), .Y(_14402_));
NOR_g _20523_ (.A(_11217_), .B(_14396_), .Y(_14403_));
NAND_g _20524_ (.A(_14397_), .B(_14403_), .Y(_14404_));
NAND_g _20525_ (.A(_11217_), .B(_14393_), .Y(_14405_));
AND_g _20526_ (.A(_14404_), .B(_14405_), .Y(_14406_));
NAND_g _20527_ (.A(_11218_), .B(_14406_), .Y(_14407_));
AND_g _20528_ (.A(_14402_), .B(_14407_), .Y(_14408_));
NAND_g _20529_ (.A(_11220_), .B(_14408_), .Y(_14409_));
AND_g _20530_ (.A(_14387_), .B(_14409_), .Y(_14410_));
NAND_g _20531_ (.A(cpuregs_13[6]), .B(_11218_), .Y(_14411_));
NAND_g _20532_ (.A(cpuregs_15[6]), .B(_00011_[1]), .Y(_14412_));
AND_g _20533_ (.A(_00011_[2]), .B(_14412_), .Y(_14413_));
NAND_g _20534_ (.A(_14411_), .B(_14413_), .Y(_14414_));
NAND_g _20535_ (.A(cpuregs_9[6]), .B(_11218_), .Y(_14415_));
NAND_g _20536_ (.A(cpuregs_11[6]), .B(_00011_[1]), .Y(_14416_));
AND_g _20537_ (.A(_11219_), .B(_14416_), .Y(_14417_));
NAND_g _20538_ (.A(_14415_), .B(_14417_), .Y(_14418_));
AND_g _20539_ (.A(_00011_[0]), .B(_14418_), .Y(_14419_));
NAND_g _20540_ (.A(_14414_), .B(_14419_), .Y(_14420_));
NAND_g _20541_ (.A(cpuregs_12[6]), .B(_11218_), .Y(_14421_));
NAND_g _20542_ (.A(cpuregs_14[6]), .B(_00011_[1]), .Y(_14422_));
AND_g _20543_ (.A(_00011_[2]), .B(_14422_), .Y(_14423_));
NAND_g _20544_ (.A(_14421_), .B(_14423_), .Y(_14424_));
NAND_g _20545_ (.A(cpuregs_8[6]), .B(_11218_), .Y(_14425_));
NAND_g _20546_ (.A(cpuregs_10[6]), .B(_00011_[1]), .Y(_14426_));
AND_g _20547_ (.A(_11219_), .B(_14426_), .Y(_14427_));
NAND_g _20548_ (.A(_14425_), .B(_14427_), .Y(_14428_));
AND_g _20549_ (.A(_11217_), .B(_14428_), .Y(_14429_));
NAND_g _20550_ (.A(_14424_), .B(_14429_), .Y(_14430_));
NAND_g _20551_ (.A(_14420_), .B(_14430_), .Y(_14431_));
NAND_g _20552_ (.A(_00011_[3]), .B(_14431_), .Y(_14432_));
NAND_g _20553_ (.A(_10939_), .B(_00011_[2]), .Y(_14433_));
NOR_g _20554_ (.A(cpuregs_2[6]), .B(_00011_[2]), .Y(_14434_));
NOR_g _20555_ (.A(_00011_[0]), .B(_14434_), .Y(_14435_));
NAND_g _20556_ (.A(_14433_), .B(_14435_), .Y(_14436_));
NAND_g _20557_ (.A(_11125_), .B(_00011_[2]), .Y(_14437_));
NOR_g _20558_ (.A(cpuregs_3[6]), .B(_00011_[2]), .Y(_14438_));
NOR_g _20559_ (.A(_11217_), .B(_14438_), .Y(_14439_));
NAND_g _20560_ (.A(_14437_), .B(_14439_), .Y(_14440_));
AND_g _20561_ (.A(_14436_), .B(_14440_), .Y(_14441_));
NAND_g _20562_ (.A(_10951_), .B(_00011_[2]), .Y(_14442_));
NOR_g _20563_ (.A(cpuregs_0[6]), .B(_00011_[2]), .Y(_14443_));
NOR_g _20564_ (.A(_00011_[0]), .B(_14443_), .Y(_14444_));
NAND_g _20565_ (.A(_14442_), .B(_14444_), .Y(_14445_));
NAND_g _20566_ (.A(_11109_), .B(_00011_[2]), .Y(_14446_));
NOR_g _20567_ (.A(cpuregs_1[6]), .B(_00011_[2]), .Y(_14447_));
NOR_g _20568_ (.A(_11217_), .B(_14447_), .Y(_14448_));
NAND_g _20569_ (.A(_14446_), .B(_14448_), .Y(_14449_));
AND_g _20570_ (.A(_14445_), .B(_14449_), .Y(_14450_));
NAND_g _20571_ (.A(_00011_[1]), .B(_14441_), .Y(_14451_));
NAND_g _20572_ (.A(_11218_), .B(_14450_), .Y(_14452_));
AND_g _20573_ (.A(_14451_), .B(_14452_), .Y(_14453_));
NAND_g _20574_ (.A(_11220_), .B(_14453_), .Y(_14454_));
AND_g _20575_ (.A(_14432_), .B(_14454_), .Y(_14455_));
NAND_g _20576_ (.A(_00011_[4]), .B(_14410_), .Y(_14456_));
NAND_g _20577_ (.A(_11221_), .B(_14455_), .Y(_14457_));
AND_g _20578_ (.A(_13734_), .B(_14457_), .Y(_14458_));
AND_g _20579_ (.A(_14456_), .B(_14458_), .Y(_14459_));
NAND_g _20580_ (.A(_14358_), .B(_14459_), .Y(_14460_));
AND_g _20581_ (.A(decoded_imm[6]), .B(_13830_), .Y(_14461_));
NAND_g _20582_ (.A(_13409_), .B(_14461_), .Y(_14462_));
AND_g _20583_ (.A(_13727_), .B(_14462_), .Y(_14463_));
NAND_g _20584_ (.A(_14460_), .B(_14463_), .Y(_14464_));
AND_g _20585_ (.A(_14364_), .B(_14464_), .Y(_00509_));
NAND_g _20586_ (.A(_10987_), .B(_13728_), .Y(_14465_));
NAND_g _20587_ (.A(cpuregs_29[7]), .B(_00011_[2]), .Y(_14466_));
NAND_g _20588_ (.A(cpuregs_25[7]), .B(_11219_), .Y(_14467_));
AND_g _20589_ (.A(_00011_[0]), .B(_14467_), .Y(_14468_));
NAND_g _20590_ (.A(_14466_), .B(_14468_), .Y(_14469_));
NAND_g _20591_ (.A(cpuregs_24[7]), .B(_11219_), .Y(_14470_));
NAND_g _20592_ (.A(cpuregs_28[7]), .B(_00011_[2]), .Y(_14471_));
AND_g _20593_ (.A(_11217_), .B(_14471_), .Y(_14472_));
NAND_g _20594_ (.A(_14470_), .B(_14472_), .Y(_14473_));
AND_g _20595_ (.A(_11218_), .B(_14473_), .Y(_14474_));
NAND_g _20596_ (.A(_14469_), .B(_14474_), .Y(_14475_));
NAND_g _20597_ (.A(cpuregs_27[7]), .B(_11219_), .Y(_14476_));
NAND_g _20598_ (.A(cpuregs_31[7]), .B(_00011_[2]), .Y(_14477_));
AND_g _20599_ (.A(_00011_[0]), .B(_14477_), .Y(_14478_));
NAND_g _20600_ (.A(_14476_), .B(_14478_), .Y(_14479_));
NAND_g _20601_ (.A(cpuregs_26[7]), .B(_11219_), .Y(_14480_));
NAND_g _20602_ (.A(cpuregs_30[7]), .B(_00011_[2]), .Y(_14481_));
AND_g _20603_ (.A(_11217_), .B(_14481_), .Y(_14482_));
NAND_g _20604_ (.A(_14480_), .B(_14482_), .Y(_14483_));
AND_g _20605_ (.A(_00011_[1]), .B(_14483_), .Y(_14484_));
NAND_g _20606_ (.A(_14479_), .B(_14484_), .Y(_14485_));
NAND_g _20607_ (.A(_14475_), .B(_14485_), .Y(_14486_));
NAND_g _20608_ (.A(_00011_[4]), .B(_14486_), .Y(_14487_));
NAND_g _20609_ (.A(cpuregs_14[7]), .B(_11217_), .Y(_14488_));
NAND_g _20610_ (.A(cpuregs_15[7]), .B(_00011_[0]), .Y(_14489_));
NAND_g _20611_ (.A(_14488_), .B(_14489_), .Y(_14490_));
NAND_g _20612_ (.A(_00011_[2]), .B(_14490_), .Y(_14491_));
NAND_g _20613_ (.A(cpuregs_10[7]), .B(_11217_), .Y(_14492_));
NAND_g _20614_ (.A(cpuregs_11[7]), .B(_00011_[0]), .Y(_14493_));
NAND_g _20615_ (.A(_14492_), .B(_14493_), .Y(_14494_));
NAND_g _20616_ (.A(_11219_), .B(_14494_), .Y(_14495_));
NAND_g _20617_ (.A(_14491_), .B(_14495_), .Y(_14496_));
NAND_g _20618_ (.A(_00011_[1]), .B(_14496_), .Y(_14497_));
NAND_g _20619_ (.A(cpuregs_12[7]), .B(_11217_), .Y(_14498_));
NAND_g _20620_ (.A(cpuregs_13[7]), .B(_00011_[0]), .Y(_14499_));
NAND_g _20621_ (.A(_14498_), .B(_14499_), .Y(_14500_));
NAND_g _20622_ (.A(_00011_[2]), .B(_14500_), .Y(_14501_));
NAND_g _20623_ (.A(cpuregs_8[7]), .B(_11217_), .Y(_14502_));
NAND_g _20624_ (.A(cpuregs_9[7]), .B(_00011_[0]), .Y(_14503_));
NAND_g _20625_ (.A(_14502_), .B(_14503_), .Y(_14504_));
NAND_g _20626_ (.A(_11219_), .B(_14504_), .Y(_14505_));
NAND_g _20627_ (.A(_14501_), .B(_14505_), .Y(_14506_));
NAND_g _20628_ (.A(_11218_), .B(_14506_), .Y(_14507_));
NAND_g _20629_ (.A(_14497_), .B(_14507_), .Y(_14508_));
AND_g _20630_ (.A(_11221_), .B(_14508_), .Y(_14509_));
NOT_g _20631_ (.A(_14509_), .Y(_14510_));
NAND_g _20632_ (.A(_14487_), .B(_14510_), .Y(_14511_));
NAND_g _20633_ (.A(_00011_[3]), .B(_14511_), .Y(_14512_));
NAND_g _20634_ (.A(cpuregs_1[7]), .B(_11219_), .Y(_14513_));
NAND_g _20635_ (.A(cpuregs_5[7]), .B(_00011_[2]), .Y(_14514_));
AND_g _20636_ (.A(_00011_[0]), .B(_14514_), .Y(_14515_));
NAND_g _20637_ (.A(_14513_), .B(_14515_), .Y(_14516_));
NAND_g _20638_ (.A(cpuregs_0[7]), .B(_11219_), .Y(_14517_));
NAND_g _20639_ (.A(cpuregs_4[7]), .B(_00011_[2]), .Y(_14518_));
AND_g _20640_ (.A(_11217_), .B(_14518_), .Y(_14519_));
NAND_g _20641_ (.A(_14517_), .B(_14519_), .Y(_14520_));
AND_g _20642_ (.A(_11218_), .B(_14520_), .Y(_14521_));
NAND_g _20643_ (.A(_14516_), .B(_14521_), .Y(_14522_));
NAND_g _20644_ (.A(cpuregs_3[7]), .B(_11219_), .Y(_14523_));
NAND_g _20645_ (.A(cpuregs_7[7]), .B(_00011_[2]), .Y(_14524_));
AND_g _20646_ (.A(_00011_[0]), .B(_14524_), .Y(_14525_));
NAND_g _20647_ (.A(_14523_), .B(_14525_), .Y(_14526_));
NAND_g _20648_ (.A(cpuregs_2[7]), .B(_11219_), .Y(_14527_));
NAND_g _20649_ (.A(cpuregs_6[7]), .B(_00011_[2]), .Y(_14528_));
AND_g _20650_ (.A(_11217_), .B(_14528_), .Y(_14529_));
NAND_g _20651_ (.A(_14527_), .B(_14529_), .Y(_14530_));
AND_g _20652_ (.A(_00011_[1]), .B(_14530_), .Y(_14531_));
NAND_g _20653_ (.A(_14526_), .B(_14531_), .Y(_14532_));
NAND_g _20654_ (.A(_14522_), .B(_14532_), .Y(_14533_));
NAND_g _20655_ (.A(_11221_), .B(_14533_), .Y(_14534_));
NAND_g _20656_ (.A(cpuregs_19[7]), .B(_00011_[1]), .Y(_14535_));
NAND_g _20657_ (.A(cpuregs_17[7]), .B(_11218_), .Y(_14536_));
NAND_g _20658_ (.A(_14535_), .B(_14536_), .Y(_14537_));
NAND_g _20659_ (.A(_11219_), .B(_14537_), .Y(_14538_));
NAND_g _20660_ (.A(cpuregs_23[7]), .B(_00011_[1]), .Y(_14539_));
NAND_g _20661_ (.A(cpuregs_21[7]), .B(_11218_), .Y(_14540_));
NAND_g _20662_ (.A(_14539_), .B(_14540_), .Y(_14541_));
NAND_g _20663_ (.A(_00011_[2]), .B(_14541_), .Y(_14542_));
AND_g _20664_ (.A(_00011_[0]), .B(_14542_), .Y(_14543_));
NAND_g _20665_ (.A(_14538_), .B(_14543_), .Y(_14544_));
NAND_g _20666_ (.A(cpuregs_18[7]), .B(_00011_[1]), .Y(_14545_));
NAND_g _20667_ (.A(cpuregs_16[7]), .B(_11218_), .Y(_14546_));
NAND_g _20668_ (.A(_14545_), .B(_14546_), .Y(_14547_));
NAND_g _20669_ (.A(_11219_), .B(_14547_), .Y(_14548_));
NAND_g _20670_ (.A(cpuregs_22[7]), .B(_00011_[1]), .Y(_14549_));
NAND_g _20671_ (.A(cpuregs_20[7]), .B(_11218_), .Y(_14550_));
NAND_g _20672_ (.A(_14549_), .B(_14550_), .Y(_14551_));
NAND_g _20673_ (.A(_00011_[2]), .B(_14551_), .Y(_14552_));
AND_g _20674_ (.A(_11217_), .B(_14552_), .Y(_14553_));
NAND_g _20675_ (.A(_14548_), .B(_14553_), .Y(_14554_));
AND_g _20676_ (.A(_00011_[4]), .B(_14554_), .Y(_14555_));
NAND_g _20677_ (.A(_14544_), .B(_14555_), .Y(_14556_));
NAND_g _20678_ (.A(_14534_), .B(_14556_), .Y(_14557_));
NAND_g _20679_ (.A(_11220_), .B(_14557_), .Y(_14558_));
NAND_g _20680_ (.A(_14512_), .B(_14558_), .Y(_14559_));
AND_g _20681_ (.A(_13734_), .B(_14559_), .Y(_14560_));
NAND_g _20682_ (.A(_14358_), .B(_14560_), .Y(_14561_));
AND_g _20683_ (.A(decoded_imm[7]), .B(_13830_), .Y(_14562_));
NAND_g _20684_ (.A(_13409_), .B(_14562_), .Y(_14563_));
AND_g _20685_ (.A(_13727_), .B(_14563_), .Y(_14564_));
NAND_g _20686_ (.A(_14561_), .B(_14564_), .Y(_14565_));
AND_g _20687_ (.A(_14465_), .B(_14565_), .Y(_00510_));
NAND_g _20688_ (.A(_10988_), .B(_13728_), .Y(_14566_));
NAND_g _20689_ (.A(cpuregs_19[8]), .B(_11219_), .Y(_14567_));
NAND_g _20690_ (.A(cpuregs_23[8]), .B(_00011_[2]), .Y(_14568_));
AND_g _20691_ (.A(_00011_[0]), .B(_14568_), .Y(_14569_));
NAND_g _20692_ (.A(_14567_), .B(_14569_), .Y(_14570_));
NAND_g _20693_ (.A(cpuregs_18[8]), .B(_11219_), .Y(_14571_));
NAND_g _20694_ (.A(cpuregs_22[8]), .B(_00011_[2]), .Y(_14572_));
AND_g _20695_ (.A(_11217_), .B(_14572_), .Y(_14573_));
NAND_g _20696_ (.A(_14571_), .B(_14573_), .Y(_14574_));
AND_g _20697_ (.A(_11220_), .B(_14574_), .Y(_14575_));
NAND_g _20698_ (.A(_14570_), .B(_14575_), .Y(_14576_));
NAND_g _20699_ (.A(cpuregs_27[8]), .B(_11219_), .Y(_14577_));
NAND_g _20700_ (.A(cpuregs_31[8]), .B(_00011_[2]), .Y(_14578_));
AND_g _20701_ (.A(_00011_[0]), .B(_14578_), .Y(_14579_));
NAND_g _20702_ (.A(_14577_), .B(_14579_), .Y(_14580_));
NAND_g _20703_ (.A(cpuregs_26[8]), .B(_11219_), .Y(_14581_));
NAND_g _20704_ (.A(cpuregs_30[8]), .B(_00011_[2]), .Y(_14582_));
AND_g _20705_ (.A(_11217_), .B(_14582_), .Y(_14583_));
NAND_g _20706_ (.A(_14581_), .B(_14583_), .Y(_14584_));
AND_g _20707_ (.A(_00011_[3]), .B(_14584_), .Y(_14585_));
NAND_g _20708_ (.A(_14580_), .B(_14585_), .Y(_14586_));
NAND_g _20709_ (.A(_14576_), .B(_14586_), .Y(_14587_));
NAND_g _20710_ (.A(_00011_[1]), .B(_14587_), .Y(_14588_));
NAND_g _20711_ (.A(cpuregs_21[8]), .B(_00011_[2]), .Y(_14589_));
NAND_g _20712_ (.A(cpuregs_17[8]), .B(_11219_), .Y(_14590_));
AND_g _20713_ (.A(_00011_[0]), .B(_14590_), .Y(_14591_));
NAND_g _20714_ (.A(_14589_), .B(_14591_), .Y(_14592_));
NAND_g _20715_ (.A(cpuregs_20[8]), .B(_00011_[2]), .Y(_14593_));
NAND_g _20716_ (.A(cpuregs_16[8]), .B(_11219_), .Y(_14594_));
AND_g _20717_ (.A(_11217_), .B(_14594_), .Y(_14595_));
NAND_g _20718_ (.A(_14593_), .B(_14595_), .Y(_14596_));
AND_g _20719_ (.A(_11220_), .B(_14596_), .Y(_14597_));
NAND_g _20720_ (.A(_14592_), .B(_14597_), .Y(_14598_));
NAND_g _20721_ (.A(cpuregs_25[8]), .B(_11219_), .Y(_14599_));
NAND_g _20722_ (.A(cpuregs_29[8]), .B(_00011_[2]), .Y(_14600_));
AND_g _20723_ (.A(_00011_[0]), .B(_14600_), .Y(_14601_));
NAND_g _20724_ (.A(_14599_), .B(_14601_), .Y(_14602_));
NAND_g _20725_ (.A(cpuregs_24[8]), .B(_11219_), .Y(_14603_));
NAND_g _20726_ (.A(cpuregs_28[8]), .B(_00011_[2]), .Y(_14604_));
AND_g _20727_ (.A(_11217_), .B(_14604_), .Y(_14605_));
NAND_g _20728_ (.A(_14603_), .B(_14605_), .Y(_14606_));
AND_g _20729_ (.A(_00011_[3]), .B(_14606_), .Y(_14607_));
NAND_g _20730_ (.A(_14602_), .B(_14607_), .Y(_14608_));
NAND_g _20731_ (.A(_14598_), .B(_14608_), .Y(_14609_));
NAND_g _20732_ (.A(_11218_), .B(_14609_), .Y(_14610_));
NAND_g _20733_ (.A(_14588_), .B(_14610_), .Y(_14611_));
NAND_g _20734_ (.A(_00011_[4]), .B(_14611_), .Y(_14612_));
NAND_g _20735_ (.A(cpuregs_6[8]), .B(_00011_[2]), .Y(_14613_));
NAND_g _20736_ (.A(cpuregs_2[8]), .B(_11219_), .Y(_14614_));
AND_g _20737_ (.A(_14613_), .B(_14614_), .Y(_14615_));
NAND_g _20738_ (.A(_11217_), .B(_14615_), .Y(_14616_));
NAND_g _20739_ (.A(cpuregs_7[8]), .B(_00011_[2]), .Y(_14617_));
NAND_g _20740_ (.A(cpuregs_3[8]), .B(_11219_), .Y(_14618_));
AND_g _20741_ (.A(_00011_[0]), .B(_14618_), .Y(_14619_));
NAND_g _20742_ (.A(_14617_), .B(_14619_), .Y(_14620_));
AND_g _20743_ (.A(_11220_), .B(_14620_), .Y(_14621_));
NAND_g _20744_ (.A(_14616_), .B(_14621_), .Y(_14622_));
NOR_g _20745_ (.A(cpuregs_10[8]), .B(_00011_[2]), .Y(_14623_));
AND_g _20746_ (.A(_11102_), .B(_00011_[2]), .Y(_14624_));
NOR_g _20747_ (.A(_14623_), .B(_14624_), .Y(_14625_));
NOR_g _20748_ (.A(cpuregs_11[8]), .B(_00011_[2]), .Y(_14626_));
NOT_g _20749_ (.A(_14626_), .Y(_14627_));
NAND_g _20750_ (.A(_11159_), .B(_00011_[2]), .Y(_14628_));
AND_g _20751_ (.A(_00011_[0]), .B(_14628_), .Y(_14629_));
NAND_g _20752_ (.A(_14627_), .B(_14629_), .Y(_14630_));
NAND_g _20753_ (.A(_11217_), .B(_14625_), .Y(_14631_));
NAND_g _20754_ (.A(_14630_), .B(_14631_), .Y(_14632_));
NAND_g _20755_ (.A(_00011_[3]), .B(_14632_), .Y(_14633_));
AND_g _20756_ (.A(_14622_), .B(_14633_), .Y(_14634_));
NAND_g _20757_ (.A(cpuregs_4[8]), .B(_00011_[2]), .Y(_14635_));
NAND_g _20758_ (.A(cpuregs_0[8]), .B(_11219_), .Y(_14636_));
AND_g _20759_ (.A(_11217_), .B(_14636_), .Y(_14637_));
NAND_g _20760_ (.A(_14635_), .B(_14637_), .Y(_14638_));
NAND_g _20761_ (.A(cpuregs_1[8]), .B(_11219_), .Y(_14639_));
NAND_g _20762_ (.A(cpuregs_5[8]), .B(_00011_[2]), .Y(_14640_));
AND_g _20763_ (.A(_00011_[0]), .B(_14640_), .Y(_14641_));
NAND_g _20764_ (.A(_14639_), .B(_14641_), .Y(_14642_));
NOR_g _20765_ (.A(cpuregs_9[8]), .B(_00011_[2]), .Y(_14643_));
NAND_g _20766_ (.A(_11144_), .B(_00011_[2]), .Y(_14644_));
NOR_g _20767_ (.A(cpuregs_8[8]), .B(_00011_[2]), .Y(_14645_));
NOR_g _20768_ (.A(cpuregs_12[8]), .B(_11219_), .Y(_14646_));
NOR_g _20769_ (.A(_14645_), .B(_14646_), .Y(_14647_));
NAND_g _20770_ (.A(_14638_), .B(_14642_), .Y(_14648_));
NAND_g _20771_ (.A(_11220_), .B(_14648_), .Y(_14649_));
NAND_g _20772_ (.A(_11217_), .B(_14647_), .Y(_14650_));
NOR_g _20773_ (.A(_11217_), .B(_14643_), .Y(_14651_));
NAND_g _20774_ (.A(_14644_), .B(_14651_), .Y(_14652_));
AND_g _20775_ (.A(_00011_[3]), .B(_14652_), .Y(_14653_));
NAND_g _20776_ (.A(_14650_), .B(_14653_), .Y(_14654_));
NAND_g _20777_ (.A(_14649_), .B(_14654_), .Y(_14655_));
NAND_g _20778_ (.A(_11218_), .B(_14655_), .Y(_14656_));
NAND_g _20779_ (.A(_00011_[1]), .B(_14634_), .Y(_14657_));
AND_g _20780_ (.A(_14656_), .B(_14657_), .Y(_14658_));
NAND_g _20781_ (.A(_11221_), .B(_14658_), .Y(_14659_));
NAND_g _20782_ (.A(_14612_), .B(_14659_), .Y(_14660_));
AND_g _20783_ (.A(_13734_), .B(_14660_), .Y(_14661_));
NAND_g _20784_ (.A(_14358_), .B(_14661_), .Y(_14662_));
AND_g _20785_ (.A(decoded_imm[8]), .B(_13830_), .Y(_14663_));
NAND_g _20786_ (.A(_13409_), .B(_14663_), .Y(_14664_));
AND_g _20787_ (.A(_13727_), .B(_14664_), .Y(_14665_));
NAND_g _20788_ (.A(_14662_), .B(_14665_), .Y(_14666_));
AND_g _20789_ (.A(_14566_), .B(_14666_), .Y(_00511_));
NAND_g _20790_ (.A(_10989_), .B(_13728_), .Y(_14667_));
NAND_g _20791_ (.A(cpuregs_19[9]), .B(_11219_), .Y(_14668_));
NAND_g _20792_ (.A(cpuregs_23[9]), .B(_00011_[2]), .Y(_14669_));
AND_g _20793_ (.A(_00011_[0]), .B(_14669_), .Y(_14670_));
NAND_g _20794_ (.A(_14668_), .B(_14670_), .Y(_14671_));
NAND_g _20795_ (.A(cpuregs_18[9]), .B(_11219_), .Y(_14672_));
NAND_g _20796_ (.A(cpuregs_22[9]), .B(_00011_[2]), .Y(_14673_));
AND_g _20797_ (.A(_11217_), .B(_14673_), .Y(_14674_));
NAND_g _20798_ (.A(_14672_), .B(_14674_), .Y(_14675_));
AND_g _20799_ (.A(_11220_), .B(_14675_), .Y(_14676_));
NAND_g _20800_ (.A(_14671_), .B(_14676_), .Y(_14677_));
NAND_g _20801_ (.A(cpuregs_27[9]), .B(_11219_), .Y(_14678_));
NAND_g _20802_ (.A(cpuregs_31[9]), .B(_00011_[2]), .Y(_14679_));
AND_g _20803_ (.A(_00011_[0]), .B(_14679_), .Y(_14680_));
NAND_g _20804_ (.A(_14678_), .B(_14680_), .Y(_14681_));
NAND_g _20805_ (.A(cpuregs_26[9]), .B(_11219_), .Y(_14682_));
NAND_g _20806_ (.A(cpuregs_30[9]), .B(_00011_[2]), .Y(_14683_));
AND_g _20807_ (.A(_11217_), .B(_14683_), .Y(_14684_));
NAND_g _20808_ (.A(_14682_), .B(_14684_), .Y(_14685_));
AND_g _20809_ (.A(_00011_[3]), .B(_14685_), .Y(_14686_));
NAND_g _20810_ (.A(_14681_), .B(_14686_), .Y(_14687_));
NAND_g _20811_ (.A(_14677_), .B(_14687_), .Y(_14688_));
NAND_g _20812_ (.A(_00011_[1]), .B(_14688_), .Y(_14689_));
NAND_g _20813_ (.A(cpuregs_21[9]), .B(_00011_[2]), .Y(_14690_));
NAND_g _20814_ (.A(cpuregs_17[9]), .B(_11219_), .Y(_14691_));
AND_g _20815_ (.A(_00011_[0]), .B(_14691_), .Y(_14692_));
NAND_g _20816_ (.A(_14690_), .B(_14692_), .Y(_14693_));
NAND_g _20817_ (.A(cpuregs_20[9]), .B(_00011_[2]), .Y(_14694_));
NAND_g _20818_ (.A(cpuregs_16[9]), .B(_11219_), .Y(_14695_));
AND_g _20819_ (.A(_11217_), .B(_14695_), .Y(_14696_));
NAND_g _20820_ (.A(_14694_), .B(_14696_), .Y(_14697_));
AND_g _20821_ (.A(_11220_), .B(_14697_), .Y(_14698_));
NAND_g _20822_ (.A(_14693_), .B(_14698_), .Y(_14699_));
NAND_g _20823_ (.A(cpuregs_25[9]), .B(_11219_), .Y(_14700_));
NAND_g _20824_ (.A(cpuregs_29[9]), .B(_00011_[2]), .Y(_14701_));
AND_g _20825_ (.A(_00011_[0]), .B(_14701_), .Y(_14702_));
NAND_g _20826_ (.A(_14700_), .B(_14702_), .Y(_14703_));
NAND_g _20827_ (.A(cpuregs_24[9]), .B(_11219_), .Y(_14704_));
NAND_g _20828_ (.A(cpuregs_28[9]), .B(_00011_[2]), .Y(_14705_));
AND_g _20829_ (.A(_11217_), .B(_14705_), .Y(_14706_));
NAND_g _20830_ (.A(_14704_), .B(_14706_), .Y(_14707_));
AND_g _20831_ (.A(_00011_[3]), .B(_14707_), .Y(_14708_));
NAND_g _20832_ (.A(_14703_), .B(_14708_), .Y(_14709_));
NAND_g _20833_ (.A(_14699_), .B(_14709_), .Y(_14710_));
NAND_g _20834_ (.A(_11218_), .B(_14710_), .Y(_14711_));
AND_g _20835_ (.A(_14689_), .B(_14711_), .Y(_14712_));
NAND_g _20836_ (.A(cpuregs_6[9]), .B(_00011_[2]), .Y(_14713_));
NAND_g _20837_ (.A(cpuregs_2[9]), .B(_11219_), .Y(_14714_));
AND_g _20838_ (.A(_11217_), .B(_14714_), .Y(_14715_));
NAND_g _20839_ (.A(_14713_), .B(_14715_), .Y(_14716_));
NAND_g _20840_ (.A(cpuregs_3[9]), .B(_11219_), .Y(_14717_));
NAND_g _20841_ (.A(cpuregs_7[9]), .B(_00011_[2]), .Y(_14718_));
AND_g _20842_ (.A(_00011_[0]), .B(_14718_), .Y(_14719_));
NAND_g _20843_ (.A(_14717_), .B(_14719_), .Y(_14720_));
NOR_g _20844_ (.A(cpuregs_10[9]), .B(_00011_[2]), .Y(_14721_));
NOR_g _20845_ (.A(cpuregs_14[9]), .B(_11219_), .Y(_14722_));
NOR_g _20846_ (.A(_14721_), .B(_14722_), .Y(_14723_));
NOR_g _20847_ (.A(cpuregs_11[9]), .B(_00011_[2]), .Y(_14724_));
NAND_g _20848_ (.A(_11160_), .B(_00011_[2]), .Y(_14725_));
NAND_g _20849_ (.A(_14716_), .B(_14720_), .Y(_14726_));
NAND_g _20850_ (.A(_11220_), .B(_14726_), .Y(_14727_));
NAND_g _20851_ (.A(_11217_), .B(_14723_), .Y(_14728_));
NOR_g _20852_ (.A(_11217_), .B(_14724_), .Y(_14729_));
NAND_g _20853_ (.A(_14725_), .B(_14729_), .Y(_14730_));
AND_g _20854_ (.A(_00011_[3]), .B(_14730_), .Y(_14731_));
NAND_g _20855_ (.A(_14728_), .B(_14731_), .Y(_14732_));
AND_g _20856_ (.A(_14727_), .B(_14732_), .Y(_14733_));
NAND_g _20857_ (.A(_00011_[1]), .B(_14733_), .Y(_14734_));
NAND_g _20858_ (.A(cpuregs_4[9]), .B(_00011_[2]), .Y(_14735_));
NAND_g _20859_ (.A(cpuregs_0[9]), .B(_11219_), .Y(_14736_));
AND_g _20860_ (.A(_11217_), .B(_14736_), .Y(_14737_));
NAND_g _20861_ (.A(_14735_), .B(_14737_), .Y(_14738_));
NAND_g _20862_ (.A(cpuregs_1[9]), .B(_11219_), .Y(_14739_));
NAND_g _20863_ (.A(cpuregs_5[9]), .B(_00011_[2]), .Y(_14740_));
AND_g _20864_ (.A(_00011_[0]), .B(_14740_), .Y(_14741_));
NAND_g _20865_ (.A(_14739_), .B(_14741_), .Y(_14742_));
NOR_g _20866_ (.A(cpuregs_8[9]), .B(_00011_[2]), .Y(_14743_));
NOR_g _20867_ (.A(cpuregs_12[9]), .B(_11219_), .Y(_14744_));
NOR_g _20868_ (.A(_14743_), .B(_14744_), .Y(_14745_));
NOR_g _20869_ (.A(cpuregs_9[9]), .B(_00011_[2]), .Y(_14746_));
NAND_g _20870_ (.A(_11145_), .B(_00011_[2]), .Y(_14747_));
NAND_g _20871_ (.A(_14738_), .B(_14742_), .Y(_14748_));
NAND_g _20872_ (.A(_11220_), .B(_14748_), .Y(_14749_));
NAND_g _20873_ (.A(_11217_), .B(_14745_), .Y(_14750_));
NOR_g _20874_ (.A(_11217_), .B(_14746_), .Y(_14751_));
NAND_g _20875_ (.A(_14747_), .B(_14751_), .Y(_14752_));
AND_g _20876_ (.A(_00011_[3]), .B(_14752_), .Y(_14753_));
NAND_g _20877_ (.A(_14750_), .B(_14753_), .Y(_14754_));
AND_g _20878_ (.A(_14749_), .B(_14754_), .Y(_14755_));
NAND_g _20879_ (.A(_11218_), .B(_14755_), .Y(_14756_));
AND_g _20880_ (.A(_14734_), .B(_14756_), .Y(_14757_));
NAND_g _20881_ (.A(_00011_[4]), .B(_14712_), .Y(_14758_));
NAND_g _20882_ (.A(_11221_), .B(_14757_), .Y(_14759_));
AND_g _20883_ (.A(_14758_), .B(_14759_), .Y(_14760_));
AND_g _20884_ (.A(_13734_), .B(_14760_), .Y(_14761_));
NAND_g _20885_ (.A(_14358_), .B(_14761_), .Y(_14762_));
AND_g _20886_ (.A(decoded_imm[9]), .B(_13830_), .Y(_14763_));
NAND_g _20887_ (.A(_13409_), .B(_14763_), .Y(_14764_));
AND_g _20888_ (.A(_13727_), .B(_14764_), .Y(_14765_));
NAND_g _20889_ (.A(_14762_), .B(_14765_), .Y(_14766_));
AND_g _20890_ (.A(_14667_), .B(_14766_), .Y(_00512_));
NAND_g _20891_ (.A(_10990_), .B(_13728_), .Y(_14767_));
NAND_g _20892_ (.A(cpuregs_31[10]), .B(_00011_[1]), .Y(_14768_));
NAND_g _20893_ (.A(cpuregs_29[10]), .B(_11218_), .Y(_14769_));
NAND_g _20894_ (.A(_14768_), .B(_14769_), .Y(_14770_));
NAND_g _20895_ (.A(_00011_[2]), .B(_14770_), .Y(_14771_));
NAND_g _20896_ (.A(cpuregs_27[10]), .B(_00011_[1]), .Y(_14772_));
NAND_g _20897_ (.A(cpuregs_25[10]), .B(_11218_), .Y(_14773_));
NAND_g _20898_ (.A(_14772_), .B(_14773_), .Y(_14774_));
NAND_g _20899_ (.A(_11219_), .B(_14774_), .Y(_14775_));
NAND_g _20900_ (.A(_14771_), .B(_14775_), .Y(_14776_));
NAND_g _20901_ (.A(_00011_[0]), .B(_14776_), .Y(_14777_));
NAND_g _20902_ (.A(cpuregs_30[10]), .B(_00011_[1]), .Y(_14778_));
NAND_g _20903_ (.A(cpuregs_28[10]), .B(_11218_), .Y(_14779_));
NAND_g _20904_ (.A(_14778_), .B(_14779_), .Y(_14780_));
NAND_g _20905_ (.A(_00011_[2]), .B(_14780_), .Y(_14781_));
NAND_g _20906_ (.A(cpuregs_26[10]), .B(_00011_[1]), .Y(_14782_));
NAND_g _20907_ (.A(cpuregs_24[10]), .B(_11218_), .Y(_14783_));
NAND_g _20908_ (.A(_14782_), .B(_14783_), .Y(_14784_));
NAND_g _20909_ (.A(_11219_), .B(_14784_), .Y(_14785_));
NAND_g _20910_ (.A(_14781_), .B(_14785_), .Y(_14786_));
AND_g _20911_ (.A(_11217_), .B(_14786_), .Y(_14787_));
NOT_g _20912_ (.A(_14787_), .Y(_14788_));
NAND_g _20913_ (.A(_14777_), .B(_14788_), .Y(_14789_));
NAND_g _20914_ (.A(_00011_[3]), .B(_14789_), .Y(_14790_));
NOR_g _20915_ (.A(cpuregs_18[10]), .B(_00011_[2]), .Y(_14791_));
AND_g _20916_ (.A(_11015_), .B(_00011_[2]), .Y(_14792_));
NOR_g _20917_ (.A(_14791_), .B(_14792_), .Y(_14793_));
NOR_g _20918_ (.A(cpuregs_16[10]), .B(_00011_[2]), .Y(_14794_));
AND_g _20919_ (.A(_11195_), .B(_00011_[2]), .Y(_14795_));
NOR_g _20920_ (.A(_14794_), .B(_14795_), .Y(_14796_));
NAND_g _20921_ (.A(_11180_), .B(_00011_[2]), .Y(_14797_));
NOR_g _20922_ (.A(cpuregs_19[10]), .B(_00011_[2]), .Y(_14798_));
NOR_g _20923_ (.A(cpuregs_17[10]), .B(_00011_[2]), .Y(_14799_));
NAND_g _20924_ (.A(_11026_), .B(_00011_[2]), .Y(_14800_));
NOR_g _20925_ (.A(_11217_), .B(_14798_), .Y(_14801_));
NAND_g _20926_ (.A(_14797_), .B(_14801_), .Y(_14802_));
NAND_g _20927_ (.A(_11217_), .B(_14793_), .Y(_14803_));
AND_g _20928_ (.A(_14802_), .B(_14803_), .Y(_14804_));
NAND_g _20929_ (.A(_00011_[1]), .B(_14804_), .Y(_14805_));
NOR_g _20930_ (.A(_11217_), .B(_14799_), .Y(_14806_));
NAND_g _20931_ (.A(_14800_), .B(_14806_), .Y(_14807_));
NAND_g _20932_ (.A(_11217_), .B(_14796_), .Y(_14808_));
AND_g _20933_ (.A(_14807_), .B(_14808_), .Y(_14809_));
NAND_g _20934_ (.A(_11218_), .B(_14809_), .Y(_14810_));
AND_g _20935_ (.A(_14805_), .B(_14810_), .Y(_14811_));
NAND_g _20936_ (.A(_11220_), .B(_14811_), .Y(_14812_));
NAND_g _20937_ (.A(_14790_), .B(_14812_), .Y(_14813_));
NAND_g _20938_ (.A(_00011_[4]), .B(_14813_), .Y(_14814_));
NAND_g _20939_ (.A(cpuregs_13[10]), .B(_11218_), .Y(_14815_));
NAND_g _20940_ (.A(cpuregs_15[10]), .B(_00011_[1]), .Y(_14816_));
AND_g _20941_ (.A(_00011_[2]), .B(_14816_), .Y(_14817_));
NAND_g _20942_ (.A(_14815_), .B(_14817_), .Y(_14818_));
NAND_g _20943_ (.A(cpuregs_9[10]), .B(_11218_), .Y(_14819_));
NAND_g _20944_ (.A(cpuregs_11[10]), .B(_00011_[1]), .Y(_14820_));
AND_g _20945_ (.A(_11219_), .B(_14820_), .Y(_14821_));
NAND_g _20946_ (.A(_14819_), .B(_14821_), .Y(_14822_));
AND_g _20947_ (.A(_00011_[0]), .B(_14822_), .Y(_14823_));
NAND_g _20948_ (.A(_14818_), .B(_14823_), .Y(_14824_));
NAND_g _20949_ (.A(cpuregs_12[10]), .B(_11218_), .Y(_14825_));
NAND_g _20950_ (.A(cpuregs_14[10]), .B(_00011_[1]), .Y(_14826_));
AND_g _20951_ (.A(_00011_[2]), .B(_14826_), .Y(_14827_));
NAND_g _20952_ (.A(_14825_), .B(_14827_), .Y(_14828_));
NAND_g _20953_ (.A(cpuregs_8[10]), .B(_11218_), .Y(_14829_));
NAND_g _20954_ (.A(cpuregs_10[10]), .B(_00011_[1]), .Y(_14830_));
AND_g _20955_ (.A(_11219_), .B(_14830_), .Y(_14831_));
NAND_g _20956_ (.A(_14829_), .B(_14831_), .Y(_14832_));
AND_g _20957_ (.A(_11217_), .B(_14832_), .Y(_14833_));
NAND_g _20958_ (.A(_14828_), .B(_14833_), .Y(_14834_));
NAND_g _20959_ (.A(_14824_), .B(_14834_), .Y(_14835_));
NAND_g _20960_ (.A(_00011_[3]), .B(_14835_), .Y(_14836_));
NAND_g _20961_ (.A(_10941_), .B(_00011_[2]), .Y(_14837_));
NOR_g _20962_ (.A(cpuregs_2[10]), .B(_00011_[2]), .Y(_14838_));
NOR_g _20963_ (.A(_00011_[0]), .B(_14838_), .Y(_14839_));
NAND_g _20964_ (.A(_14837_), .B(_14839_), .Y(_14840_));
NAND_g _20965_ (.A(_11127_), .B(_00011_[2]), .Y(_14841_));
NOR_g _20966_ (.A(cpuregs_3[10]), .B(_00011_[2]), .Y(_14842_));
NOR_g _20967_ (.A(_11217_), .B(_14842_), .Y(_14843_));
NAND_g _20968_ (.A(_14841_), .B(_14843_), .Y(_14844_));
AND_g _20969_ (.A(_14840_), .B(_14844_), .Y(_14845_));
NAND_g _20970_ (.A(_10953_), .B(_00011_[2]), .Y(_14846_));
NOR_g _20971_ (.A(cpuregs_0[10]), .B(_00011_[2]), .Y(_14847_));
NOR_g _20972_ (.A(_00011_[0]), .B(_14847_), .Y(_14848_));
NAND_g _20973_ (.A(_14846_), .B(_14848_), .Y(_14849_));
NAND_g _20974_ (.A(_11111_), .B(_00011_[2]), .Y(_14850_));
NOR_g _20975_ (.A(cpuregs_1[10]), .B(_00011_[2]), .Y(_14851_));
NOR_g _20976_ (.A(_11217_), .B(_14851_), .Y(_14852_));
NAND_g _20977_ (.A(_14850_), .B(_14852_), .Y(_14853_));
AND_g _20978_ (.A(_14849_), .B(_14853_), .Y(_14854_));
NAND_g _20979_ (.A(_00011_[1]), .B(_14845_), .Y(_14855_));
NAND_g _20980_ (.A(_11218_), .B(_14854_), .Y(_14856_));
AND_g _20981_ (.A(_14855_), .B(_14856_), .Y(_14857_));
NAND_g _20982_ (.A(_11220_), .B(_14857_), .Y(_14858_));
NAND_g _20983_ (.A(_14836_), .B(_14858_), .Y(_14859_));
NAND_g _20984_ (.A(_11221_), .B(_14859_), .Y(_14860_));
NAND_g _20985_ (.A(_14814_), .B(_14860_), .Y(_14861_));
AND_g _20986_ (.A(_13734_), .B(_14861_), .Y(_14862_));
NAND_g _20987_ (.A(_13833_), .B(_14862_), .Y(_14863_));
NAND_g _20988_ (.A(decoded_imm[10]), .B(_13830_), .Y(_14864_));
NAND_g _20989_ (.A(_14863_), .B(_14864_), .Y(_14865_));
NAND_g _20990_ (.A(_13409_), .B(_14865_), .Y(_14866_));
NAND_g _20991_ (.A(_13724_), .B(_14862_), .Y(_14867_));
AND_g _20992_ (.A(_13727_), .B(_14867_), .Y(_14868_));
NAND_g _20993_ (.A(_14866_), .B(_14868_), .Y(_14869_));
AND_g _20994_ (.A(_14767_), .B(_14869_), .Y(_00513_));
NAND_g _20995_ (.A(_10991_), .B(_13728_), .Y(_14870_));
NAND_g _20996_ (.A(cpuregs_25[11]), .B(_11219_), .Y(_14871_));
NAND_g _20997_ (.A(cpuregs_29[11]), .B(_00011_[2]), .Y(_14872_));
AND_g _20998_ (.A(_00011_[0]), .B(_14872_), .Y(_14873_));
NAND_g _20999_ (.A(_14871_), .B(_14873_), .Y(_14874_));
NAND_g _21000_ (.A(cpuregs_24[11]), .B(_11219_), .Y(_14875_));
NAND_g _21001_ (.A(cpuregs_28[11]), .B(_00011_[2]), .Y(_14876_));
AND_g _21002_ (.A(_11217_), .B(_14876_), .Y(_14877_));
NAND_g _21003_ (.A(_14875_), .B(_14877_), .Y(_14878_));
AND_g _21004_ (.A(_11218_), .B(_14878_), .Y(_14879_));
NAND_g _21005_ (.A(_14874_), .B(_14879_), .Y(_14880_));
NAND_g _21006_ (.A(cpuregs_31[11]), .B(_00011_[2]), .Y(_14881_));
NAND_g _21007_ (.A(cpuregs_27[11]), .B(_11219_), .Y(_14882_));
AND_g _21008_ (.A(_00011_[0]), .B(_14882_), .Y(_14883_));
NAND_g _21009_ (.A(_14881_), .B(_14883_), .Y(_14884_));
NAND_g _21010_ (.A(cpuregs_26[11]), .B(_11219_), .Y(_14885_));
NAND_g _21011_ (.A(cpuregs_30[11]), .B(_00011_[2]), .Y(_14886_));
AND_g _21012_ (.A(_11217_), .B(_14886_), .Y(_14887_));
NAND_g _21013_ (.A(_14885_), .B(_14887_), .Y(_14888_));
AND_g _21014_ (.A(_00011_[1]), .B(_14888_), .Y(_14889_));
NAND_g _21015_ (.A(_14884_), .B(_14889_), .Y(_14890_));
NAND_g _21016_ (.A(_14880_), .B(_14890_), .Y(_14891_));
NAND_g _21017_ (.A(_00011_[3]), .B(_14891_), .Y(_14892_));
NAND_g _21018_ (.A(cpuregs_22[11]), .B(_00011_[2]), .Y(_14893_));
NAND_g _21019_ (.A(cpuregs_18[11]), .B(_11219_), .Y(_14894_));
AND_g _21020_ (.A(_11217_), .B(_14894_), .Y(_14895_));
NAND_g _21021_ (.A(_14893_), .B(_14895_), .Y(_14896_));
NAND_g _21022_ (.A(cpuregs_19[11]), .B(_11219_), .Y(_14897_));
NAND_g _21023_ (.A(cpuregs_23[11]), .B(_00011_[2]), .Y(_14898_));
AND_g _21024_ (.A(_00011_[0]), .B(_14898_), .Y(_14899_));
NAND_g _21025_ (.A(_14897_), .B(_14899_), .Y(_14900_));
AND_g _21026_ (.A(_00011_[1]), .B(_14900_), .Y(_14901_));
NAND_g _21027_ (.A(_14896_), .B(_14901_), .Y(_14902_));
NAND_g _21028_ (.A(cpuregs_21[11]), .B(_00011_[0]), .Y(_14903_));
NAND_g _21029_ (.A(cpuregs_20[11]), .B(_11217_), .Y(_14904_));
NAND_g _21030_ (.A(_14903_), .B(_14904_), .Y(_14905_));
NAND_g _21031_ (.A(_00011_[2]), .B(_14905_), .Y(_14906_));
NAND_g _21032_ (.A(cpuregs_17[11]), .B(_00011_[0]), .Y(_14907_));
NAND_g _21033_ (.A(cpuregs_16[11]), .B(_11217_), .Y(_14908_));
NAND_g _21034_ (.A(_14907_), .B(_14908_), .Y(_14909_));
NAND_g _21035_ (.A(_11219_), .B(_14909_), .Y(_14910_));
NAND_g _21036_ (.A(_14906_), .B(_14910_), .Y(_14911_));
NAND_g _21037_ (.A(_11218_), .B(_14911_), .Y(_14912_));
NAND_g _21038_ (.A(_14902_), .B(_14912_), .Y(_14913_));
NAND_g _21039_ (.A(_11220_), .B(_14913_), .Y(_14914_));
AND_g _21040_ (.A(_14892_), .B(_14914_), .Y(_14915_));
NAND_g _21041_ (.A(cpuregs_1[11]), .B(_11219_), .Y(_14916_));
NAND_g _21042_ (.A(cpuregs_5[11]), .B(_00011_[2]), .Y(_14917_));
AND_g _21043_ (.A(_00011_[0]), .B(_14917_), .Y(_14918_));
NAND_g _21044_ (.A(_14916_), .B(_14918_), .Y(_14919_));
NAND_g _21045_ (.A(cpuregs_0[11]), .B(_11219_), .Y(_14920_));
NAND_g _21046_ (.A(cpuregs_4[11]), .B(_00011_[2]), .Y(_14921_));
AND_g _21047_ (.A(_11217_), .B(_14921_), .Y(_14922_));
NAND_g _21048_ (.A(_14920_), .B(_14922_), .Y(_14923_));
AND_g _21049_ (.A(_11218_), .B(_14923_), .Y(_14924_));
NAND_g _21050_ (.A(_14919_), .B(_14924_), .Y(_14925_));
NAND_g _21051_ (.A(cpuregs_3[11]), .B(_11219_), .Y(_14926_));
NAND_g _21052_ (.A(cpuregs_7[11]), .B(_00011_[2]), .Y(_14927_));
AND_g _21053_ (.A(_00011_[0]), .B(_14927_), .Y(_14928_));
NAND_g _21054_ (.A(_14926_), .B(_14928_), .Y(_14929_));
NAND_g _21055_ (.A(cpuregs_2[11]), .B(_11219_), .Y(_14930_));
NAND_g _21056_ (.A(cpuregs_6[11]), .B(_00011_[2]), .Y(_14931_));
AND_g _21057_ (.A(_11217_), .B(_14931_), .Y(_14932_));
NAND_g _21058_ (.A(_14930_), .B(_14932_), .Y(_14933_));
AND_g _21059_ (.A(_00011_[1]), .B(_14933_), .Y(_14934_));
NAND_g _21060_ (.A(_14929_), .B(_14934_), .Y(_14935_));
NAND_g _21061_ (.A(_14925_), .B(_14935_), .Y(_14936_));
NAND_g _21062_ (.A(_11220_), .B(_14936_), .Y(_14937_));
NAND_g _21063_ (.A(cpuregs_14[11]), .B(_11217_), .Y(_14938_));
NAND_g _21064_ (.A(cpuregs_15[11]), .B(_00011_[0]), .Y(_14939_));
NAND_g _21065_ (.A(_14938_), .B(_14939_), .Y(_14940_));
NAND_g _21066_ (.A(_00011_[2]), .B(_14940_), .Y(_14941_));
NAND_g _21067_ (.A(cpuregs_10[11]), .B(_11217_), .Y(_14942_));
NAND_g _21068_ (.A(cpuregs_11[11]), .B(_00011_[0]), .Y(_14943_));
NAND_g _21069_ (.A(_14942_), .B(_14943_), .Y(_14944_));
NAND_g _21070_ (.A(_11219_), .B(_14944_), .Y(_14945_));
AND_g _21071_ (.A(_14941_), .B(_14945_), .Y(_14946_));
NAND_g _21072_ (.A(cpuregs_12[11]), .B(_11217_), .Y(_14947_));
NAND_g _21073_ (.A(cpuregs_13[11]), .B(_00011_[0]), .Y(_14948_));
NAND_g _21074_ (.A(_14947_), .B(_14948_), .Y(_14949_));
NAND_g _21075_ (.A(_00011_[2]), .B(_14949_), .Y(_14950_));
NAND_g _21076_ (.A(cpuregs_8[11]), .B(_11217_), .Y(_14951_));
NAND_g _21077_ (.A(cpuregs_9[11]), .B(_00011_[0]), .Y(_14952_));
NAND_g _21078_ (.A(_14951_), .B(_14952_), .Y(_14953_));
NAND_g _21079_ (.A(_11219_), .B(_14953_), .Y(_14954_));
AND_g _21080_ (.A(_14950_), .B(_14954_), .Y(_14955_));
NAND_g _21081_ (.A(_11218_), .B(_14955_), .Y(_14956_));
NAND_g _21082_ (.A(_00011_[1]), .B(_14946_), .Y(_14957_));
AND_g _21083_ (.A(_00011_[3]), .B(_14956_), .Y(_14958_));
NAND_g _21084_ (.A(_14957_), .B(_14958_), .Y(_14959_));
NAND_g _21085_ (.A(_00011_[4]), .B(_14915_), .Y(_14960_));
AND_g _21086_ (.A(_11221_), .B(_14937_), .Y(_14961_));
NAND_g _21087_ (.A(_14959_), .B(_14961_), .Y(_14962_));
AND_g _21088_ (.A(_13734_), .B(_14962_), .Y(_14963_));
AND_g _21089_ (.A(_14960_), .B(_14963_), .Y(_14964_));
NAND_g _21090_ (.A(_14358_), .B(_14964_), .Y(_14965_));
AND_g _21091_ (.A(decoded_imm[11]), .B(_13830_), .Y(_14966_));
NAND_g _21092_ (.A(_13409_), .B(_14966_), .Y(_14967_));
AND_g _21093_ (.A(_13727_), .B(_14967_), .Y(_14968_));
NAND_g _21094_ (.A(_14965_), .B(_14968_), .Y(_14969_));
AND_g _21095_ (.A(_14870_), .B(_14969_), .Y(_00514_));
NAND_g _21096_ (.A(_10992_), .B(_13728_), .Y(_14970_));
NOR_g _21097_ (.A(cpuregs_16[12]), .B(_00011_[2]), .Y(_14971_));
AND_g _21098_ (.A(_11197_), .B(_00011_[2]), .Y(_14972_));
NOR_g _21099_ (.A(_14971_), .B(_14972_), .Y(_14973_));
NOR_g _21100_ (.A(cpuregs_18[12]), .B(_00011_[2]), .Y(_14974_));
NOR_g _21101_ (.A(cpuregs_22[12]), .B(_11219_), .Y(_14975_));
NOR_g _21102_ (.A(_14974_), .B(_14975_), .Y(_14976_));
NOR_g _21103_ (.A(cpuregs_17[12]), .B(_00011_[2]), .Y(_14977_));
NAND_g _21104_ (.A(_11028_), .B(_00011_[2]), .Y(_14978_));
NAND_g _21105_ (.A(_11182_), .B(_00011_[2]), .Y(_14979_));
NOR_g _21106_ (.A(cpuregs_19[12]), .B(_00011_[2]), .Y(_14980_));
NOR_g _21107_ (.A(_11217_), .B(_14980_), .Y(_14981_));
NAND_g _21108_ (.A(_14979_), .B(_14981_), .Y(_14982_));
NAND_g _21109_ (.A(_11217_), .B(_14976_), .Y(_14983_));
AND_g _21110_ (.A(_14982_), .B(_14983_), .Y(_14984_));
NAND_g _21111_ (.A(_00011_[1]), .B(_14984_), .Y(_14985_));
NOR_g _21112_ (.A(_11217_), .B(_14977_), .Y(_14986_));
NAND_g _21113_ (.A(_14978_), .B(_14986_), .Y(_14987_));
NAND_g _21114_ (.A(_11217_), .B(_14973_), .Y(_14988_));
AND_g _21115_ (.A(_14987_), .B(_14988_), .Y(_14989_));
NAND_g _21116_ (.A(_11218_), .B(_14989_), .Y(_14990_));
AND_g _21117_ (.A(_11220_), .B(_14990_), .Y(_14991_));
NAND_g _21118_ (.A(_14985_), .B(_14991_), .Y(_14992_));
NAND_g _21119_ (.A(cpuregs_27[12]), .B(_00011_[1]), .Y(_14993_));
NAND_g _21120_ (.A(cpuregs_25[12]), .B(_11218_), .Y(_14994_));
NAND_g _21121_ (.A(_14993_), .B(_14994_), .Y(_14995_));
NAND_g _21122_ (.A(_11219_), .B(_14995_), .Y(_14996_));
NAND_g _21123_ (.A(cpuregs_31[12]), .B(_00011_[1]), .Y(_14997_));
NAND_g _21124_ (.A(cpuregs_29[12]), .B(_11218_), .Y(_14998_));
NAND_g _21125_ (.A(_14997_), .B(_14998_), .Y(_14999_));
NAND_g _21126_ (.A(_00011_[2]), .B(_14999_), .Y(_15000_));
AND_g _21127_ (.A(_00011_[0]), .B(_15000_), .Y(_15001_));
NAND_g _21128_ (.A(_14996_), .B(_15001_), .Y(_15002_));
NAND_g _21129_ (.A(cpuregs_26[12]), .B(_00011_[1]), .Y(_15003_));
NAND_g _21130_ (.A(cpuregs_24[12]), .B(_11218_), .Y(_15004_));
NAND_g _21131_ (.A(_15003_), .B(_15004_), .Y(_15005_));
NAND_g _21132_ (.A(_11219_), .B(_15005_), .Y(_15006_));
NAND_g _21133_ (.A(cpuregs_30[12]), .B(_00011_[1]), .Y(_15007_));
NAND_g _21134_ (.A(cpuregs_28[12]), .B(_11218_), .Y(_15008_));
NAND_g _21135_ (.A(_15007_), .B(_15008_), .Y(_15009_));
NAND_g _21136_ (.A(_00011_[2]), .B(_15009_), .Y(_15010_));
AND_g _21137_ (.A(_11217_), .B(_15010_), .Y(_15011_));
NAND_g _21138_ (.A(_15006_), .B(_15011_), .Y(_15012_));
AND_g _21139_ (.A(_00011_[3]), .B(_15012_), .Y(_15013_));
NAND_g _21140_ (.A(_15002_), .B(_15013_), .Y(_15014_));
AND_g _21141_ (.A(_14992_), .B(_15014_), .Y(_15015_));
NAND_g _21142_ (.A(cpuregs_1[12]), .B(_11219_), .Y(_15016_));
NAND_g _21143_ (.A(cpuregs_5[12]), .B(_00011_[2]), .Y(_15017_));
AND_g _21144_ (.A(_00011_[0]), .B(_15017_), .Y(_15018_));
NAND_g _21145_ (.A(_15016_), .B(_15018_), .Y(_15019_));
NAND_g _21146_ (.A(cpuregs_0[12]), .B(_11219_), .Y(_15020_));
NAND_g _21147_ (.A(cpuregs_4[12]), .B(_00011_[2]), .Y(_15021_));
AND_g _21148_ (.A(_11217_), .B(_15021_), .Y(_15022_));
NAND_g _21149_ (.A(_15020_), .B(_15022_), .Y(_15023_));
AND_g _21150_ (.A(_11218_), .B(_15023_), .Y(_15024_));
NAND_g _21151_ (.A(_15019_), .B(_15024_), .Y(_15025_));
NAND_g _21152_ (.A(cpuregs_3[12]), .B(_11219_), .Y(_15026_));
NAND_g _21153_ (.A(cpuregs_7[12]), .B(_00011_[2]), .Y(_15027_));
AND_g _21154_ (.A(_00011_[0]), .B(_15027_), .Y(_15028_));
NAND_g _21155_ (.A(_15026_), .B(_15028_), .Y(_15029_));
NAND_g _21156_ (.A(cpuregs_2[12]), .B(_11219_), .Y(_15030_));
NAND_g _21157_ (.A(cpuregs_6[12]), .B(_00011_[2]), .Y(_15031_));
AND_g _21158_ (.A(_11217_), .B(_15031_), .Y(_15032_));
NAND_g _21159_ (.A(_15030_), .B(_15032_), .Y(_15033_));
AND_g _21160_ (.A(_00011_[1]), .B(_15033_), .Y(_15034_));
NAND_g _21161_ (.A(_15029_), .B(_15034_), .Y(_15035_));
NAND_g _21162_ (.A(_15025_), .B(_15035_), .Y(_15036_));
NAND_g _21163_ (.A(_11220_), .B(_15036_), .Y(_15037_));
NAND_g _21164_ (.A(cpuregs_14[12]), .B(_11217_), .Y(_15038_));
NAND_g _21165_ (.A(cpuregs_15[12]), .B(_00011_[0]), .Y(_15039_));
NAND_g _21166_ (.A(_15038_), .B(_15039_), .Y(_15040_));
NAND_g _21167_ (.A(_00011_[2]), .B(_15040_), .Y(_15041_));
NAND_g _21168_ (.A(cpuregs_10[12]), .B(_11217_), .Y(_15042_));
NAND_g _21169_ (.A(cpuregs_11[12]), .B(_00011_[0]), .Y(_15043_));
NAND_g _21170_ (.A(_15042_), .B(_15043_), .Y(_15044_));
NAND_g _21171_ (.A(_11219_), .B(_15044_), .Y(_15045_));
AND_g _21172_ (.A(_15041_), .B(_15045_), .Y(_15046_));
NAND_g _21173_ (.A(cpuregs_12[12]), .B(_11217_), .Y(_15047_));
NAND_g _21174_ (.A(cpuregs_13[12]), .B(_00011_[0]), .Y(_15048_));
NAND_g _21175_ (.A(_15047_), .B(_15048_), .Y(_15049_));
NAND_g _21176_ (.A(_00011_[2]), .B(_15049_), .Y(_15050_));
NAND_g _21177_ (.A(cpuregs_8[12]), .B(_11217_), .Y(_15051_));
NAND_g _21178_ (.A(cpuregs_9[12]), .B(_00011_[0]), .Y(_15052_));
NAND_g _21179_ (.A(_15051_), .B(_15052_), .Y(_15053_));
NAND_g _21180_ (.A(_11219_), .B(_15053_), .Y(_15054_));
AND_g _21181_ (.A(_15050_), .B(_15054_), .Y(_15055_));
NAND_g _21182_ (.A(_11218_), .B(_15055_), .Y(_15056_));
NAND_g _21183_ (.A(_00011_[1]), .B(_15046_), .Y(_15057_));
AND_g _21184_ (.A(_00011_[3]), .B(_15056_), .Y(_15058_));
NAND_g _21185_ (.A(_15057_), .B(_15058_), .Y(_15059_));
NAND_g _21186_ (.A(_00011_[4]), .B(_15015_), .Y(_15060_));
AND_g _21187_ (.A(_11221_), .B(_15037_), .Y(_15061_));
NAND_g _21188_ (.A(_15059_), .B(_15061_), .Y(_15062_));
AND_g _21189_ (.A(_13734_), .B(_15062_), .Y(_15063_));
AND_g _21190_ (.A(_15060_), .B(_15063_), .Y(_15064_));
NAND_g _21191_ (.A(_14358_), .B(_15064_), .Y(_15065_));
AND_g _21192_ (.A(decoded_imm[12]), .B(_13830_), .Y(_15066_));
NAND_g _21193_ (.A(_13409_), .B(_15066_), .Y(_15067_));
AND_g _21194_ (.A(_13727_), .B(_15067_), .Y(_15068_));
NAND_g _21195_ (.A(_15065_), .B(_15068_), .Y(_15069_));
AND_g _21196_ (.A(_14970_), .B(_15069_), .Y(_00515_));
NAND_g _21197_ (.A(_10993_), .B(_13728_), .Y(_15070_));
NAND_g _21198_ (.A(cpuregs_29[13]), .B(_00011_[2]), .Y(_15071_));
NAND_g _21199_ (.A(cpuregs_25[13]), .B(_11219_), .Y(_15072_));
AND_g _21200_ (.A(_00011_[0]), .B(_15072_), .Y(_15073_));
NAND_g _21201_ (.A(_15071_), .B(_15073_), .Y(_15074_));
NAND_g _21202_ (.A(cpuregs_24[13]), .B(_11219_), .Y(_15075_));
NAND_g _21203_ (.A(cpuregs_28[13]), .B(_00011_[2]), .Y(_15076_));
AND_g _21204_ (.A(_11217_), .B(_15076_), .Y(_15077_));
NAND_g _21205_ (.A(_15075_), .B(_15077_), .Y(_15078_));
AND_g _21206_ (.A(_11218_), .B(_15078_), .Y(_15079_));
NAND_g _21207_ (.A(_15074_), .B(_15079_), .Y(_15080_));
NAND_g _21208_ (.A(cpuregs_27[13]), .B(_11219_), .Y(_15081_));
NAND_g _21209_ (.A(cpuregs_31[13]), .B(_00011_[2]), .Y(_15082_));
AND_g _21210_ (.A(_00011_[0]), .B(_15082_), .Y(_15083_));
NAND_g _21211_ (.A(_15081_), .B(_15083_), .Y(_15084_));
NAND_g _21212_ (.A(cpuregs_26[13]), .B(_11219_), .Y(_15085_));
NAND_g _21213_ (.A(cpuregs_30[13]), .B(_00011_[2]), .Y(_15086_));
AND_g _21214_ (.A(_11217_), .B(_15086_), .Y(_15087_));
NAND_g _21215_ (.A(_15085_), .B(_15087_), .Y(_15088_));
AND_g _21216_ (.A(_00011_[1]), .B(_15088_), .Y(_15089_));
NAND_g _21217_ (.A(_15084_), .B(_15089_), .Y(_15090_));
NAND_g _21218_ (.A(_15080_), .B(_15090_), .Y(_15091_));
NAND_g _21219_ (.A(_00011_[4]), .B(_15091_), .Y(_15092_));
NAND_g _21220_ (.A(cpuregs_14[13]), .B(_11217_), .Y(_15093_));
NAND_g _21221_ (.A(cpuregs_15[13]), .B(_00011_[0]), .Y(_15094_));
NAND_g _21222_ (.A(_15093_), .B(_15094_), .Y(_15095_));
NAND_g _21223_ (.A(_00011_[2]), .B(_15095_), .Y(_15096_));
NAND_g _21224_ (.A(cpuregs_10[13]), .B(_11217_), .Y(_15097_));
NAND_g _21225_ (.A(cpuregs_11[13]), .B(_00011_[0]), .Y(_15098_));
NAND_g _21226_ (.A(_15097_), .B(_15098_), .Y(_15099_));
NAND_g _21227_ (.A(_11219_), .B(_15099_), .Y(_15100_));
NAND_g _21228_ (.A(_15096_), .B(_15100_), .Y(_15101_));
NAND_g _21229_ (.A(_00011_[1]), .B(_15101_), .Y(_15102_));
NAND_g _21230_ (.A(cpuregs_12[13]), .B(_11217_), .Y(_15103_));
NAND_g _21231_ (.A(cpuregs_13[13]), .B(_00011_[0]), .Y(_15104_));
NAND_g _21232_ (.A(_15103_), .B(_15104_), .Y(_15105_));
NAND_g _21233_ (.A(_00011_[2]), .B(_15105_), .Y(_15106_));
NAND_g _21234_ (.A(cpuregs_8[13]), .B(_11217_), .Y(_15107_));
NAND_g _21235_ (.A(cpuregs_9[13]), .B(_00011_[0]), .Y(_15108_));
NAND_g _21236_ (.A(_15107_), .B(_15108_), .Y(_15109_));
NAND_g _21237_ (.A(_11219_), .B(_15109_), .Y(_15110_));
NAND_g _21238_ (.A(_15106_), .B(_15110_), .Y(_15111_));
NAND_g _21239_ (.A(_11218_), .B(_15111_), .Y(_15112_));
NAND_g _21240_ (.A(_15102_), .B(_15112_), .Y(_15113_));
NAND_g _21241_ (.A(_11221_), .B(_15113_), .Y(_15114_));
NAND_g _21242_ (.A(_15092_), .B(_15114_), .Y(_15115_));
NAND_g _21243_ (.A(_00011_[3]), .B(_15115_), .Y(_15116_));
NAND_g _21244_ (.A(cpuregs_1[13]), .B(_11219_), .Y(_15117_));
NAND_g _21245_ (.A(cpuregs_5[13]), .B(_00011_[2]), .Y(_15118_));
AND_g _21246_ (.A(_00011_[0]), .B(_15118_), .Y(_15119_));
NAND_g _21247_ (.A(_15117_), .B(_15119_), .Y(_15120_));
NAND_g _21248_ (.A(cpuregs_0[13]), .B(_11219_), .Y(_15121_));
NAND_g _21249_ (.A(cpuregs_4[13]), .B(_00011_[2]), .Y(_15122_));
AND_g _21250_ (.A(_11217_), .B(_15122_), .Y(_15123_));
NAND_g _21251_ (.A(_15121_), .B(_15123_), .Y(_15124_));
AND_g _21252_ (.A(_11218_), .B(_15124_), .Y(_15125_));
NAND_g _21253_ (.A(_15120_), .B(_15125_), .Y(_15126_));
NAND_g _21254_ (.A(cpuregs_3[13]), .B(_11219_), .Y(_15127_));
NAND_g _21255_ (.A(cpuregs_7[13]), .B(_00011_[2]), .Y(_15128_));
AND_g _21256_ (.A(_00011_[0]), .B(_15128_), .Y(_15129_));
NAND_g _21257_ (.A(_15127_), .B(_15129_), .Y(_15130_));
NAND_g _21258_ (.A(cpuregs_2[13]), .B(_11219_), .Y(_15131_));
NAND_g _21259_ (.A(cpuregs_6[13]), .B(_00011_[2]), .Y(_15132_));
AND_g _21260_ (.A(_11217_), .B(_15132_), .Y(_15133_));
NAND_g _21261_ (.A(_15131_), .B(_15133_), .Y(_15134_));
AND_g _21262_ (.A(_00011_[1]), .B(_15134_), .Y(_15135_));
NAND_g _21263_ (.A(_15130_), .B(_15135_), .Y(_15136_));
NAND_g _21264_ (.A(_15126_), .B(_15136_), .Y(_15137_));
NAND_g _21265_ (.A(_11221_), .B(_15137_), .Y(_15138_));
NAND_g _21266_ (.A(cpuregs_19[13]), .B(_00011_[1]), .Y(_15139_));
NAND_g _21267_ (.A(cpuregs_17[13]), .B(_11218_), .Y(_15140_));
NAND_g _21268_ (.A(_15139_), .B(_15140_), .Y(_15141_));
NAND_g _21269_ (.A(_11219_), .B(_15141_), .Y(_15142_));
NAND_g _21270_ (.A(cpuregs_23[13]), .B(_00011_[1]), .Y(_15143_));
NAND_g _21271_ (.A(cpuregs_21[13]), .B(_11218_), .Y(_15144_));
NAND_g _21272_ (.A(_15143_), .B(_15144_), .Y(_15145_));
NAND_g _21273_ (.A(_00011_[2]), .B(_15145_), .Y(_15146_));
AND_g _21274_ (.A(_00011_[0]), .B(_15146_), .Y(_15147_));
NAND_g _21275_ (.A(_15142_), .B(_15147_), .Y(_15148_));
NAND_g _21276_ (.A(cpuregs_18[13]), .B(_00011_[1]), .Y(_15149_));
NAND_g _21277_ (.A(cpuregs_16[13]), .B(_11218_), .Y(_15150_));
NAND_g _21278_ (.A(_15149_), .B(_15150_), .Y(_15151_));
NAND_g _21279_ (.A(_11219_), .B(_15151_), .Y(_15152_));
NAND_g _21280_ (.A(cpuregs_22[13]), .B(_00011_[1]), .Y(_15153_));
NAND_g _21281_ (.A(cpuregs_20[13]), .B(_11218_), .Y(_15154_));
NAND_g _21282_ (.A(_15153_), .B(_15154_), .Y(_15155_));
NAND_g _21283_ (.A(_00011_[2]), .B(_15155_), .Y(_15156_));
AND_g _21284_ (.A(_11217_), .B(_15156_), .Y(_15157_));
NAND_g _21285_ (.A(_15152_), .B(_15157_), .Y(_15158_));
AND_g _21286_ (.A(_00011_[4]), .B(_15158_), .Y(_15159_));
NAND_g _21287_ (.A(_15148_), .B(_15159_), .Y(_15160_));
NAND_g _21288_ (.A(_15138_), .B(_15160_), .Y(_15161_));
NAND_g _21289_ (.A(_11220_), .B(_15161_), .Y(_15162_));
NAND_g _21290_ (.A(_15116_), .B(_15162_), .Y(_15163_));
AND_g _21291_ (.A(_13734_), .B(_15163_), .Y(_15164_));
NAND_g _21292_ (.A(_13833_), .B(_15164_), .Y(_15165_));
NAND_g _21293_ (.A(decoded_imm[13]), .B(_13830_), .Y(_15166_));
NAND_g _21294_ (.A(_15165_), .B(_15166_), .Y(_15167_));
NAND_g _21295_ (.A(_13409_), .B(_15167_), .Y(_15168_));
AND_g _21296_ (.A(_13724_), .B(_15164_), .Y(_15169_));
NOR_g _21297_ (.A(_13728_), .B(_15169_), .Y(_15170_));
NAND_g _21298_ (.A(_15168_), .B(_15170_), .Y(_15171_));
AND_g _21299_ (.A(_15070_), .B(_15171_), .Y(_00516_));
NAND_g _21300_ (.A(_10994_), .B(_13728_), .Y(_15172_));
NAND_g _21301_ (.A(cpuregs_31[14]), .B(_00011_[1]), .Y(_15173_));
NAND_g _21302_ (.A(cpuregs_29[14]), .B(_11218_), .Y(_15174_));
NAND_g _21303_ (.A(_15173_), .B(_15174_), .Y(_15175_));
NAND_g _21304_ (.A(_00011_[2]), .B(_15175_), .Y(_15176_));
NAND_g _21305_ (.A(cpuregs_27[14]), .B(_00011_[1]), .Y(_15177_));
NAND_g _21306_ (.A(cpuregs_25[14]), .B(_11218_), .Y(_15178_));
NAND_g _21307_ (.A(_15177_), .B(_15178_), .Y(_15179_));
NAND_g _21308_ (.A(_11219_), .B(_15179_), .Y(_15180_));
NAND_g _21309_ (.A(_15176_), .B(_15180_), .Y(_15181_));
NAND_g _21310_ (.A(_00011_[0]), .B(_15181_), .Y(_15182_));
NAND_g _21311_ (.A(cpuregs_30[14]), .B(_00011_[1]), .Y(_15183_));
NAND_g _21312_ (.A(cpuregs_28[14]), .B(_11218_), .Y(_15184_));
NAND_g _21313_ (.A(_15183_), .B(_15184_), .Y(_15185_));
NAND_g _21314_ (.A(_00011_[2]), .B(_15185_), .Y(_15186_));
NAND_g _21315_ (.A(cpuregs_26[14]), .B(_00011_[1]), .Y(_15187_));
NAND_g _21316_ (.A(cpuregs_24[14]), .B(_11218_), .Y(_15188_));
NAND_g _21317_ (.A(_15187_), .B(_15188_), .Y(_15189_));
NAND_g _21318_ (.A(_11219_), .B(_15189_), .Y(_15190_));
NAND_g _21319_ (.A(_15186_), .B(_15190_), .Y(_15191_));
AND_g _21320_ (.A(_11217_), .B(_15191_), .Y(_15192_));
NOT_g _21321_ (.A(_15192_), .Y(_15193_));
NAND_g _21322_ (.A(_15182_), .B(_15193_), .Y(_15194_));
NAND_g _21323_ (.A(_00011_[3]), .B(_15194_), .Y(_15195_));
NOR_g _21324_ (.A(cpuregs_18[14]), .B(_00011_[2]), .Y(_15196_));
NOR_g _21325_ (.A(cpuregs_22[14]), .B(_11219_), .Y(_15197_));
NOR_g _21326_ (.A(_15196_), .B(_15197_), .Y(_15198_));
NOR_g _21327_ (.A(cpuregs_16[14]), .B(_00011_[2]), .Y(_15199_));
NOR_g _21328_ (.A(cpuregs_20[14]), .B(_11219_), .Y(_15200_));
NOR_g _21329_ (.A(_15199_), .B(_15200_), .Y(_15201_));
NAND_g _21330_ (.A(_11183_), .B(_00011_[2]), .Y(_15202_));
NOR_g _21331_ (.A(cpuregs_19[14]), .B(_00011_[2]), .Y(_15203_));
NOR_g _21332_ (.A(cpuregs_17[14]), .B(_00011_[2]), .Y(_15204_));
NAND_g _21333_ (.A(_11029_), .B(_00011_[2]), .Y(_15205_));
NOR_g _21334_ (.A(_11217_), .B(_15203_), .Y(_15206_));
NAND_g _21335_ (.A(_15202_), .B(_15206_), .Y(_15207_));
NAND_g _21336_ (.A(_11217_), .B(_15198_), .Y(_15208_));
AND_g _21337_ (.A(_15207_), .B(_15208_), .Y(_15209_));
NAND_g _21338_ (.A(_00011_[1]), .B(_15209_), .Y(_15210_));
NOR_g _21339_ (.A(_11217_), .B(_15204_), .Y(_15211_));
NAND_g _21340_ (.A(_15205_), .B(_15211_), .Y(_15212_));
NAND_g _21341_ (.A(_11217_), .B(_15201_), .Y(_15213_));
AND_g _21342_ (.A(_15212_), .B(_15213_), .Y(_15214_));
NAND_g _21343_ (.A(_11218_), .B(_15214_), .Y(_15215_));
AND_g _21344_ (.A(_15210_), .B(_15215_), .Y(_15216_));
NAND_g _21345_ (.A(_11220_), .B(_15216_), .Y(_15217_));
NAND_g _21346_ (.A(_15195_), .B(_15217_), .Y(_15218_));
NAND_g _21347_ (.A(_00011_[4]), .B(_15218_), .Y(_15219_));
NAND_g _21348_ (.A(cpuregs_13[14]), .B(_11218_), .Y(_15220_));
NAND_g _21349_ (.A(cpuregs_15[14]), .B(_00011_[1]), .Y(_15221_));
AND_g _21350_ (.A(_00011_[2]), .B(_15221_), .Y(_15222_));
NAND_g _21351_ (.A(_15220_), .B(_15222_), .Y(_15223_));
NAND_g _21352_ (.A(cpuregs_9[14]), .B(_11218_), .Y(_15224_));
NAND_g _21353_ (.A(cpuregs_11[14]), .B(_00011_[1]), .Y(_15225_));
AND_g _21354_ (.A(_11219_), .B(_15225_), .Y(_15226_));
NAND_g _21355_ (.A(_15224_), .B(_15226_), .Y(_15227_));
AND_g _21356_ (.A(_00011_[0]), .B(_15227_), .Y(_15228_));
NAND_g _21357_ (.A(_15223_), .B(_15228_), .Y(_15229_));
NAND_g _21358_ (.A(cpuregs_12[14]), .B(_11218_), .Y(_15230_));
NAND_g _21359_ (.A(cpuregs_14[14]), .B(_00011_[1]), .Y(_15231_));
AND_g _21360_ (.A(_00011_[2]), .B(_15231_), .Y(_15232_));
NAND_g _21361_ (.A(_15230_), .B(_15232_), .Y(_15233_));
NAND_g _21362_ (.A(cpuregs_8[14]), .B(_11218_), .Y(_15234_));
NAND_g _21363_ (.A(cpuregs_10[14]), .B(_00011_[1]), .Y(_15235_));
AND_g _21364_ (.A(_11219_), .B(_15235_), .Y(_15236_));
NAND_g _21365_ (.A(_15234_), .B(_15236_), .Y(_15237_));
AND_g _21366_ (.A(_11217_), .B(_15237_), .Y(_15238_));
NAND_g _21367_ (.A(_15233_), .B(_15238_), .Y(_15239_));
NAND_g _21368_ (.A(_15229_), .B(_15239_), .Y(_15240_));
NAND_g _21369_ (.A(_00011_[3]), .B(_15240_), .Y(_15241_));
NAND_g _21370_ (.A(_10943_), .B(_00011_[2]), .Y(_15242_));
NOR_g _21371_ (.A(cpuregs_2[14]), .B(_00011_[2]), .Y(_15243_));
NOR_g _21372_ (.A(_00011_[0]), .B(_15243_), .Y(_15244_));
NAND_g _21373_ (.A(_15242_), .B(_15244_), .Y(_15245_));
NAND_g _21374_ (.A(_11129_), .B(_00011_[2]), .Y(_15246_));
NOR_g _21375_ (.A(cpuregs_3[14]), .B(_00011_[2]), .Y(_15247_));
NOR_g _21376_ (.A(_11217_), .B(_15247_), .Y(_15248_));
NAND_g _21377_ (.A(_15246_), .B(_15248_), .Y(_15249_));
AND_g _21378_ (.A(_15245_), .B(_15249_), .Y(_15250_));
NAND_g _21379_ (.A(_10955_), .B(_00011_[2]), .Y(_15251_));
NOR_g _21380_ (.A(cpuregs_0[14]), .B(_00011_[2]), .Y(_15252_));
NOR_g _21381_ (.A(_00011_[0]), .B(_15252_), .Y(_15253_));
NAND_g _21382_ (.A(_15251_), .B(_15253_), .Y(_15254_));
NAND_g _21383_ (.A(_11113_), .B(_00011_[2]), .Y(_15255_));
NOR_g _21384_ (.A(cpuregs_1[14]), .B(_00011_[2]), .Y(_15256_));
NOR_g _21385_ (.A(_11217_), .B(_15256_), .Y(_15257_));
NAND_g _21386_ (.A(_15255_), .B(_15257_), .Y(_15258_));
AND_g _21387_ (.A(_15254_), .B(_15258_), .Y(_15259_));
NAND_g _21388_ (.A(_00011_[1]), .B(_15250_), .Y(_15260_));
NAND_g _21389_ (.A(_11218_), .B(_15259_), .Y(_15261_));
AND_g _21390_ (.A(_15260_), .B(_15261_), .Y(_15262_));
NAND_g _21391_ (.A(_11220_), .B(_15262_), .Y(_15263_));
NAND_g _21392_ (.A(_15241_), .B(_15263_), .Y(_15264_));
NAND_g _21393_ (.A(_11221_), .B(_15264_), .Y(_15265_));
NAND_g _21394_ (.A(_15219_), .B(_15265_), .Y(_15266_));
AND_g _21395_ (.A(_13734_), .B(_15266_), .Y(_15267_));
NAND_g _21396_ (.A(_14358_), .B(_15267_), .Y(_15268_));
AND_g _21397_ (.A(decoded_imm[14]), .B(_13830_), .Y(_15269_));
NAND_g _21398_ (.A(_13409_), .B(_15269_), .Y(_15270_));
AND_g _21399_ (.A(_13727_), .B(_15270_), .Y(_15271_));
NAND_g _21400_ (.A(_15268_), .B(_15271_), .Y(_15272_));
AND_g _21401_ (.A(_15172_), .B(_15272_), .Y(_00517_));
NAND_g _21402_ (.A(_10995_), .B(_13728_), .Y(_15273_));
NAND_g _21403_ (.A(cpuregs_19[15]), .B(_11219_), .Y(_15274_));
NAND_g _21404_ (.A(cpuregs_23[15]), .B(_00011_[2]), .Y(_15275_));
AND_g _21405_ (.A(_00011_[0]), .B(_15275_), .Y(_15276_));
NAND_g _21406_ (.A(_15274_), .B(_15276_), .Y(_15277_));
NAND_g _21407_ (.A(cpuregs_18[15]), .B(_11219_), .Y(_15278_));
NAND_g _21408_ (.A(cpuregs_22[15]), .B(_00011_[2]), .Y(_15279_));
AND_g _21409_ (.A(_11217_), .B(_15279_), .Y(_15280_));
NAND_g _21410_ (.A(_15278_), .B(_15280_), .Y(_15281_));
AND_g _21411_ (.A(_11220_), .B(_15281_), .Y(_15282_));
NAND_g _21412_ (.A(_15277_), .B(_15282_), .Y(_15283_));
NAND_g _21413_ (.A(cpuregs_27[15]), .B(_11219_), .Y(_15284_));
NAND_g _21414_ (.A(cpuregs_31[15]), .B(_00011_[2]), .Y(_15285_));
AND_g _21415_ (.A(_00011_[0]), .B(_15285_), .Y(_15286_));
NAND_g _21416_ (.A(_15284_), .B(_15286_), .Y(_15287_));
NAND_g _21417_ (.A(cpuregs_26[15]), .B(_11219_), .Y(_15288_));
NAND_g _21418_ (.A(cpuregs_30[15]), .B(_00011_[2]), .Y(_15289_));
AND_g _21419_ (.A(_11217_), .B(_15289_), .Y(_15290_));
NAND_g _21420_ (.A(_15288_), .B(_15290_), .Y(_15291_));
AND_g _21421_ (.A(_00011_[3]), .B(_15291_), .Y(_15292_));
NAND_g _21422_ (.A(_15287_), .B(_15292_), .Y(_15293_));
NAND_g _21423_ (.A(_15283_), .B(_15293_), .Y(_15294_));
NAND_g _21424_ (.A(_00011_[1]), .B(_15294_), .Y(_15295_));
NOR_g _21425_ (.A(cpuregs_16[15]), .B(_00011_[2]), .Y(_15296_));
NOR_g _21426_ (.A(cpuregs_20[15]), .B(_11219_), .Y(_15297_));
NOR_g _21427_ (.A(_15296_), .B(_15297_), .Y(_15298_));
NOR_g _21428_ (.A(cpuregs_17[15]), .B(_00011_[2]), .Y(_15299_));
NAND_g _21429_ (.A(_11030_), .B(_00011_[2]), .Y(_15300_));
NOR_g _21430_ (.A(cpuregs_24[15]), .B(_00011_[2]), .Y(_15301_));
NOR_g _21431_ (.A(cpuregs_28[15]), .B(_11219_), .Y(_15302_));
NOR_g _21432_ (.A(_15301_), .B(_15302_), .Y(_15303_));
NOR_g _21433_ (.A(cpuregs_25[15]), .B(_00011_[2]), .Y(_15304_));
NAND_g _21434_ (.A(_10929_), .B(_00011_[2]), .Y(_15305_));
NAND_g _21435_ (.A(_11217_), .B(_15298_), .Y(_15306_));
NOR_g _21436_ (.A(_11217_), .B(_15299_), .Y(_15307_));
NAND_g _21437_ (.A(_15300_), .B(_15307_), .Y(_15308_));
AND_g _21438_ (.A(_15306_), .B(_15308_), .Y(_15309_));
NAND_g _21439_ (.A(_11220_), .B(_15309_), .Y(_15310_));
NOR_g _21440_ (.A(_11217_), .B(_15304_), .Y(_15311_));
NAND_g _21441_ (.A(_15305_), .B(_15311_), .Y(_15312_));
NAND_g _21442_ (.A(_11217_), .B(_15303_), .Y(_15313_));
AND_g _21443_ (.A(_15312_), .B(_15313_), .Y(_15314_));
NAND_g _21444_ (.A(_00011_[3]), .B(_15314_), .Y(_15315_));
AND_g _21445_ (.A(_15310_), .B(_15315_), .Y(_15316_));
NAND_g _21446_ (.A(_11218_), .B(_15316_), .Y(_15317_));
NAND_g _21447_ (.A(cpuregs_14[15]), .B(_11217_), .Y(_15318_));
NAND_g _21448_ (.A(cpuregs_15[15]), .B(_00011_[0]), .Y(_15319_));
NAND_g _21449_ (.A(_15318_), .B(_15319_), .Y(_15320_));
NAND_g _21450_ (.A(_00011_[2]), .B(_15320_), .Y(_15321_));
NAND_g _21451_ (.A(cpuregs_10[15]), .B(_11217_), .Y(_15322_));
NAND_g _21452_ (.A(cpuregs_11[15]), .B(_00011_[0]), .Y(_15323_));
NAND_g _21453_ (.A(_15322_), .B(_15323_), .Y(_15324_));
NAND_g _21454_ (.A(_11219_), .B(_15324_), .Y(_15325_));
NAND_g _21455_ (.A(_15321_), .B(_15325_), .Y(_15326_));
NAND_g _21456_ (.A(_00011_[3]), .B(_15326_), .Y(_15327_));
NAND_g _21457_ (.A(cpuregs_6[15]), .B(_11217_), .Y(_15328_));
NAND_g _21458_ (.A(cpuregs_7[15]), .B(_00011_[0]), .Y(_15329_));
NAND_g _21459_ (.A(_15328_), .B(_15329_), .Y(_15330_));
NAND_g _21460_ (.A(_00011_[2]), .B(_15330_), .Y(_15331_));
NAND_g _21461_ (.A(cpuregs_2[15]), .B(_11217_), .Y(_15332_));
NAND_g _21462_ (.A(cpuregs_3[15]), .B(_00011_[0]), .Y(_15333_));
NAND_g _21463_ (.A(_15332_), .B(_15333_), .Y(_15334_));
NAND_g _21464_ (.A(_11219_), .B(_15334_), .Y(_15335_));
NAND_g _21465_ (.A(_15331_), .B(_15335_), .Y(_15336_));
NAND_g _21466_ (.A(_11220_), .B(_15336_), .Y(_15337_));
NAND_g _21467_ (.A(_15327_), .B(_15337_), .Y(_15338_));
NAND_g _21468_ (.A(_00011_[1]), .B(_15338_), .Y(_15339_));
NOR_g _21469_ (.A(cpuregs_9[15]), .B(_00011_[2]), .Y(_15340_));
NOT_g _21470_ (.A(_15340_), .Y(_15341_));
NAND_g _21471_ (.A(_11148_), .B(_00011_[2]), .Y(_15342_));
AND_g _21472_ (.A(_00011_[0]), .B(_15342_), .Y(_15343_));
NAND_g _21473_ (.A(_15341_), .B(_15343_), .Y(_15344_));
NOR_g _21474_ (.A(cpuregs_8[15]), .B(_00011_[2]), .Y(_15345_));
AND_g _21475_ (.A(_11119_), .B(_00011_[2]), .Y(_15346_));
NOR_g _21476_ (.A(_15345_), .B(_15346_), .Y(_15347_));
NAND_g _21477_ (.A(_11217_), .B(_15347_), .Y(_15348_));
NAND_g _21478_ (.A(_15344_), .B(_15348_), .Y(_15349_));
NAND_g _21479_ (.A(_00011_[3]), .B(_15349_), .Y(_15350_));
NAND_g _21480_ (.A(cpuregs_4[15]), .B(_00011_[2]), .Y(_15351_));
NAND_g _21481_ (.A(cpuregs_0[15]), .B(_11219_), .Y(_15352_));
AND_g _21482_ (.A(_15351_), .B(_15352_), .Y(_15353_));
NAND_g _21483_ (.A(_11217_), .B(_15353_), .Y(_15354_));
NAND_g _21484_ (.A(cpuregs_5[15]), .B(_00011_[2]), .Y(_15355_));
NAND_g _21485_ (.A(cpuregs_1[15]), .B(_11219_), .Y(_15356_));
AND_g _21486_ (.A(_00011_[0]), .B(_15356_), .Y(_15357_));
NAND_g _21487_ (.A(_15355_), .B(_15357_), .Y(_15358_));
AND_g _21488_ (.A(_11220_), .B(_15358_), .Y(_15359_));
NAND_g _21489_ (.A(_15354_), .B(_15359_), .Y(_15360_));
NAND_g _21490_ (.A(_15350_), .B(_15360_), .Y(_15361_));
NAND_g _21491_ (.A(_11218_), .B(_15361_), .Y(_15362_));
NAND_g _21492_ (.A(_15339_), .B(_15362_), .Y(_15363_));
AND_g _21493_ (.A(_00011_[4]), .B(_15295_), .Y(_15364_));
AND_g _21494_ (.A(_15317_), .B(_15364_), .Y(_15365_));
NOR_g _21495_ (.A(_00011_[4]), .B(_15363_), .Y(_15366_));
NOR_g _21496_ (.A(_15365_), .B(_15366_), .Y(_15367_));
AND_g _21497_ (.A(_13734_), .B(_15367_), .Y(_15368_));
NAND_g _21498_ (.A(_14358_), .B(_15368_), .Y(_15369_));
AND_g _21499_ (.A(decoded_imm[15]), .B(_13830_), .Y(_15370_));
NAND_g _21500_ (.A(_13409_), .B(_15370_), .Y(_15371_));
AND_g _21501_ (.A(_13727_), .B(_15371_), .Y(_15372_));
NAND_g _21502_ (.A(_15369_), .B(_15372_), .Y(_15373_));
AND_g _21503_ (.A(_15273_), .B(_15373_), .Y(_00518_));
NAND_g _21504_ (.A(_10996_), .B(_13728_), .Y(_15374_));
NAND_g _21505_ (.A(cpuregs_29[16]), .B(_00011_[2]), .Y(_15375_));
NAND_g _21506_ (.A(cpuregs_25[16]), .B(_11219_), .Y(_15376_));
AND_g _21507_ (.A(_00011_[0]), .B(_15376_), .Y(_15377_));
NAND_g _21508_ (.A(_15375_), .B(_15377_), .Y(_15378_));
NAND_g _21509_ (.A(cpuregs_24[16]), .B(_11219_), .Y(_15379_));
NAND_g _21510_ (.A(cpuregs_28[16]), .B(_00011_[2]), .Y(_15380_));
AND_g _21511_ (.A(_11217_), .B(_15380_), .Y(_15381_));
NAND_g _21512_ (.A(_15379_), .B(_15381_), .Y(_15382_));
AND_g _21513_ (.A(_11218_), .B(_15382_), .Y(_15383_));
NAND_g _21514_ (.A(_15378_), .B(_15383_), .Y(_15384_));
NAND_g _21515_ (.A(cpuregs_27[16]), .B(_11219_), .Y(_15385_));
NAND_g _21516_ (.A(cpuregs_31[16]), .B(_00011_[2]), .Y(_15386_));
AND_g _21517_ (.A(_00011_[0]), .B(_15386_), .Y(_15387_));
NAND_g _21518_ (.A(_15385_), .B(_15387_), .Y(_15388_));
NAND_g _21519_ (.A(cpuregs_26[16]), .B(_11219_), .Y(_15389_));
NAND_g _21520_ (.A(cpuregs_30[16]), .B(_00011_[2]), .Y(_15390_));
AND_g _21521_ (.A(_11217_), .B(_15390_), .Y(_15391_));
NAND_g _21522_ (.A(_15389_), .B(_15391_), .Y(_15392_));
AND_g _21523_ (.A(_00011_[1]), .B(_15392_), .Y(_15393_));
NAND_g _21524_ (.A(_15388_), .B(_15393_), .Y(_15394_));
NAND_g _21525_ (.A(_15384_), .B(_15394_), .Y(_15395_));
NAND_g _21526_ (.A(_00011_[4]), .B(_15395_), .Y(_15396_));
NAND_g _21527_ (.A(cpuregs_14[16]), .B(_11217_), .Y(_15397_));
NAND_g _21528_ (.A(cpuregs_15[16]), .B(_00011_[0]), .Y(_15398_));
NAND_g _21529_ (.A(_15397_), .B(_15398_), .Y(_15399_));
NAND_g _21530_ (.A(_00011_[2]), .B(_15399_), .Y(_15400_));
NAND_g _21531_ (.A(cpuregs_10[16]), .B(_11217_), .Y(_15401_));
NAND_g _21532_ (.A(cpuregs_11[16]), .B(_00011_[0]), .Y(_15402_));
NAND_g _21533_ (.A(_15401_), .B(_15402_), .Y(_15403_));
NAND_g _21534_ (.A(_11219_), .B(_15403_), .Y(_15404_));
NAND_g _21535_ (.A(_15400_), .B(_15404_), .Y(_15405_));
NAND_g _21536_ (.A(_00011_[1]), .B(_15405_), .Y(_15406_));
NAND_g _21537_ (.A(cpuregs_12[16]), .B(_11217_), .Y(_15407_));
NAND_g _21538_ (.A(cpuregs_13[16]), .B(_00011_[0]), .Y(_15408_));
NAND_g _21539_ (.A(_15407_), .B(_15408_), .Y(_15409_));
NAND_g _21540_ (.A(_00011_[2]), .B(_15409_), .Y(_15410_));
NAND_g _21541_ (.A(cpuregs_8[16]), .B(_11217_), .Y(_15411_));
NAND_g _21542_ (.A(cpuregs_9[16]), .B(_00011_[0]), .Y(_15412_));
NAND_g _21543_ (.A(_15411_), .B(_15412_), .Y(_15413_));
NAND_g _21544_ (.A(_11219_), .B(_15413_), .Y(_15414_));
NAND_g _21545_ (.A(_15410_), .B(_15414_), .Y(_15415_));
NAND_g _21546_ (.A(_11218_), .B(_15415_), .Y(_15416_));
NAND_g _21547_ (.A(_15406_), .B(_15416_), .Y(_15417_));
NAND_g _21548_ (.A(_11221_), .B(_15417_), .Y(_15418_));
NAND_g _21549_ (.A(_15396_), .B(_15418_), .Y(_15419_));
NAND_g _21550_ (.A(_00011_[3]), .B(_15419_), .Y(_15420_));
NAND_g _21551_ (.A(cpuregs_1[16]), .B(_11219_), .Y(_15421_));
NAND_g _21552_ (.A(cpuregs_5[16]), .B(_00011_[2]), .Y(_15422_));
AND_g _21553_ (.A(_00011_[0]), .B(_15422_), .Y(_15423_));
NAND_g _21554_ (.A(_15421_), .B(_15423_), .Y(_15424_));
NAND_g _21555_ (.A(cpuregs_0[16]), .B(_11219_), .Y(_15425_));
NAND_g _21556_ (.A(cpuregs_4[16]), .B(_00011_[2]), .Y(_15426_));
AND_g _21557_ (.A(_11217_), .B(_15426_), .Y(_15427_));
NAND_g _21558_ (.A(_15425_), .B(_15427_), .Y(_15428_));
AND_g _21559_ (.A(_11218_), .B(_15428_), .Y(_15429_));
NAND_g _21560_ (.A(_15424_), .B(_15429_), .Y(_15430_));
NAND_g _21561_ (.A(cpuregs_3[16]), .B(_11219_), .Y(_15431_));
NAND_g _21562_ (.A(cpuregs_7[16]), .B(_00011_[2]), .Y(_15432_));
AND_g _21563_ (.A(_00011_[0]), .B(_15432_), .Y(_15433_));
NAND_g _21564_ (.A(_15431_), .B(_15433_), .Y(_15434_));
NAND_g _21565_ (.A(cpuregs_2[16]), .B(_11219_), .Y(_15435_));
NAND_g _21566_ (.A(cpuregs_6[16]), .B(_00011_[2]), .Y(_15436_));
AND_g _21567_ (.A(_11217_), .B(_15436_), .Y(_15437_));
NAND_g _21568_ (.A(_15435_), .B(_15437_), .Y(_15438_));
AND_g _21569_ (.A(_00011_[1]), .B(_15438_), .Y(_15439_));
NAND_g _21570_ (.A(_15434_), .B(_15439_), .Y(_15440_));
NAND_g _21571_ (.A(_15430_), .B(_15440_), .Y(_15441_));
NAND_g _21572_ (.A(_11221_), .B(_15441_), .Y(_15442_));
NAND_g _21573_ (.A(cpuregs_19[16]), .B(_00011_[1]), .Y(_15443_));
NAND_g _21574_ (.A(cpuregs_17[16]), .B(_11218_), .Y(_15444_));
NAND_g _21575_ (.A(_15443_), .B(_15444_), .Y(_15445_));
NAND_g _21576_ (.A(_11219_), .B(_15445_), .Y(_15446_));
NAND_g _21577_ (.A(cpuregs_23[16]), .B(_00011_[1]), .Y(_15447_));
NAND_g _21578_ (.A(cpuregs_21[16]), .B(_11218_), .Y(_15448_));
NAND_g _21579_ (.A(_15447_), .B(_15448_), .Y(_15449_));
NAND_g _21580_ (.A(_00011_[2]), .B(_15449_), .Y(_15450_));
AND_g _21581_ (.A(_00011_[0]), .B(_15450_), .Y(_15451_));
NAND_g _21582_ (.A(_15446_), .B(_15451_), .Y(_15452_));
NAND_g _21583_ (.A(cpuregs_18[16]), .B(_00011_[1]), .Y(_15453_));
NAND_g _21584_ (.A(cpuregs_16[16]), .B(_11218_), .Y(_15454_));
NAND_g _21585_ (.A(_15453_), .B(_15454_), .Y(_15455_));
NAND_g _21586_ (.A(_11219_), .B(_15455_), .Y(_15456_));
NAND_g _21587_ (.A(cpuregs_22[16]), .B(_00011_[1]), .Y(_15457_));
NAND_g _21588_ (.A(cpuregs_20[16]), .B(_11218_), .Y(_15458_));
NAND_g _21589_ (.A(_15457_), .B(_15458_), .Y(_15459_));
NAND_g _21590_ (.A(_00011_[2]), .B(_15459_), .Y(_15460_));
AND_g _21591_ (.A(_11217_), .B(_15460_), .Y(_15461_));
NAND_g _21592_ (.A(_15456_), .B(_15461_), .Y(_15462_));
AND_g _21593_ (.A(_00011_[4]), .B(_15462_), .Y(_15463_));
NAND_g _21594_ (.A(_15452_), .B(_15463_), .Y(_15464_));
NAND_g _21595_ (.A(_15442_), .B(_15464_), .Y(_15465_));
NAND_g _21596_ (.A(_11220_), .B(_15465_), .Y(_15466_));
NAND_g _21597_ (.A(_15420_), .B(_15466_), .Y(_15467_));
AND_g _21598_ (.A(_13734_), .B(_15467_), .Y(_15468_));
NAND_g _21599_ (.A(_14358_), .B(_15468_), .Y(_15469_));
AND_g _21600_ (.A(decoded_imm[16]), .B(_13830_), .Y(_15470_));
NAND_g _21601_ (.A(_13409_), .B(_15470_), .Y(_15471_));
AND_g _21602_ (.A(_13727_), .B(_15471_), .Y(_15472_));
NAND_g _21603_ (.A(_15469_), .B(_15472_), .Y(_15473_));
AND_g _21604_ (.A(_15374_), .B(_15473_), .Y(_00519_));
NAND_g _21605_ (.A(_10997_), .B(_13728_), .Y(_15474_));
NAND_g _21606_ (.A(cpuregs_19[17]), .B(_11219_), .Y(_15475_));
NAND_g _21607_ (.A(cpuregs_23[17]), .B(_00011_[2]), .Y(_15476_));
AND_g _21608_ (.A(_00011_[0]), .B(_15476_), .Y(_15477_));
NAND_g _21609_ (.A(_15475_), .B(_15477_), .Y(_15478_));
NAND_g _21610_ (.A(cpuregs_18[17]), .B(_11219_), .Y(_15479_));
NAND_g _21611_ (.A(cpuregs_22[17]), .B(_00011_[2]), .Y(_15480_));
AND_g _21612_ (.A(_11217_), .B(_15480_), .Y(_15481_));
NAND_g _21613_ (.A(_15479_), .B(_15481_), .Y(_15482_));
AND_g _21614_ (.A(_11220_), .B(_15482_), .Y(_15483_));
NAND_g _21615_ (.A(_15478_), .B(_15483_), .Y(_15484_));
NAND_g _21616_ (.A(cpuregs_27[17]), .B(_11219_), .Y(_15485_));
NAND_g _21617_ (.A(cpuregs_31[17]), .B(_00011_[2]), .Y(_15486_));
AND_g _21618_ (.A(_00011_[0]), .B(_15486_), .Y(_15487_));
NAND_g _21619_ (.A(_15485_), .B(_15487_), .Y(_15488_));
NAND_g _21620_ (.A(cpuregs_26[17]), .B(_11219_), .Y(_15489_));
NAND_g _21621_ (.A(cpuregs_30[17]), .B(_00011_[2]), .Y(_15490_));
AND_g _21622_ (.A(_11217_), .B(_15490_), .Y(_15491_));
NAND_g _21623_ (.A(_15489_), .B(_15491_), .Y(_15492_));
AND_g _21624_ (.A(_00011_[3]), .B(_15492_), .Y(_15493_));
NAND_g _21625_ (.A(_15488_), .B(_15493_), .Y(_15494_));
NAND_g _21626_ (.A(_15484_), .B(_15494_), .Y(_15495_));
NAND_g _21627_ (.A(_00011_[1]), .B(_15495_), .Y(_15496_));
NOR_g _21628_ (.A(cpuregs_16[17]), .B(_00011_[2]), .Y(_15497_));
AND_g _21629_ (.A(_11198_), .B(_00011_[2]), .Y(_15498_));
NOR_g _21630_ (.A(_15497_), .B(_15498_), .Y(_15499_));
NOR_g _21631_ (.A(cpuregs_17[17]), .B(_00011_[2]), .Y(_15500_));
NAND_g _21632_ (.A(_11031_), .B(_00011_[2]), .Y(_15501_));
NOR_g _21633_ (.A(cpuregs_24[17]), .B(_00011_[2]), .Y(_15502_));
AND_g _21634_ (.A(_11098_), .B(_00011_[2]), .Y(_15503_));
NOR_g _21635_ (.A(_15502_), .B(_15503_), .Y(_15504_));
NOR_g _21636_ (.A(cpuregs_25[17]), .B(_00011_[2]), .Y(_15505_));
NAND_g _21637_ (.A(_10930_), .B(_00011_[2]), .Y(_15506_));
NAND_g _21638_ (.A(_11217_), .B(_15499_), .Y(_15507_));
NOR_g _21639_ (.A(_11217_), .B(_15500_), .Y(_15508_));
NAND_g _21640_ (.A(_15501_), .B(_15508_), .Y(_15509_));
AND_g _21641_ (.A(_15507_), .B(_15509_), .Y(_15510_));
NAND_g _21642_ (.A(_11220_), .B(_15510_), .Y(_15511_));
NOR_g _21643_ (.A(_11217_), .B(_15505_), .Y(_15512_));
NAND_g _21644_ (.A(_15506_), .B(_15512_), .Y(_15513_));
NAND_g _21645_ (.A(_11217_), .B(_15504_), .Y(_15514_));
AND_g _21646_ (.A(_15513_), .B(_15514_), .Y(_15515_));
NAND_g _21647_ (.A(_00011_[3]), .B(_15515_), .Y(_15516_));
AND_g _21648_ (.A(_15511_), .B(_15516_), .Y(_15517_));
NAND_g _21649_ (.A(_11218_), .B(_15517_), .Y(_15518_));
NAND_g _21650_ (.A(cpuregs_6[17]), .B(_00011_[2]), .Y(_15519_));
NAND_g _21651_ (.A(cpuregs_2[17]), .B(_11219_), .Y(_15520_));
AND_g _21652_ (.A(_15519_), .B(_15520_), .Y(_15521_));
NAND_g _21653_ (.A(_11217_), .B(_15521_), .Y(_15522_));
NAND_g _21654_ (.A(cpuregs_7[17]), .B(_00011_[2]), .Y(_15523_));
NAND_g _21655_ (.A(cpuregs_3[17]), .B(_11219_), .Y(_15524_));
AND_g _21656_ (.A(_00011_[0]), .B(_15524_), .Y(_15525_));
NAND_g _21657_ (.A(_15523_), .B(_15525_), .Y(_15526_));
AND_g _21658_ (.A(_11220_), .B(_15526_), .Y(_15527_));
NAND_g _21659_ (.A(_15522_), .B(_15527_), .Y(_15528_));
NOR_g _21660_ (.A(cpuregs_10[17]), .B(_00011_[2]), .Y(_15529_));
NOR_g _21661_ (.A(cpuregs_14[17]), .B(_11219_), .Y(_15530_));
NOR_g _21662_ (.A(_15529_), .B(_15530_), .Y(_15531_));
NOR_g _21663_ (.A(cpuregs_11[17]), .B(_00011_[2]), .Y(_15532_));
NOT_g _21664_ (.A(_15532_), .Y(_15533_));
NAND_g _21665_ (.A(_11165_), .B(_00011_[2]), .Y(_15534_));
AND_g _21666_ (.A(_00011_[0]), .B(_15534_), .Y(_15535_));
NAND_g _21667_ (.A(_15533_), .B(_15535_), .Y(_15536_));
NAND_g _21668_ (.A(_11217_), .B(_15531_), .Y(_15537_));
NAND_g _21669_ (.A(_15536_), .B(_15537_), .Y(_15538_));
NAND_g _21670_ (.A(_00011_[3]), .B(_15538_), .Y(_15539_));
NAND_g _21671_ (.A(_15528_), .B(_15539_), .Y(_15540_));
NAND_g _21672_ (.A(_00011_[1]), .B(_15540_), .Y(_15541_));
NAND_g _21673_ (.A(cpuregs_4[17]), .B(_00011_[2]), .Y(_15542_));
NAND_g _21674_ (.A(cpuregs_0[17]), .B(_11219_), .Y(_15543_));
AND_g _21675_ (.A(_11217_), .B(_15543_), .Y(_15544_));
NAND_g _21676_ (.A(_15542_), .B(_15544_), .Y(_15545_));
NAND_g _21677_ (.A(cpuregs_1[17]), .B(_11219_), .Y(_15546_));
NAND_g _21678_ (.A(cpuregs_5[17]), .B(_00011_[2]), .Y(_15547_));
AND_g _21679_ (.A(_00011_[0]), .B(_15547_), .Y(_15548_));
NAND_g _21680_ (.A(_15546_), .B(_15548_), .Y(_15549_));
NOR_g _21681_ (.A(cpuregs_9[17]), .B(_00011_[2]), .Y(_15550_));
NAND_g _21682_ (.A(_11149_), .B(_00011_[2]), .Y(_15551_));
NOR_g _21683_ (.A(cpuregs_8[17]), .B(_00011_[2]), .Y(_15552_));
NOR_g _21684_ (.A(cpuregs_12[17]), .B(_11219_), .Y(_15553_));
NOR_g _21685_ (.A(_15552_), .B(_15553_), .Y(_15554_));
NAND_g _21686_ (.A(_15545_), .B(_15549_), .Y(_15555_));
NAND_g _21687_ (.A(_11220_), .B(_15555_), .Y(_15556_));
NAND_g _21688_ (.A(_11217_), .B(_15554_), .Y(_15557_));
NOR_g _21689_ (.A(_11217_), .B(_15550_), .Y(_15558_));
NAND_g _21690_ (.A(_15551_), .B(_15558_), .Y(_15559_));
AND_g _21691_ (.A(_00011_[3]), .B(_15559_), .Y(_15560_));
NAND_g _21692_ (.A(_15557_), .B(_15560_), .Y(_15561_));
AND_g _21693_ (.A(_15556_), .B(_15561_), .Y(_15562_));
NAND_g _21694_ (.A(_11218_), .B(_15562_), .Y(_15563_));
AND_g _21695_ (.A(_15541_), .B(_15563_), .Y(_15564_));
AND_g _21696_ (.A(_00011_[4]), .B(_15496_), .Y(_15565_));
NAND_g _21697_ (.A(_15518_), .B(_15565_), .Y(_15566_));
NAND_g _21698_ (.A(_11221_), .B(_15564_), .Y(_15567_));
AND_g _21699_ (.A(_15566_), .B(_15567_), .Y(_15568_));
AND_g _21700_ (.A(_13734_), .B(_15568_), .Y(_15569_));
NAND_g _21701_ (.A(_14358_), .B(_15569_), .Y(_15570_));
AND_g _21702_ (.A(decoded_imm[17]), .B(_13830_), .Y(_15571_));
NAND_g _21703_ (.A(_13409_), .B(_15571_), .Y(_15572_));
AND_g _21704_ (.A(_13727_), .B(_15572_), .Y(_15573_));
NAND_g _21705_ (.A(_15570_), .B(_15573_), .Y(_15574_));
AND_g _21706_ (.A(_15474_), .B(_15574_), .Y(_00520_));
NAND_g _21707_ (.A(_10998_), .B(_13728_), .Y(_15575_));
NAND_g _21708_ (.A(_10931_), .B(_00011_[2]), .Y(_15576_));
NOR_g _21709_ (.A(cpuregs_25[18]), .B(_00011_[2]), .Y(_15577_));
NAND_g _21710_ (.A(_00011_[0]), .B(_15576_), .Y(_15578_));
NOR_g _21711_ (.A(_15577_), .B(_15578_), .Y(_15579_));
NOR_g _21712_ (.A(cpuregs_24[18]), .B(_00011_[2]), .Y(_15580_));
AND_g _21713_ (.A(_11099_), .B(_00011_[2]), .Y(_15581_));
NOR_g _21714_ (.A(_15580_), .B(_15581_), .Y(_15582_));
AND_g _21715_ (.A(_11217_), .B(_15582_), .Y(_15583_));
NOR_g _21716_ (.A(_15579_), .B(_15583_), .Y(_15584_));
NAND_g _21717_ (.A(_11218_), .B(_15584_), .Y(_15585_));
NOR_g _21718_ (.A(cpuregs_26[18]), .B(_00011_[2]), .Y(_15586_));
AND_g _21719_ (.A(_11175_), .B(_00011_[2]), .Y(_15587_));
NOR_g _21720_ (.A(_15586_), .B(_15587_), .Y(_15588_));
AND_g _21721_ (.A(_11217_), .B(_15588_), .Y(_15589_));
NAND_g _21722_ (.A(_11091_), .B(_00011_[2]), .Y(_15590_));
NOR_g _21723_ (.A(cpuregs_27[18]), .B(_00011_[2]), .Y(_15591_));
NAND_g _21724_ (.A(_00011_[0]), .B(_15590_), .Y(_15592_));
NOR_g _21725_ (.A(_15591_), .B(_15592_), .Y(_15593_));
NOR_g _21726_ (.A(_15589_), .B(_15593_), .Y(_15594_));
NAND_g _21727_ (.A(_00011_[1]), .B(_15594_), .Y(_15595_));
AND_g _21728_ (.A(_00011_[3]), .B(_15585_), .Y(_15596_));
NAND_g _21729_ (.A(_15595_), .B(_15596_), .Y(_15597_));
NOR_g _21730_ (.A(cpuregs_18[18]), .B(_00011_[2]), .Y(_15598_));
AND_g _21731_ (.A(_11018_), .B(_00011_[2]), .Y(_15599_));
NOR_g _21732_ (.A(_15598_), .B(_15599_), .Y(_15600_));
NOR_g _21733_ (.A(cpuregs_16[18]), .B(_00011_[2]), .Y(_15601_));
AND_g _21734_ (.A(_11199_), .B(_00011_[2]), .Y(_15602_));
NOR_g _21735_ (.A(_15601_), .B(_15602_), .Y(_15603_));
NAND_g _21736_ (.A(_11185_), .B(_00011_[2]), .Y(_15604_));
NOR_g _21737_ (.A(cpuregs_19[18]), .B(_00011_[2]), .Y(_15605_));
NOR_g _21738_ (.A(cpuregs_17[18]), .B(_00011_[2]), .Y(_15606_));
NAND_g _21739_ (.A(_11032_), .B(_00011_[2]), .Y(_15607_));
NOR_g _21740_ (.A(_11217_), .B(_15605_), .Y(_15608_));
NAND_g _21741_ (.A(_15604_), .B(_15608_), .Y(_15609_));
NAND_g _21742_ (.A(_11217_), .B(_15600_), .Y(_15610_));
AND_g _21743_ (.A(_15609_), .B(_15610_), .Y(_15611_));
NAND_g _21744_ (.A(_00011_[1]), .B(_15611_), .Y(_15612_));
NOR_g _21745_ (.A(_11217_), .B(_15606_), .Y(_15613_));
NAND_g _21746_ (.A(_15607_), .B(_15613_), .Y(_15614_));
NAND_g _21747_ (.A(_11217_), .B(_15603_), .Y(_15615_));
AND_g _21748_ (.A(_15614_), .B(_15615_), .Y(_15616_));
NAND_g _21749_ (.A(_11218_), .B(_15616_), .Y(_15617_));
AND_g _21750_ (.A(_15612_), .B(_15617_), .Y(_15618_));
NAND_g _21751_ (.A(_11220_), .B(_15618_), .Y(_15619_));
NAND_g _21752_ (.A(_15597_), .B(_15619_), .Y(_15620_));
NAND_g _21753_ (.A(_00011_[4]), .B(_15620_), .Y(_15621_));
NAND_g _21754_ (.A(cpuregs_13[18]), .B(_11218_), .Y(_15622_));
NAND_g _21755_ (.A(cpuregs_15[18]), .B(_00011_[1]), .Y(_15623_));
AND_g _21756_ (.A(_00011_[2]), .B(_15623_), .Y(_15624_));
NAND_g _21757_ (.A(_15622_), .B(_15624_), .Y(_15625_));
NAND_g _21758_ (.A(cpuregs_9[18]), .B(_11218_), .Y(_15626_));
NAND_g _21759_ (.A(cpuregs_11[18]), .B(_00011_[1]), .Y(_15627_));
AND_g _21760_ (.A(_11219_), .B(_15627_), .Y(_15628_));
NAND_g _21761_ (.A(_15626_), .B(_15628_), .Y(_15629_));
AND_g _21762_ (.A(_00011_[0]), .B(_15629_), .Y(_15630_));
NAND_g _21763_ (.A(_15625_), .B(_15630_), .Y(_15631_));
NAND_g _21764_ (.A(cpuregs_12[18]), .B(_11218_), .Y(_15632_));
NAND_g _21765_ (.A(cpuregs_14[18]), .B(_00011_[1]), .Y(_15633_));
AND_g _21766_ (.A(_00011_[2]), .B(_15633_), .Y(_15634_));
NAND_g _21767_ (.A(_15632_), .B(_15634_), .Y(_15635_));
NAND_g _21768_ (.A(cpuregs_8[18]), .B(_11218_), .Y(_15636_));
NAND_g _21769_ (.A(cpuregs_10[18]), .B(_00011_[1]), .Y(_15637_));
AND_g _21770_ (.A(_11219_), .B(_15637_), .Y(_15638_));
NAND_g _21771_ (.A(_15636_), .B(_15638_), .Y(_15639_));
AND_g _21772_ (.A(_11217_), .B(_15639_), .Y(_15640_));
NAND_g _21773_ (.A(_15635_), .B(_15640_), .Y(_15641_));
NAND_g _21774_ (.A(_15631_), .B(_15641_), .Y(_15642_));
NAND_g _21775_ (.A(_00011_[3]), .B(_15642_), .Y(_15643_));
NAND_g _21776_ (.A(_10944_), .B(_00011_[2]), .Y(_15644_));
NOR_g _21777_ (.A(cpuregs_2[18]), .B(_00011_[2]), .Y(_15645_));
NOR_g _21778_ (.A(_00011_[0]), .B(_15645_), .Y(_15646_));
NAND_g _21779_ (.A(_15644_), .B(_15646_), .Y(_15647_));
NAND_g _21780_ (.A(_11130_), .B(_00011_[2]), .Y(_15648_));
NOR_g _21781_ (.A(cpuregs_3[18]), .B(_00011_[2]), .Y(_15649_));
NOR_g _21782_ (.A(_11217_), .B(_15649_), .Y(_15650_));
NAND_g _21783_ (.A(_15648_), .B(_15650_), .Y(_15651_));
AND_g _21784_ (.A(_15647_), .B(_15651_), .Y(_15652_));
NAND_g _21785_ (.A(_10956_), .B(_00011_[2]), .Y(_15653_));
NOR_g _21786_ (.A(cpuregs_0[18]), .B(_00011_[2]), .Y(_15654_));
NOR_g _21787_ (.A(_00011_[0]), .B(_15654_), .Y(_15655_));
NAND_g _21788_ (.A(_15653_), .B(_15655_), .Y(_15656_));
NAND_g _21789_ (.A(_11114_), .B(_00011_[2]), .Y(_15657_));
NOR_g _21790_ (.A(cpuregs_1[18]), .B(_00011_[2]), .Y(_15658_));
NOR_g _21791_ (.A(_11217_), .B(_15658_), .Y(_15659_));
NAND_g _21792_ (.A(_15657_), .B(_15659_), .Y(_15660_));
AND_g _21793_ (.A(_15656_), .B(_15660_), .Y(_15661_));
NAND_g _21794_ (.A(_00011_[1]), .B(_15652_), .Y(_15662_));
NAND_g _21795_ (.A(_11218_), .B(_15661_), .Y(_15663_));
AND_g _21796_ (.A(_15662_), .B(_15663_), .Y(_15664_));
NAND_g _21797_ (.A(_11220_), .B(_15664_), .Y(_15665_));
NAND_g _21798_ (.A(_15643_), .B(_15665_), .Y(_15666_));
NAND_g _21799_ (.A(_11221_), .B(_15666_), .Y(_15667_));
NAND_g _21800_ (.A(_15621_), .B(_15667_), .Y(_15668_));
AND_g _21801_ (.A(_13734_), .B(_15668_), .Y(_15669_));
NAND_g _21802_ (.A(_14358_), .B(_15669_), .Y(_15670_));
AND_g _21803_ (.A(decoded_imm[18]), .B(_13830_), .Y(_15671_));
NAND_g _21804_ (.A(_13409_), .B(_15671_), .Y(_15672_));
AND_g _21805_ (.A(_13727_), .B(_15672_), .Y(_15673_));
NAND_g _21806_ (.A(_15670_), .B(_15673_), .Y(_15674_));
AND_g _21807_ (.A(_15575_), .B(_15674_), .Y(_00521_));
NAND_g _21808_ (.A(_10999_), .B(_13728_), .Y(_15675_));
NAND_g _21809_ (.A(cpuregs_19[19]), .B(_11219_), .Y(_15676_));
NAND_g _21810_ (.A(cpuregs_23[19]), .B(_00011_[2]), .Y(_15677_));
AND_g _21811_ (.A(_00011_[0]), .B(_15677_), .Y(_15678_));
NAND_g _21812_ (.A(_15676_), .B(_15678_), .Y(_15679_));
NAND_g _21813_ (.A(cpuregs_18[19]), .B(_11219_), .Y(_15680_));
NAND_g _21814_ (.A(cpuregs_22[19]), .B(_00011_[2]), .Y(_15681_));
AND_g _21815_ (.A(_11217_), .B(_15681_), .Y(_15682_));
NAND_g _21816_ (.A(_15680_), .B(_15682_), .Y(_15683_));
AND_g _21817_ (.A(_11220_), .B(_15683_), .Y(_15684_));
NAND_g _21818_ (.A(_15679_), .B(_15684_), .Y(_15685_));
NAND_g _21819_ (.A(cpuregs_27[19]), .B(_11219_), .Y(_15686_));
NAND_g _21820_ (.A(cpuregs_31[19]), .B(_00011_[2]), .Y(_15687_));
AND_g _21821_ (.A(_00011_[0]), .B(_15687_), .Y(_15688_));
NAND_g _21822_ (.A(_15686_), .B(_15688_), .Y(_15689_));
NAND_g _21823_ (.A(cpuregs_26[19]), .B(_11219_), .Y(_15690_));
NAND_g _21824_ (.A(cpuregs_30[19]), .B(_00011_[2]), .Y(_15691_));
AND_g _21825_ (.A(_11217_), .B(_15691_), .Y(_15692_));
NAND_g _21826_ (.A(_15690_), .B(_15692_), .Y(_15693_));
AND_g _21827_ (.A(_00011_[3]), .B(_15693_), .Y(_15694_));
NAND_g _21828_ (.A(_15689_), .B(_15694_), .Y(_15695_));
NAND_g _21829_ (.A(_15685_), .B(_15695_), .Y(_15696_));
NAND_g _21830_ (.A(_00011_[1]), .B(_15696_), .Y(_15697_));
NAND_g _21831_ (.A(cpuregs_21[19]), .B(_00011_[2]), .Y(_15698_));
NAND_g _21832_ (.A(cpuregs_17[19]), .B(_11219_), .Y(_15699_));
AND_g _21833_ (.A(_00011_[0]), .B(_15699_), .Y(_15700_));
NAND_g _21834_ (.A(_15698_), .B(_15700_), .Y(_15701_));
NAND_g _21835_ (.A(cpuregs_20[19]), .B(_00011_[2]), .Y(_15702_));
NAND_g _21836_ (.A(cpuregs_16[19]), .B(_11219_), .Y(_15703_));
AND_g _21837_ (.A(_11217_), .B(_15703_), .Y(_15704_));
NAND_g _21838_ (.A(_15702_), .B(_15704_), .Y(_15705_));
AND_g _21839_ (.A(_11220_), .B(_15705_), .Y(_15706_));
NAND_g _21840_ (.A(_15701_), .B(_15706_), .Y(_15707_));
NAND_g _21841_ (.A(cpuregs_25[19]), .B(_11219_), .Y(_15708_));
NAND_g _21842_ (.A(cpuregs_29[19]), .B(_00011_[2]), .Y(_15709_));
AND_g _21843_ (.A(_00011_[0]), .B(_15709_), .Y(_15710_));
NAND_g _21844_ (.A(_15708_), .B(_15710_), .Y(_15711_));
NAND_g _21845_ (.A(cpuregs_24[19]), .B(_11219_), .Y(_15712_));
NAND_g _21846_ (.A(cpuregs_28[19]), .B(_00011_[2]), .Y(_15713_));
AND_g _21847_ (.A(_11217_), .B(_15713_), .Y(_15714_));
NAND_g _21848_ (.A(_15712_), .B(_15714_), .Y(_15715_));
AND_g _21849_ (.A(_00011_[3]), .B(_15715_), .Y(_15716_));
NAND_g _21850_ (.A(_15711_), .B(_15716_), .Y(_15717_));
NAND_g _21851_ (.A(_15707_), .B(_15717_), .Y(_15718_));
NAND_g _21852_ (.A(_11218_), .B(_15718_), .Y(_15719_));
NAND_g _21853_ (.A(_15697_), .B(_15719_), .Y(_15720_));
NAND_g _21854_ (.A(_00011_[4]), .B(_15720_), .Y(_15721_));
NAND_g _21855_ (.A(cpuregs_6[19]), .B(_00011_[2]), .Y(_15722_));
NAND_g _21856_ (.A(cpuregs_2[19]), .B(_11219_), .Y(_15723_));
AND_g _21857_ (.A(_15722_), .B(_15723_), .Y(_15724_));
NAND_g _21858_ (.A(_11217_), .B(_15724_), .Y(_15725_));
NAND_g _21859_ (.A(cpuregs_7[19]), .B(_00011_[2]), .Y(_15726_));
NAND_g _21860_ (.A(cpuregs_3[19]), .B(_11219_), .Y(_15727_));
AND_g _21861_ (.A(_00011_[0]), .B(_15727_), .Y(_15728_));
NAND_g _21862_ (.A(_15726_), .B(_15728_), .Y(_15729_));
AND_g _21863_ (.A(_11220_), .B(_15729_), .Y(_15730_));
NAND_g _21864_ (.A(_15725_), .B(_15730_), .Y(_15731_));
NOR_g _21865_ (.A(cpuregs_10[19]), .B(_00011_[2]), .Y(_15732_));
AND_g _21866_ (.A(_11105_), .B(_00011_[2]), .Y(_15733_));
NOR_g _21867_ (.A(_15732_), .B(_15733_), .Y(_15734_));
NOR_g _21868_ (.A(cpuregs_11[19]), .B(_00011_[2]), .Y(_15735_));
NOT_g _21869_ (.A(_15735_), .Y(_15736_));
NAND_g _21870_ (.A(_11167_), .B(_00011_[2]), .Y(_15737_));
AND_g _21871_ (.A(_00011_[0]), .B(_15737_), .Y(_15738_));
NAND_g _21872_ (.A(_15736_), .B(_15738_), .Y(_15739_));
NAND_g _21873_ (.A(_11217_), .B(_15734_), .Y(_15740_));
NAND_g _21874_ (.A(_15739_), .B(_15740_), .Y(_15741_));
NAND_g _21875_ (.A(_00011_[3]), .B(_15741_), .Y(_15742_));
AND_g _21876_ (.A(_15731_), .B(_15742_), .Y(_15743_));
NAND_g _21877_ (.A(cpuregs_4[19]), .B(_00011_[2]), .Y(_15744_));
NAND_g _21878_ (.A(cpuregs_0[19]), .B(_11219_), .Y(_15745_));
AND_g _21879_ (.A(_15744_), .B(_15745_), .Y(_15746_));
NAND_g _21880_ (.A(_11217_), .B(_15746_), .Y(_15747_));
NAND_g _21881_ (.A(cpuregs_5[19]), .B(_00011_[2]), .Y(_15748_));
NAND_g _21882_ (.A(cpuregs_1[19]), .B(_11219_), .Y(_15749_));
AND_g _21883_ (.A(_00011_[0]), .B(_15749_), .Y(_15750_));
NAND_g _21884_ (.A(_15748_), .B(_15750_), .Y(_15751_));
AND_g _21885_ (.A(_11220_), .B(_15751_), .Y(_15752_));
AND_g _21886_ (.A(_15747_), .B(_15752_), .Y(_15753_));
NAND_g _21887_ (.A(_10934_), .B(_11219_), .Y(_15754_));
NAND_g _21888_ (.A(_11151_), .B(_00011_[2]), .Y(_15755_));
NOR_g _21889_ (.A(cpuregs_8[19]), .B(_00011_[2]), .Y(_15756_));
AND_g _21890_ (.A(_11121_), .B(_00011_[2]), .Y(_15757_));
NOR_g _21891_ (.A(_15756_), .B(_15757_), .Y(_15758_));
AND_g _21892_ (.A(_00011_[0]), .B(_15755_), .Y(_15759_));
NAND_g _21893_ (.A(_15754_), .B(_15759_), .Y(_15760_));
NAND_g _21894_ (.A(_11217_), .B(_15758_), .Y(_15761_));
NAND_g _21895_ (.A(_15760_), .B(_15761_), .Y(_15762_));
AND_g _21896_ (.A(_00011_[3]), .B(_15762_), .Y(_15763_));
NOR_g _21897_ (.A(_15753_), .B(_15763_), .Y(_15764_));
NAND_g _21898_ (.A(_11218_), .B(_15764_), .Y(_15765_));
NAND_g _21899_ (.A(_00011_[1]), .B(_15743_), .Y(_15766_));
AND_g _21900_ (.A(_15765_), .B(_15766_), .Y(_15767_));
NAND_g _21901_ (.A(_11221_), .B(_15767_), .Y(_15768_));
NAND_g _21902_ (.A(_15721_), .B(_15768_), .Y(_15769_));
AND_g _21903_ (.A(_13734_), .B(_15769_), .Y(_15770_));
NAND_g _21904_ (.A(_14358_), .B(_15770_), .Y(_15771_));
AND_g _21905_ (.A(decoded_imm[19]), .B(_13830_), .Y(_15772_));
NAND_g _21906_ (.A(_13409_), .B(_15772_), .Y(_15773_));
AND_g _21907_ (.A(_13727_), .B(_15773_), .Y(_15774_));
NAND_g _21908_ (.A(_15771_), .B(_15774_), .Y(_15775_));
AND_g _21909_ (.A(_15675_), .B(_15775_), .Y(_00522_));
NAND_g _21910_ (.A(_11000_), .B(_13728_), .Y(_15776_));
NAND_g _21911_ (.A(cpuregs_16[20]), .B(_11217_), .Y(_15777_));
NAND_g _21912_ (.A(cpuregs_17[20]), .B(_00011_[0]), .Y(_15778_));
AND_g _21913_ (.A(_11219_), .B(_15778_), .Y(_15779_));
NAND_g _21914_ (.A(_15777_), .B(_15779_), .Y(_15780_));
NAND_g _21915_ (.A(cpuregs_20[20]), .B(_11217_), .Y(_15781_));
NAND_g _21916_ (.A(cpuregs_21[20]), .B(_00011_[0]), .Y(_15782_));
AND_g _21917_ (.A(_00011_[2]), .B(_15782_), .Y(_15783_));
NAND_g _21918_ (.A(_15781_), .B(_15783_), .Y(_15784_));
NAND_g _21919_ (.A(_15780_), .B(_15784_), .Y(_15785_));
NAND_g _21920_ (.A(_11218_), .B(_15785_), .Y(_15786_));
NAND_g _21921_ (.A(cpuregs_18[20]), .B(_11217_), .Y(_15787_));
NAND_g _21922_ (.A(cpuregs_19[20]), .B(_00011_[0]), .Y(_15788_));
AND_g _21923_ (.A(_11219_), .B(_15788_), .Y(_15789_));
NAND_g _21924_ (.A(_15787_), .B(_15789_), .Y(_15790_));
NAND_g _21925_ (.A(cpuregs_22[20]), .B(_11217_), .Y(_15791_));
NAND_g _21926_ (.A(cpuregs_23[20]), .B(_00011_[0]), .Y(_15792_));
AND_g _21927_ (.A(_00011_[2]), .B(_15792_), .Y(_15793_));
NAND_g _21928_ (.A(_15791_), .B(_15793_), .Y(_15794_));
NAND_g _21929_ (.A(_15790_), .B(_15794_), .Y(_15795_));
NAND_g _21930_ (.A(_00011_[1]), .B(_15795_), .Y(_15796_));
AND_g _21931_ (.A(_11220_), .B(_15796_), .Y(_15797_));
NAND_g _21932_ (.A(_15786_), .B(_15797_), .Y(_15798_));
NOR_g _21933_ (.A(cpuregs_26[20]), .B(_00011_[2]), .Y(_15799_));
AND_g _21934_ (.A(_11176_), .B(_00011_[2]), .Y(_15800_));
NOR_g _21935_ (.A(_15799_), .B(_15800_), .Y(_15801_));
NAND_g _21936_ (.A(_11217_), .B(_15801_), .Y(_15802_));
NAND_g _21937_ (.A(_11092_), .B(_00011_[2]), .Y(_15803_));
NOR_g _21938_ (.A(cpuregs_27[20]), .B(_00011_[2]), .Y(_15804_));
NOR_g _21939_ (.A(_11217_), .B(_15804_), .Y(_15805_));
NAND_g _21940_ (.A(_15803_), .B(_15805_), .Y(_15806_));
AND_g _21941_ (.A(_15802_), .B(_15806_), .Y(_15807_));
NAND_g _21942_ (.A(_00011_[1]), .B(_15807_), .Y(_15808_));
NOR_g _21943_ (.A(cpuregs_24[20]), .B(_00011_[2]), .Y(_15809_));
AND_g _21944_ (.A(_11100_), .B(_00011_[2]), .Y(_15810_));
NOR_g _21945_ (.A(_15809_), .B(_15810_), .Y(_15811_));
NAND_g _21946_ (.A(_11217_), .B(_15811_), .Y(_15812_));
NAND_g _21947_ (.A(_10932_), .B(_00011_[2]), .Y(_15813_));
NOR_g _21948_ (.A(cpuregs_25[20]), .B(_00011_[2]), .Y(_15814_));
NOR_g _21949_ (.A(_11217_), .B(_15814_), .Y(_15815_));
AND_g _21950_ (.A(_15813_), .B(_15815_), .Y(_15816_));
NOR_g _21951_ (.A(_00011_[1]), .B(_15816_), .Y(_15817_));
NAND_g _21952_ (.A(_15812_), .B(_15817_), .Y(_15818_));
AND_g _21953_ (.A(_00011_[3]), .B(_15818_), .Y(_15819_));
NAND_g _21954_ (.A(_15808_), .B(_15819_), .Y(_15820_));
NAND_g _21955_ (.A(_15798_), .B(_15820_), .Y(_15821_));
NAND_g _21956_ (.A(_00011_[4]), .B(_15821_), .Y(_15822_));
NAND_g _21957_ (.A(cpuregs_13[20]), .B(_11218_), .Y(_15823_));
NAND_g _21958_ (.A(cpuregs_15[20]), .B(_00011_[1]), .Y(_15824_));
AND_g _21959_ (.A(_00011_[2]), .B(_15824_), .Y(_15825_));
NAND_g _21960_ (.A(_15823_), .B(_15825_), .Y(_15826_));
NAND_g _21961_ (.A(cpuregs_9[20]), .B(_11218_), .Y(_15827_));
NAND_g _21962_ (.A(cpuregs_11[20]), .B(_00011_[1]), .Y(_15828_));
AND_g _21963_ (.A(_11219_), .B(_15828_), .Y(_15829_));
NAND_g _21964_ (.A(_15827_), .B(_15829_), .Y(_15830_));
AND_g _21965_ (.A(_00011_[0]), .B(_15830_), .Y(_15831_));
NAND_g _21966_ (.A(_15826_), .B(_15831_), .Y(_15832_));
NAND_g _21967_ (.A(cpuregs_12[20]), .B(_11218_), .Y(_15833_));
NAND_g _21968_ (.A(cpuregs_14[20]), .B(_00011_[1]), .Y(_15834_));
AND_g _21969_ (.A(_00011_[2]), .B(_15834_), .Y(_15835_));
NAND_g _21970_ (.A(_15833_), .B(_15835_), .Y(_15836_));
NAND_g _21971_ (.A(cpuregs_8[20]), .B(_11218_), .Y(_15837_));
NAND_g _21972_ (.A(cpuregs_10[20]), .B(_00011_[1]), .Y(_15838_));
AND_g _21973_ (.A(_11219_), .B(_15838_), .Y(_15839_));
NAND_g _21974_ (.A(_15837_), .B(_15839_), .Y(_15840_));
AND_g _21975_ (.A(_11217_), .B(_15840_), .Y(_15841_));
NAND_g _21976_ (.A(_15836_), .B(_15841_), .Y(_15842_));
NAND_g _21977_ (.A(_15832_), .B(_15842_), .Y(_15843_));
NAND_g _21978_ (.A(_00011_[3]), .B(_15843_), .Y(_15844_));
NAND_g _21979_ (.A(_10945_), .B(_00011_[2]), .Y(_15845_));
NOR_g _21980_ (.A(cpuregs_2[20]), .B(_00011_[2]), .Y(_15846_));
NOR_g _21981_ (.A(_00011_[0]), .B(_15846_), .Y(_15847_));
NAND_g _21982_ (.A(_15845_), .B(_15847_), .Y(_15848_));
NAND_g _21983_ (.A(_11131_), .B(_00011_[2]), .Y(_15849_));
NOR_g _21984_ (.A(cpuregs_3[20]), .B(_00011_[2]), .Y(_15850_));
NOR_g _21985_ (.A(_11217_), .B(_15850_), .Y(_15851_));
NAND_g _21986_ (.A(_15849_), .B(_15851_), .Y(_15852_));
AND_g _21987_ (.A(_15848_), .B(_15852_), .Y(_15853_));
NAND_g _21988_ (.A(_10957_), .B(_00011_[2]), .Y(_15854_));
NOR_g _21989_ (.A(cpuregs_0[20]), .B(_00011_[2]), .Y(_15855_));
NOR_g _21990_ (.A(_00011_[0]), .B(_15855_), .Y(_15856_));
NAND_g _21991_ (.A(_15854_), .B(_15856_), .Y(_15857_));
NAND_g _21992_ (.A(_11115_), .B(_00011_[2]), .Y(_15858_));
NOR_g _21993_ (.A(cpuregs_1[20]), .B(_00011_[2]), .Y(_15859_));
NOR_g _21994_ (.A(_11217_), .B(_15859_), .Y(_15860_));
NAND_g _21995_ (.A(_15858_), .B(_15860_), .Y(_15861_));
AND_g _21996_ (.A(_15857_), .B(_15861_), .Y(_15862_));
NAND_g _21997_ (.A(_00011_[1]), .B(_15853_), .Y(_15863_));
NAND_g _21998_ (.A(_11218_), .B(_15862_), .Y(_15864_));
AND_g _21999_ (.A(_15863_), .B(_15864_), .Y(_15865_));
NAND_g _22000_ (.A(_11220_), .B(_15865_), .Y(_15866_));
NAND_g _22001_ (.A(_15844_), .B(_15866_), .Y(_15867_));
NAND_g _22002_ (.A(_11221_), .B(_15867_), .Y(_15868_));
NAND_g _22003_ (.A(_15822_), .B(_15868_), .Y(_15869_));
AND_g _22004_ (.A(_13734_), .B(_15869_), .Y(_15870_));
NAND_g _22005_ (.A(_14358_), .B(_15870_), .Y(_15871_));
AND_g _22006_ (.A(decoded_imm[20]), .B(_13830_), .Y(_15872_));
NAND_g _22007_ (.A(_13409_), .B(_15872_), .Y(_15873_));
AND_g _22008_ (.A(_13727_), .B(_15873_), .Y(_15874_));
NAND_g _22009_ (.A(_15871_), .B(_15874_), .Y(_15875_));
AND_g _22010_ (.A(_15776_), .B(_15875_), .Y(_00523_));
NAND_g _22011_ (.A(_11001_), .B(_13728_), .Y(_15876_));
NOR_g _22012_ (.A(cpuregs_16[21]), .B(_00011_[2]), .Y(_15877_));
AND_g _22013_ (.A(_11200_), .B(_00011_[2]), .Y(_15878_));
NOR_g _22014_ (.A(_15877_), .B(_15878_), .Y(_15879_));
NOR_g _22015_ (.A(cpuregs_18[21]), .B(_00011_[2]), .Y(_15880_));
AND_g _22016_ (.A(_11019_), .B(_00011_[2]), .Y(_15881_));
NOR_g _22017_ (.A(_15880_), .B(_15881_), .Y(_15882_));
NOR_g _22018_ (.A(cpuregs_17[21]), .B(_00011_[2]), .Y(_15883_));
NAND_g _22019_ (.A(_11033_), .B(_00011_[2]), .Y(_15884_));
NAND_g _22020_ (.A(_11186_), .B(_00011_[2]), .Y(_15885_));
NOR_g _22021_ (.A(cpuregs_19[21]), .B(_00011_[2]), .Y(_15886_));
NOR_g _22022_ (.A(_11217_), .B(_15886_), .Y(_15887_));
NAND_g _22023_ (.A(_15885_), .B(_15887_), .Y(_15888_));
NAND_g _22024_ (.A(_11217_), .B(_15882_), .Y(_15889_));
AND_g _22025_ (.A(_15888_), .B(_15889_), .Y(_15890_));
NAND_g _22026_ (.A(_00011_[1]), .B(_15890_), .Y(_15891_));
NOR_g _22027_ (.A(_11217_), .B(_15883_), .Y(_15892_));
NAND_g _22028_ (.A(_15884_), .B(_15892_), .Y(_15893_));
NAND_g _22029_ (.A(_11217_), .B(_15879_), .Y(_15894_));
AND_g _22030_ (.A(_15893_), .B(_15894_), .Y(_15895_));
NAND_g _22031_ (.A(_11218_), .B(_15895_), .Y(_15896_));
AND_g _22032_ (.A(_15891_), .B(_15896_), .Y(_15897_));
NAND_g _22033_ (.A(_11220_), .B(_15897_), .Y(_15898_));
NAND_g _22034_ (.A(cpuregs_27[21]), .B(_00011_[1]), .Y(_15899_));
NAND_g _22035_ (.A(cpuregs_25[21]), .B(_11218_), .Y(_15900_));
NAND_g _22036_ (.A(_15899_), .B(_15900_), .Y(_15901_));
NAND_g _22037_ (.A(_11219_), .B(_15901_), .Y(_15902_));
NAND_g _22038_ (.A(cpuregs_31[21]), .B(_00011_[1]), .Y(_15903_));
NAND_g _22039_ (.A(cpuregs_29[21]), .B(_11218_), .Y(_15904_));
NAND_g _22040_ (.A(_15903_), .B(_15904_), .Y(_15905_));
NAND_g _22041_ (.A(_00011_[2]), .B(_15905_), .Y(_15906_));
AND_g _22042_ (.A(_00011_[0]), .B(_15906_), .Y(_15907_));
NAND_g _22043_ (.A(_15902_), .B(_15907_), .Y(_15908_));
NAND_g _22044_ (.A(cpuregs_26[21]), .B(_00011_[1]), .Y(_15909_));
NAND_g _22045_ (.A(cpuregs_24[21]), .B(_11218_), .Y(_15910_));
NAND_g _22046_ (.A(_15909_), .B(_15910_), .Y(_15911_));
NAND_g _22047_ (.A(_11219_), .B(_15911_), .Y(_15912_));
NAND_g _22048_ (.A(cpuregs_30[21]), .B(_00011_[1]), .Y(_15913_));
NAND_g _22049_ (.A(cpuregs_28[21]), .B(_11218_), .Y(_15914_));
NAND_g _22050_ (.A(_15913_), .B(_15914_), .Y(_15915_));
NAND_g _22051_ (.A(_00011_[2]), .B(_15915_), .Y(_15916_));
AND_g _22052_ (.A(_11217_), .B(_15916_), .Y(_15917_));
NAND_g _22053_ (.A(_15912_), .B(_15917_), .Y(_15918_));
AND_g _22054_ (.A(_00011_[3]), .B(_15918_), .Y(_15919_));
NAND_g _22055_ (.A(_15908_), .B(_15919_), .Y(_15920_));
AND_g _22056_ (.A(_15898_), .B(_15920_), .Y(_15921_));
NAND_g _22057_ (.A(cpuregs_1[21]), .B(_11219_), .Y(_15922_));
NAND_g _22058_ (.A(cpuregs_5[21]), .B(_00011_[2]), .Y(_15923_));
AND_g _22059_ (.A(_00011_[0]), .B(_15923_), .Y(_15924_));
NAND_g _22060_ (.A(_15922_), .B(_15924_), .Y(_15925_));
NAND_g _22061_ (.A(cpuregs_0[21]), .B(_11219_), .Y(_15926_));
NAND_g _22062_ (.A(cpuregs_4[21]), .B(_00011_[2]), .Y(_15927_));
AND_g _22063_ (.A(_11217_), .B(_15927_), .Y(_15928_));
NAND_g _22064_ (.A(_15926_), .B(_15928_), .Y(_15929_));
AND_g _22065_ (.A(_11218_), .B(_15929_), .Y(_15930_));
NAND_g _22066_ (.A(_15925_), .B(_15930_), .Y(_15931_));
NAND_g _22067_ (.A(cpuregs_3[21]), .B(_11219_), .Y(_15932_));
NAND_g _22068_ (.A(cpuregs_7[21]), .B(_00011_[2]), .Y(_15933_));
AND_g _22069_ (.A(_00011_[0]), .B(_15933_), .Y(_15934_));
NAND_g _22070_ (.A(_15932_), .B(_15934_), .Y(_15935_));
NAND_g _22071_ (.A(cpuregs_2[21]), .B(_11219_), .Y(_15936_));
NAND_g _22072_ (.A(cpuregs_6[21]), .B(_00011_[2]), .Y(_15937_));
AND_g _22073_ (.A(_11217_), .B(_15937_), .Y(_15938_));
NAND_g _22074_ (.A(_15936_), .B(_15938_), .Y(_15939_));
AND_g _22075_ (.A(_00011_[1]), .B(_15939_), .Y(_15940_));
NAND_g _22076_ (.A(_15935_), .B(_15940_), .Y(_15941_));
NAND_g _22077_ (.A(_15931_), .B(_15941_), .Y(_15942_));
NAND_g _22078_ (.A(_11220_), .B(_15942_), .Y(_15943_));
NAND_g _22079_ (.A(cpuregs_14[21]), .B(_11217_), .Y(_15944_));
NAND_g _22080_ (.A(cpuregs_15[21]), .B(_00011_[0]), .Y(_15945_));
NAND_g _22081_ (.A(_15944_), .B(_15945_), .Y(_15946_));
NAND_g _22082_ (.A(_00011_[2]), .B(_15946_), .Y(_15947_));
NAND_g _22083_ (.A(cpuregs_10[21]), .B(_11217_), .Y(_15948_));
NAND_g _22084_ (.A(cpuregs_11[21]), .B(_00011_[0]), .Y(_15949_));
NAND_g _22085_ (.A(_15948_), .B(_15949_), .Y(_15950_));
NAND_g _22086_ (.A(_11219_), .B(_15950_), .Y(_15951_));
AND_g _22087_ (.A(_15947_), .B(_15951_), .Y(_15952_));
NAND_g _22088_ (.A(cpuregs_12[21]), .B(_11217_), .Y(_15953_));
NAND_g _22089_ (.A(cpuregs_13[21]), .B(_00011_[0]), .Y(_15954_));
NAND_g _22090_ (.A(_15953_), .B(_15954_), .Y(_15955_));
NAND_g _22091_ (.A(_00011_[2]), .B(_15955_), .Y(_15956_));
NAND_g _22092_ (.A(cpuregs_8[21]), .B(_11217_), .Y(_15957_));
NAND_g _22093_ (.A(cpuregs_9[21]), .B(_00011_[0]), .Y(_15958_));
NAND_g _22094_ (.A(_15957_), .B(_15958_), .Y(_15959_));
NAND_g _22095_ (.A(_11219_), .B(_15959_), .Y(_15960_));
AND_g _22096_ (.A(_15956_), .B(_15960_), .Y(_15961_));
NAND_g _22097_ (.A(_11218_), .B(_15961_), .Y(_15962_));
NAND_g _22098_ (.A(_00011_[1]), .B(_15952_), .Y(_15963_));
AND_g _22099_ (.A(_00011_[3]), .B(_15962_), .Y(_15964_));
NAND_g _22100_ (.A(_15963_), .B(_15964_), .Y(_15965_));
NAND_g _22101_ (.A(_00011_[4]), .B(_15921_), .Y(_15966_));
AND_g _22102_ (.A(_11221_), .B(_15943_), .Y(_15967_));
NAND_g _22103_ (.A(_15965_), .B(_15967_), .Y(_15968_));
AND_g _22104_ (.A(_13734_), .B(_15968_), .Y(_15969_));
AND_g _22105_ (.A(_15966_), .B(_15969_), .Y(_15970_));
NAND_g _22106_ (.A(_14358_), .B(_15970_), .Y(_15971_));
AND_g _22107_ (.A(decoded_imm[21]), .B(_13830_), .Y(_15972_));
NAND_g _22108_ (.A(_13409_), .B(_15972_), .Y(_15973_));
AND_g _22109_ (.A(_13727_), .B(_15973_), .Y(_15974_));
NAND_g _22110_ (.A(_15971_), .B(_15974_), .Y(_15975_));
AND_g _22111_ (.A(_15876_), .B(_15975_), .Y(_00524_));
NAND_g _22112_ (.A(_11002_), .B(_13728_), .Y(_15976_));
NAND_g _22113_ (.A(cpuregs_31[22]), .B(_00011_[1]), .Y(_15977_));
NAND_g _22114_ (.A(cpuregs_29[22]), .B(_11218_), .Y(_15978_));
NAND_g _22115_ (.A(_15977_), .B(_15978_), .Y(_15979_));
NAND_g _22116_ (.A(_00011_[2]), .B(_15979_), .Y(_15980_));
NAND_g _22117_ (.A(cpuregs_27[22]), .B(_00011_[1]), .Y(_15981_));
NAND_g _22118_ (.A(cpuregs_25[22]), .B(_11218_), .Y(_15982_));
NAND_g _22119_ (.A(_15981_), .B(_15982_), .Y(_15983_));
NAND_g _22120_ (.A(_11219_), .B(_15983_), .Y(_15984_));
NAND_g _22121_ (.A(_15980_), .B(_15984_), .Y(_15985_));
NAND_g _22122_ (.A(_00011_[0]), .B(_15985_), .Y(_15986_));
NAND_g _22123_ (.A(cpuregs_30[22]), .B(_00011_[1]), .Y(_15987_));
NAND_g _22124_ (.A(cpuregs_28[22]), .B(_11218_), .Y(_15988_));
NAND_g _22125_ (.A(_15987_), .B(_15988_), .Y(_15989_));
NAND_g _22126_ (.A(_00011_[2]), .B(_15989_), .Y(_15990_));
NAND_g _22127_ (.A(cpuregs_26[22]), .B(_00011_[1]), .Y(_15991_));
NAND_g _22128_ (.A(cpuregs_24[22]), .B(_11218_), .Y(_15992_));
NAND_g _22129_ (.A(_15991_), .B(_15992_), .Y(_15993_));
NAND_g _22130_ (.A(_11219_), .B(_15993_), .Y(_15994_));
NAND_g _22131_ (.A(_15990_), .B(_15994_), .Y(_15995_));
AND_g _22132_ (.A(_11217_), .B(_15995_), .Y(_15996_));
NOT_g _22133_ (.A(_15996_), .Y(_15997_));
NAND_g _22134_ (.A(_15986_), .B(_15997_), .Y(_15998_));
NAND_g _22135_ (.A(_00011_[3]), .B(_15998_), .Y(_15999_));
NOR_g _22136_ (.A(cpuregs_18[22]), .B(_00011_[2]), .Y(_16000_));
NOR_g _22137_ (.A(cpuregs_22[22]), .B(_11219_), .Y(_16001_));
NOR_g _22138_ (.A(_16000_), .B(_16001_), .Y(_16002_));
NOR_g _22139_ (.A(cpuregs_16[22]), .B(_00011_[2]), .Y(_16003_));
NOR_g _22140_ (.A(cpuregs_20[22]), .B(_11219_), .Y(_16004_));
NOR_g _22141_ (.A(_16003_), .B(_16004_), .Y(_16005_));
NAND_g _22142_ (.A(_11187_), .B(_00011_[2]), .Y(_16006_));
NOR_g _22143_ (.A(cpuregs_19[22]), .B(_00011_[2]), .Y(_16007_));
NOR_g _22144_ (.A(cpuregs_17[22]), .B(_00011_[2]), .Y(_16008_));
NAND_g _22145_ (.A(_11034_), .B(_00011_[2]), .Y(_16009_));
NOR_g _22146_ (.A(_11217_), .B(_16007_), .Y(_16010_));
NAND_g _22147_ (.A(_16006_), .B(_16010_), .Y(_16011_));
NAND_g _22148_ (.A(_11217_), .B(_16002_), .Y(_16012_));
AND_g _22149_ (.A(_16011_), .B(_16012_), .Y(_16013_));
NAND_g _22150_ (.A(_00011_[1]), .B(_16013_), .Y(_16014_));
NOR_g _22151_ (.A(_11217_), .B(_16008_), .Y(_16015_));
NAND_g _22152_ (.A(_16009_), .B(_16015_), .Y(_16016_));
NAND_g _22153_ (.A(_11217_), .B(_16005_), .Y(_16017_));
AND_g _22154_ (.A(_16016_), .B(_16017_), .Y(_16018_));
NAND_g _22155_ (.A(_11218_), .B(_16018_), .Y(_16019_));
AND_g _22156_ (.A(_16014_), .B(_16019_), .Y(_16020_));
NAND_g _22157_ (.A(_11220_), .B(_16020_), .Y(_16021_));
NAND_g _22158_ (.A(_15999_), .B(_16021_), .Y(_16022_));
NAND_g _22159_ (.A(_00011_[4]), .B(_16022_), .Y(_16023_));
NAND_g _22160_ (.A(cpuregs_13[22]), .B(_11218_), .Y(_16024_));
NAND_g _22161_ (.A(cpuregs_15[22]), .B(_00011_[1]), .Y(_16025_));
AND_g _22162_ (.A(_00011_[2]), .B(_16025_), .Y(_16026_));
NAND_g _22163_ (.A(_16024_), .B(_16026_), .Y(_16027_));
NAND_g _22164_ (.A(cpuregs_9[22]), .B(_11218_), .Y(_16028_));
NAND_g _22165_ (.A(cpuregs_11[22]), .B(_00011_[1]), .Y(_16029_));
AND_g _22166_ (.A(_11219_), .B(_16029_), .Y(_16030_));
NAND_g _22167_ (.A(_16028_), .B(_16030_), .Y(_16031_));
AND_g _22168_ (.A(_00011_[0]), .B(_16031_), .Y(_16032_));
NAND_g _22169_ (.A(_16027_), .B(_16032_), .Y(_16033_));
NAND_g _22170_ (.A(cpuregs_12[22]), .B(_11218_), .Y(_16034_));
NAND_g _22171_ (.A(cpuregs_14[22]), .B(_00011_[1]), .Y(_16035_));
AND_g _22172_ (.A(_00011_[2]), .B(_16035_), .Y(_16036_));
NAND_g _22173_ (.A(_16034_), .B(_16036_), .Y(_16037_));
NAND_g _22174_ (.A(cpuregs_8[22]), .B(_11218_), .Y(_16038_));
NAND_g _22175_ (.A(cpuregs_10[22]), .B(_00011_[1]), .Y(_16039_));
AND_g _22176_ (.A(_11219_), .B(_16039_), .Y(_16040_));
NAND_g _22177_ (.A(_16038_), .B(_16040_), .Y(_16041_));
AND_g _22178_ (.A(_11217_), .B(_16041_), .Y(_16042_));
NAND_g _22179_ (.A(_16037_), .B(_16042_), .Y(_16043_));
NAND_g _22180_ (.A(_16033_), .B(_16043_), .Y(_16044_));
NAND_g _22181_ (.A(_00011_[3]), .B(_16044_), .Y(_16045_));
NAND_g _22182_ (.A(_10946_), .B(_00011_[2]), .Y(_16046_));
NOR_g _22183_ (.A(cpuregs_2[22]), .B(_00011_[2]), .Y(_16047_));
NOR_g _22184_ (.A(_00011_[0]), .B(_16047_), .Y(_16048_));
NAND_g _22185_ (.A(_16046_), .B(_16048_), .Y(_16049_));
NAND_g _22186_ (.A(_11132_), .B(_00011_[2]), .Y(_16050_));
NOR_g _22187_ (.A(cpuregs_3[22]), .B(_00011_[2]), .Y(_16051_));
NOR_g _22188_ (.A(_11217_), .B(_16051_), .Y(_16052_));
NAND_g _22189_ (.A(_16050_), .B(_16052_), .Y(_16053_));
AND_g _22190_ (.A(_16049_), .B(_16053_), .Y(_16054_));
NAND_g _22191_ (.A(_10958_), .B(_00011_[2]), .Y(_16055_));
NOR_g _22192_ (.A(cpuregs_0[22]), .B(_00011_[2]), .Y(_16056_));
NOR_g _22193_ (.A(_00011_[0]), .B(_16056_), .Y(_16057_));
NAND_g _22194_ (.A(_16055_), .B(_16057_), .Y(_16058_));
NAND_g _22195_ (.A(_11116_), .B(_00011_[2]), .Y(_16059_));
NOR_g _22196_ (.A(cpuregs_1[22]), .B(_00011_[2]), .Y(_16060_));
NOR_g _22197_ (.A(_11217_), .B(_16060_), .Y(_16061_));
NAND_g _22198_ (.A(_16059_), .B(_16061_), .Y(_16062_));
AND_g _22199_ (.A(_16058_), .B(_16062_), .Y(_16063_));
NAND_g _22200_ (.A(_00011_[1]), .B(_16054_), .Y(_16064_));
NAND_g _22201_ (.A(_11218_), .B(_16063_), .Y(_16065_));
AND_g _22202_ (.A(_16064_), .B(_16065_), .Y(_16066_));
NAND_g _22203_ (.A(_11220_), .B(_16066_), .Y(_16067_));
NAND_g _22204_ (.A(_16045_), .B(_16067_), .Y(_16068_));
NAND_g _22205_ (.A(_11221_), .B(_16068_), .Y(_16069_));
NAND_g _22206_ (.A(_16023_), .B(_16069_), .Y(_16070_));
AND_g _22207_ (.A(_13734_), .B(_16070_), .Y(_16071_));
NAND_g _22208_ (.A(_13833_), .B(_16071_), .Y(_16072_));
NAND_g _22209_ (.A(decoded_imm[22]), .B(_13830_), .Y(_16073_));
NAND_g _22210_ (.A(_16072_), .B(_16073_), .Y(_16074_));
NAND_g _22211_ (.A(_13409_), .B(_16074_), .Y(_16075_));
AND_g _22212_ (.A(_13724_), .B(_16071_), .Y(_16076_));
NOR_g _22213_ (.A(_13728_), .B(_16076_), .Y(_16077_));
NAND_g _22214_ (.A(_16075_), .B(_16077_), .Y(_16078_));
AND_g _22215_ (.A(_15976_), .B(_16078_), .Y(_00525_));
NAND_g _22216_ (.A(_11003_), .B(_13728_), .Y(_16079_));
NAND_g _22217_ (.A(cpuregs_24[23]), .B(_11219_), .Y(_16080_));
NAND_g _22218_ (.A(cpuregs_28[23]), .B(_00011_[2]), .Y(_16081_));
AND_g _22219_ (.A(_11217_), .B(_16081_), .Y(_16082_));
NAND_g _22220_ (.A(_16080_), .B(_16082_), .Y(_16083_));
NAND_g _22221_ (.A(cpuregs_25[23]), .B(_11219_), .Y(_16084_));
NAND_g _22222_ (.A(cpuregs_29[23]), .B(_00011_[2]), .Y(_16085_));
AND_g _22223_ (.A(_00011_[0]), .B(_16085_), .Y(_16086_));
NAND_g _22224_ (.A(_16084_), .B(_16086_), .Y(_16087_));
NAND_g _22225_ (.A(_16083_), .B(_16087_), .Y(_16088_));
NAND_g _22226_ (.A(_11218_), .B(_16088_), .Y(_16089_));
NAND_g _22227_ (.A(cpuregs_26[23]), .B(_11219_), .Y(_16090_));
NAND_g _22228_ (.A(cpuregs_30[23]), .B(_00011_[2]), .Y(_16091_));
AND_g _22229_ (.A(_11217_), .B(_16091_), .Y(_16092_));
NAND_g _22230_ (.A(_16090_), .B(_16092_), .Y(_16093_));
NAND_g _22231_ (.A(cpuregs_31[23]), .B(_00011_[2]), .Y(_16094_));
NAND_g _22232_ (.A(cpuregs_27[23]), .B(_11219_), .Y(_16095_));
AND_g _22233_ (.A(_00011_[0]), .B(_16095_), .Y(_16096_));
NAND_g _22234_ (.A(_16094_), .B(_16096_), .Y(_16097_));
NAND_g _22235_ (.A(_16093_), .B(_16097_), .Y(_16098_));
NAND_g _22236_ (.A(_00011_[1]), .B(_16098_), .Y(_16099_));
AND_g _22237_ (.A(_00011_[3]), .B(_16089_), .Y(_16100_));
NAND_g _22238_ (.A(_16099_), .B(_16100_), .Y(_16101_));
NAND_g _22239_ (.A(cpuregs_20[23]), .B(_00011_[2]), .Y(_16102_));
NAND_g _22240_ (.A(cpuregs_16[23]), .B(_11219_), .Y(_16103_));
AND_g _22241_ (.A(_16102_), .B(_16103_), .Y(_16104_));
NAND_g _22242_ (.A(_11217_), .B(_16104_), .Y(_16105_));
NAND_g _22243_ (.A(cpuregs_21[23]), .B(_00011_[2]), .Y(_16106_));
NAND_g _22244_ (.A(cpuregs_17[23]), .B(_11219_), .Y(_16107_));
AND_g _22245_ (.A(_00011_[0]), .B(_16107_), .Y(_16108_));
NAND_g _22246_ (.A(_16106_), .B(_16108_), .Y(_16109_));
AND_g _22247_ (.A(_11218_), .B(_16109_), .Y(_16110_));
NAND_g _22248_ (.A(_16105_), .B(_16110_), .Y(_16111_));
NAND_g _22249_ (.A(cpuregs_23[23]), .B(_00011_[2]), .Y(_16112_));
NAND_g _22250_ (.A(cpuregs_19[23]), .B(_11219_), .Y(_16113_));
AND_g _22251_ (.A(_00011_[0]), .B(_16113_), .Y(_16114_));
NAND_g _22252_ (.A(_16112_), .B(_16114_), .Y(_16115_));
NAND_g _22253_ (.A(cpuregs_22[23]), .B(_00011_[2]), .Y(_16116_));
NAND_g _22254_ (.A(cpuregs_18[23]), .B(_11219_), .Y(_16117_));
AND_g _22255_ (.A(_16116_), .B(_16117_), .Y(_16118_));
NAND_g _22256_ (.A(_11217_), .B(_16118_), .Y(_16119_));
AND_g _22257_ (.A(_00011_[1]), .B(_16119_), .Y(_16120_));
NAND_g _22258_ (.A(_16115_), .B(_16120_), .Y(_16121_));
NAND_g _22259_ (.A(_16111_), .B(_16121_), .Y(_16122_));
NAND_g _22260_ (.A(_11220_), .B(_16122_), .Y(_16123_));
AND_g _22261_ (.A(_16101_), .B(_16123_), .Y(_16124_));
NAND_g _22262_ (.A(cpuregs_13[23]), .B(_11218_), .Y(_16125_));
NAND_g _22263_ (.A(cpuregs_15[23]), .B(_00011_[1]), .Y(_16126_));
AND_g _22264_ (.A(_00011_[2]), .B(_16126_), .Y(_16127_));
NAND_g _22265_ (.A(_16125_), .B(_16127_), .Y(_16128_));
NAND_g _22266_ (.A(cpuregs_9[23]), .B(_11218_), .Y(_16129_));
NAND_g _22267_ (.A(cpuregs_11[23]), .B(_00011_[1]), .Y(_16130_));
AND_g _22268_ (.A(_11219_), .B(_16130_), .Y(_16131_));
NAND_g _22269_ (.A(_16129_), .B(_16131_), .Y(_16132_));
AND_g _22270_ (.A(_00011_[0]), .B(_16132_), .Y(_16133_));
NAND_g _22271_ (.A(_16128_), .B(_16133_), .Y(_16134_));
NAND_g _22272_ (.A(cpuregs_12[23]), .B(_11218_), .Y(_16135_));
NAND_g _22273_ (.A(cpuregs_14[23]), .B(_00011_[1]), .Y(_16136_));
AND_g _22274_ (.A(_00011_[2]), .B(_16136_), .Y(_16137_));
NAND_g _22275_ (.A(_16135_), .B(_16137_), .Y(_16138_));
NAND_g _22276_ (.A(cpuregs_8[23]), .B(_11218_), .Y(_16139_));
NAND_g _22277_ (.A(cpuregs_10[23]), .B(_00011_[1]), .Y(_16140_));
AND_g _22278_ (.A(_11219_), .B(_16140_), .Y(_16141_));
NAND_g _22279_ (.A(_16139_), .B(_16141_), .Y(_16142_));
AND_g _22280_ (.A(_11217_), .B(_16142_), .Y(_16143_));
NAND_g _22281_ (.A(_16138_), .B(_16143_), .Y(_16144_));
NAND_g _22282_ (.A(_16134_), .B(_16144_), .Y(_16145_));
NAND_g _22283_ (.A(_00011_[3]), .B(_16145_), .Y(_16146_));
NAND_g _22284_ (.A(_10947_), .B(_00011_[2]), .Y(_16147_));
NOR_g _22285_ (.A(cpuregs_2[23]), .B(_00011_[2]), .Y(_16148_));
NOR_g _22286_ (.A(_00011_[0]), .B(_16148_), .Y(_16149_));
NAND_g _22287_ (.A(_16147_), .B(_16149_), .Y(_16150_));
NAND_g _22288_ (.A(_11133_), .B(_00011_[2]), .Y(_16151_));
NOR_g _22289_ (.A(cpuregs_3[23]), .B(_00011_[2]), .Y(_16152_));
NOR_g _22290_ (.A(_11217_), .B(_16152_), .Y(_16153_));
NAND_g _22291_ (.A(_16151_), .B(_16153_), .Y(_16154_));
AND_g _22292_ (.A(_16150_), .B(_16154_), .Y(_16155_));
NAND_g _22293_ (.A(_10959_), .B(_00011_[2]), .Y(_16156_));
NOR_g _22294_ (.A(cpuregs_0[23]), .B(_00011_[2]), .Y(_16157_));
NOR_g _22295_ (.A(_00011_[0]), .B(_16157_), .Y(_16158_));
NAND_g _22296_ (.A(_16156_), .B(_16158_), .Y(_16159_));
NAND_g _22297_ (.A(_11117_), .B(_00011_[2]), .Y(_16160_));
NOR_g _22298_ (.A(cpuregs_1[23]), .B(_00011_[2]), .Y(_16161_));
NOR_g _22299_ (.A(_11217_), .B(_16161_), .Y(_16162_));
NAND_g _22300_ (.A(_16160_), .B(_16162_), .Y(_16163_));
NAND_g _22301_ (.A(_00011_[1]), .B(_16155_), .Y(_16164_));
AND_g _22302_ (.A(_11218_), .B(_16159_), .Y(_16165_));
NAND_g _22303_ (.A(_16163_), .B(_16165_), .Y(_16166_));
AND_g _22304_ (.A(_16164_), .B(_16166_), .Y(_16167_));
NAND_g _22305_ (.A(_11220_), .B(_16167_), .Y(_16168_));
NAND_g _22306_ (.A(_16146_), .B(_16168_), .Y(_16169_));
NAND_g _22307_ (.A(_00011_[4]), .B(_16124_), .Y(_16170_));
NOR_g _22308_ (.A(_00011_[4]), .B(_16169_), .Y(_16171_));
NOR_g _22309_ (.A(_13733_), .B(_16171_), .Y(_16172_));
AND_g _22310_ (.A(_16170_), .B(_16172_), .Y(_16173_));
NAND_g _22311_ (.A(_14358_), .B(_16173_), .Y(_16174_));
AND_g _22312_ (.A(decoded_imm[23]), .B(_13830_), .Y(_16175_));
NAND_g _22313_ (.A(_13409_), .B(_16175_), .Y(_16176_));
AND_g _22314_ (.A(_13727_), .B(_16176_), .Y(_16177_));
NAND_g _22315_ (.A(_16174_), .B(_16177_), .Y(_16178_));
AND_g _22316_ (.A(_16079_), .B(_16178_), .Y(_00526_));
NAND_g _22317_ (.A(_11004_), .B(_13728_), .Y(_16179_));
NAND_g _22318_ (.A(cpuregs_29[24]), .B(_00011_[2]), .Y(_16180_));
NAND_g _22319_ (.A(cpuregs_25[24]), .B(_11219_), .Y(_16181_));
AND_g _22320_ (.A(_00011_[0]), .B(_16181_), .Y(_16182_));
NAND_g _22321_ (.A(_16180_), .B(_16182_), .Y(_16183_));
NAND_g _22322_ (.A(cpuregs_24[24]), .B(_11219_), .Y(_16184_));
NAND_g _22323_ (.A(cpuregs_28[24]), .B(_00011_[2]), .Y(_16185_));
AND_g _22324_ (.A(_11217_), .B(_16185_), .Y(_16186_));
NAND_g _22325_ (.A(_16184_), .B(_16186_), .Y(_16187_));
AND_g _22326_ (.A(_11218_), .B(_16187_), .Y(_16188_));
NAND_g _22327_ (.A(_16183_), .B(_16188_), .Y(_16189_));
NAND_g _22328_ (.A(cpuregs_27[24]), .B(_11219_), .Y(_16190_));
NAND_g _22329_ (.A(cpuregs_31[24]), .B(_00011_[2]), .Y(_16191_));
AND_g _22330_ (.A(_00011_[0]), .B(_16191_), .Y(_16192_));
NAND_g _22331_ (.A(_16190_), .B(_16192_), .Y(_16193_));
NAND_g _22332_ (.A(cpuregs_26[24]), .B(_11219_), .Y(_16194_));
NAND_g _22333_ (.A(cpuregs_30[24]), .B(_00011_[2]), .Y(_16195_));
AND_g _22334_ (.A(_11217_), .B(_16195_), .Y(_16196_));
NAND_g _22335_ (.A(_16194_), .B(_16196_), .Y(_16197_));
AND_g _22336_ (.A(_00011_[1]), .B(_16197_), .Y(_16198_));
NAND_g _22337_ (.A(_16193_), .B(_16198_), .Y(_16199_));
NAND_g _22338_ (.A(_16189_), .B(_16199_), .Y(_16200_));
NAND_g _22339_ (.A(_00011_[4]), .B(_16200_), .Y(_16201_));
NAND_g _22340_ (.A(cpuregs_14[24]), .B(_11217_), .Y(_16202_));
NAND_g _22341_ (.A(cpuregs_15[24]), .B(_00011_[0]), .Y(_16203_));
NAND_g _22342_ (.A(_16202_), .B(_16203_), .Y(_16204_));
NAND_g _22343_ (.A(_00011_[2]), .B(_16204_), .Y(_16205_));
NAND_g _22344_ (.A(cpuregs_10[24]), .B(_11217_), .Y(_16206_));
NAND_g _22345_ (.A(cpuregs_11[24]), .B(_00011_[0]), .Y(_16207_));
NAND_g _22346_ (.A(_16206_), .B(_16207_), .Y(_16208_));
NAND_g _22347_ (.A(_11219_), .B(_16208_), .Y(_16209_));
NAND_g _22348_ (.A(_16205_), .B(_16209_), .Y(_16210_));
NAND_g _22349_ (.A(_00011_[1]), .B(_16210_), .Y(_16211_));
NAND_g _22350_ (.A(cpuregs_12[24]), .B(_11217_), .Y(_16212_));
NAND_g _22351_ (.A(cpuregs_13[24]), .B(_00011_[0]), .Y(_16213_));
NAND_g _22352_ (.A(_16212_), .B(_16213_), .Y(_16214_));
NAND_g _22353_ (.A(_00011_[2]), .B(_16214_), .Y(_16215_));
NAND_g _22354_ (.A(cpuregs_8[24]), .B(_11217_), .Y(_16216_));
NAND_g _22355_ (.A(cpuregs_9[24]), .B(_00011_[0]), .Y(_16217_));
NAND_g _22356_ (.A(_16216_), .B(_16217_), .Y(_16218_));
NAND_g _22357_ (.A(_11219_), .B(_16218_), .Y(_16219_));
NAND_g _22358_ (.A(_16215_), .B(_16219_), .Y(_16220_));
NAND_g _22359_ (.A(_11218_), .B(_16220_), .Y(_16221_));
NAND_g _22360_ (.A(_16211_), .B(_16221_), .Y(_16222_));
NAND_g _22361_ (.A(_11221_), .B(_16222_), .Y(_16223_));
NAND_g _22362_ (.A(_16201_), .B(_16223_), .Y(_16224_));
NAND_g _22363_ (.A(_00011_[3]), .B(_16224_), .Y(_16225_));
NAND_g _22364_ (.A(cpuregs_1[24]), .B(_11219_), .Y(_16226_));
NAND_g _22365_ (.A(cpuregs_5[24]), .B(_00011_[2]), .Y(_16227_));
AND_g _22366_ (.A(_00011_[0]), .B(_16227_), .Y(_16228_));
NAND_g _22367_ (.A(_16226_), .B(_16228_), .Y(_16229_));
NAND_g _22368_ (.A(cpuregs_0[24]), .B(_11219_), .Y(_16230_));
NAND_g _22369_ (.A(cpuregs_4[24]), .B(_00011_[2]), .Y(_16231_));
AND_g _22370_ (.A(_11217_), .B(_16231_), .Y(_16232_));
NAND_g _22371_ (.A(_16230_), .B(_16232_), .Y(_16233_));
AND_g _22372_ (.A(_11218_), .B(_16233_), .Y(_16234_));
NAND_g _22373_ (.A(_16229_), .B(_16234_), .Y(_16235_));
NAND_g _22374_ (.A(cpuregs_3[24]), .B(_11219_), .Y(_16236_));
NAND_g _22375_ (.A(cpuregs_7[24]), .B(_00011_[2]), .Y(_16237_));
AND_g _22376_ (.A(_00011_[0]), .B(_16237_), .Y(_16238_));
NAND_g _22377_ (.A(_16236_), .B(_16238_), .Y(_16239_));
NAND_g _22378_ (.A(cpuregs_2[24]), .B(_11219_), .Y(_16240_));
NAND_g _22379_ (.A(cpuregs_6[24]), .B(_00011_[2]), .Y(_16241_));
AND_g _22380_ (.A(_11217_), .B(_16241_), .Y(_16242_));
NAND_g _22381_ (.A(_16240_), .B(_16242_), .Y(_16243_));
AND_g _22382_ (.A(_00011_[1]), .B(_16243_), .Y(_16244_));
NAND_g _22383_ (.A(_16239_), .B(_16244_), .Y(_16245_));
NAND_g _22384_ (.A(_16235_), .B(_16245_), .Y(_16246_));
NAND_g _22385_ (.A(_11221_), .B(_16246_), .Y(_16247_));
NAND_g _22386_ (.A(cpuregs_19[24]), .B(_00011_[1]), .Y(_16248_));
NAND_g _22387_ (.A(cpuregs_17[24]), .B(_11218_), .Y(_16249_));
NAND_g _22388_ (.A(_16248_), .B(_16249_), .Y(_16250_));
NAND_g _22389_ (.A(_11219_), .B(_16250_), .Y(_16251_));
NAND_g _22390_ (.A(cpuregs_23[24]), .B(_00011_[1]), .Y(_16252_));
NAND_g _22391_ (.A(cpuregs_21[24]), .B(_11218_), .Y(_16253_));
NAND_g _22392_ (.A(_16252_), .B(_16253_), .Y(_16254_));
NAND_g _22393_ (.A(_00011_[2]), .B(_16254_), .Y(_16255_));
AND_g _22394_ (.A(_00011_[0]), .B(_16255_), .Y(_16256_));
NAND_g _22395_ (.A(_16251_), .B(_16256_), .Y(_16257_));
NAND_g _22396_ (.A(cpuregs_18[24]), .B(_00011_[1]), .Y(_16258_));
NAND_g _22397_ (.A(cpuregs_16[24]), .B(_11218_), .Y(_16259_));
NAND_g _22398_ (.A(_16258_), .B(_16259_), .Y(_16260_));
NAND_g _22399_ (.A(_11219_), .B(_16260_), .Y(_16261_));
NAND_g _22400_ (.A(cpuregs_22[24]), .B(_00011_[1]), .Y(_16262_));
NAND_g _22401_ (.A(cpuregs_20[24]), .B(_11218_), .Y(_16263_));
NAND_g _22402_ (.A(_16262_), .B(_16263_), .Y(_16264_));
NAND_g _22403_ (.A(_00011_[2]), .B(_16264_), .Y(_16265_));
AND_g _22404_ (.A(_11217_), .B(_16265_), .Y(_16266_));
NAND_g _22405_ (.A(_16261_), .B(_16266_), .Y(_16267_));
AND_g _22406_ (.A(_00011_[4]), .B(_16267_), .Y(_16268_));
NAND_g _22407_ (.A(_16257_), .B(_16268_), .Y(_16269_));
NAND_g _22408_ (.A(_16247_), .B(_16269_), .Y(_16270_));
NAND_g _22409_ (.A(_11220_), .B(_16270_), .Y(_16271_));
NAND_g _22410_ (.A(_16225_), .B(_16271_), .Y(_16272_));
AND_g _22411_ (.A(_13734_), .B(_16272_), .Y(_16273_));
NAND_g _22412_ (.A(_14358_), .B(_16273_), .Y(_16274_));
AND_g _22413_ (.A(decoded_imm[24]), .B(_13830_), .Y(_16275_));
NAND_g _22414_ (.A(_13409_), .B(_16275_), .Y(_16276_));
AND_g _22415_ (.A(_13727_), .B(_16276_), .Y(_16277_));
NAND_g _22416_ (.A(_16274_), .B(_16277_), .Y(_16278_));
AND_g _22417_ (.A(_16179_), .B(_16278_), .Y(_00527_));
NAND_g _22418_ (.A(_11005_), .B(_13728_), .Y(_16279_));
NOR_g _22419_ (.A(cpuregs_16[25]), .B(_00011_[2]), .Y(_16280_));
NOR_g _22420_ (.A(cpuregs_20[25]), .B(_11219_), .Y(_16281_));
NOR_g _22421_ (.A(_16280_), .B(_16281_), .Y(_16282_));
NOR_g _22422_ (.A(cpuregs_18[25]), .B(_00011_[2]), .Y(_16283_));
NOR_g _22423_ (.A(cpuregs_22[25]), .B(_11219_), .Y(_16284_));
NOR_g _22424_ (.A(_16283_), .B(_16284_), .Y(_16285_));
NOR_g _22425_ (.A(cpuregs_17[25]), .B(_00011_[2]), .Y(_16286_));
NAND_g _22426_ (.A(_11035_), .B(_00011_[2]), .Y(_16287_));
NAND_g _22427_ (.A(_11188_), .B(_00011_[2]), .Y(_16288_));
NOR_g _22428_ (.A(cpuregs_19[25]), .B(_00011_[2]), .Y(_16289_));
NOR_g _22429_ (.A(_11217_), .B(_16289_), .Y(_16290_));
NAND_g _22430_ (.A(_16288_), .B(_16290_), .Y(_16291_));
NAND_g _22431_ (.A(_11217_), .B(_16285_), .Y(_16292_));
AND_g _22432_ (.A(_16291_), .B(_16292_), .Y(_16293_));
NAND_g _22433_ (.A(_00011_[1]), .B(_16293_), .Y(_16294_));
NOR_g _22434_ (.A(_11217_), .B(_16286_), .Y(_16295_));
NAND_g _22435_ (.A(_16287_), .B(_16295_), .Y(_16296_));
NAND_g _22436_ (.A(_11217_), .B(_16282_), .Y(_16297_));
AND_g _22437_ (.A(_16296_), .B(_16297_), .Y(_16298_));
NAND_g _22438_ (.A(_11218_), .B(_16298_), .Y(_16299_));
AND_g _22439_ (.A(_16294_), .B(_16299_), .Y(_16300_));
NAND_g _22440_ (.A(_11220_), .B(_16300_), .Y(_16301_));
NAND_g _22441_ (.A(cpuregs_27[25]), .B(_00011_[1]), .Y(_16302_));
NAND_g _22442_ (.A(cpuregs_25[25]), .B(_11218_), .Y(_16303_));
NAND_g _22443_ (.A(_16302_), .B(_16303_), .Y(_16304_));
NAND_g _22444_ (.A(_11219_), .B(_16304_), .Y(_16305_));
NAND_g _22445_ (.A(cpuregs_31[25]), .B(_00011_[1]), .Y(_16306_));
NAND_g _22446_ (.A(cpuregs_29[25]), .B(_11218_), .Y(_16307_));
NAND_g _22447_ (.A(_16306_), .B(_16307_), .Y(_16308_));
NAND_g _22448_ (.A(_00011_[2]), .B(_16308_), .Y(_16309_));
AND_g _22449_ (.A(_00011_[0]), .B(_16309_), .Y(_16310_));
NAND_g _22450_ (.A(_16305_), .B(_16310_), .Y(_16311_));
NAND_g _22451_ (.A(cpuregs_26[25]), .B(_00011_[1]), .Y(_16312_));
NAND_g _22452_ (.A(cpuregs_24[25]), .B(_11218_), .Y(_16313_));
NAND_g _22453_ (.A(_16312_), .B(_16313_), .Y(_16314_));
NAND_g _22454_ (.A(_11219_), .B(_16314_), .Y(_16315_));
NAND_g _22455_ (.A(cpuregs_30[25]), .B(_00011_[1]), .Y(_16316_));
NAND_g _22456_ (.A(cpuregs_28[25]), .B(_11218_), .Y(_16317_));
NAND_g _22457_ (.A(_16316_), .B(_16317_), .Y(_16318_));
NAND_g _22458_ (.A(_00011_[2]), .B(_16318_), .Y(_16319_));
AND_g _22459_ (.A(_11217_), .B(_16319_), .Y(_16320_));
NAND_g _22460_ (.A(_16315_), .B(_16320_), .Y(_16321_));
AND_g _22461_ (.A(_00011_[3]), .B(_16321_), .Y(_16322_));
NAND_g _22462_ (.A(_16311_), .B(_16322_), .Y(_16323_));
AND_g _22463_ (.A(_16301_), .B(_16323_), .Y(_16324_));
NAND_g _22464_ (.A(cpuregs_1[25]), .B(_11219_), .Y(_16325_));
NAND_g _22465_ (.A(cpuregs_5[25]), .B(_00011_[2]), .Y(_16326_));
AND_g _22466_ (.A(_00011_[0]), .B(_16326_), .Y(_16327_));
NAND_g _22467_ (.A(_16325_), .B(_16327_), .Y(_16328_));
NAND_g _22468_ (.A(cpuregs_0[25]), .B(_11219_), .Y(_16329_));
NAND_g _22469_ (.A(cpuregs_4[25]), .B(_00011_[2]), .Y(_16330_));
AND_g _22470_ (.A(_11217_), .B(_16330_), .Y(_16331_));
NAND_g _22471_ (.A(_16329_), .B(_16331_), .Y(_16332_));
AND_g _22472_ (.A(_11218_), .B(_16332_), .Y(_16333_));
NAND_g _22473_ (.A(_16328_), .B(_16333_), .Y(_16334_));
NAND_g _22474_ (.A(cpuregs_3[25]), .B(_11219_), .Y(_16335_));
NAND_g _22475_ (.A(cpuregs_7[25]), .B(_00011_[2]), .Y(_16336_));
AND_g _22476_ (.A(_00011_[0]), .B(_16336_), .Y(_16337_));
NAND_g _22477_ (.A(_16335_), .B(_16337_), .Y(_16338_));
NAND_g _22478_ (.A(cpuregs_2[25]), .B(_11219_), .Y(_16339_));
NAND_g _22479_ (.A(cpuregs_6[25]), .B(_00011_[2]), .Y(_16340_));
AND_g _22480_ (.A(_11217_), .B(_16340_), .Y(_16341_));
NAND_g _22481_ (.A(_16339_), .B(_16341_), .Y(_16342_));
AND_g _22482_ (.A(_00011_[1]), .B(_16342_), .Y(_16343_));
NAND_g _22483_ (.A(_16338_), .B(_16343_), .Y(_16344_));
NAND_g _22484_ (.A(_16334_), .B(_16344_), .Y(_16345_));
NAND_g _22485_ (.A(_11220_), .B(_16345_), .Y(_16346_));
NAND_g _22486_ (.A(cpuregs_14[25]), .B(_11217_), .Y(_16347_));
NAND_g _22487_ (.A(cpuregs_15[25]), .B(_00011_[0]), .Y(_16348_));
NAND_g _22488_ (.A(_16347_), .B(_16348_), .Y(_16349_));
NAND_g _22489_ (.A(_00011_[2]), .B(_16349_), .Y(_16350_));
NAND_g _22490_ (.A(cpuregs_10[25]), .B(_11217_), .Y(_16351_));
NAND_g _22491_ (.A(cpuregs_11[25]), .B(_00011_[0]), .Y(_16352_));
NAND_g _22492_ (.A(_16351_), .B(_16352_), .Y(_16353_));
NAND_g _22493_ (.A(_11219_), .B(_16353_), .Y(_16354_));
AND_g _22494_ (.A(_16350_), .B(_16354_), .Y(_16355_));
NAND_g _22495_ (.A(cpuregs_12[25]), .B(_11217_), .Y(_16356_));
NAND_g _22496_ (.A(cpuregs_13[25]), .B(_00011_[0]), .Y(_16357_));
NAND_g _22497_ (.A(_16356_), .B(_16357_), .Y(_16358_));
NAND_g _22498_ (.A(_00011_[2]), .B(_16358_), .Y(_16359_));
NAND_g _22499_ (.A(cpuregs_8[25]), .B(_11217_), .Y(_16360_));
NAND_g _22500_ (.A(cpuregs_9[25]), .B(_00011_[0]), .Y(_16361_));
NAND_g _22501_ (.A(_16360_), .B(_16361_), .Y(_16362_));
NAND_g _22502_ (.A(_11219_), .B(_16362_), .Y(_16363_));
AND_g _22503_ (.A(_16359_), .B(_16363_), .Y(_16364_));
NAND_g _22504_ (.A(_11218_), .B(_16364_), .Y(_16365_));
NAND_g _22505_ (.A(_00011_[1]), .B(_16355_), .Y(_16366_));
AND_g _22506_ (.A(_00011_[3]), .B(_16365_), .Y(_16367_));
NAND_g _22507_ (.A(_16366_), .B(_16367_), .Y(_16368_));
NAND_g _22508_ (.A(_00011_[4]), .B(_16324_), .Y(_16369_));
AND_g _22509_ (.A(_11221_), .B(_16346_), .Y(_16370_));
NAND_g _22510_ (.A(_16368_), .B(_16370_), .Y(_16371_));
AND_g _22511_ (.A(_13734_), .B(_16371_), .Y(_16372_));
AND_g _22512_ (.A(_16369_), .B(_16372_), .Y(_16373_));
NAND_g _22513_ (.A(_13833_), .B(_16373_), .Y(_16374_));
NAND_g _22514_ (.A(decoded_imm[25]), .B(_13830_), .Y(_16375_));
NAND_g _22515_ (.A(_16374_), .B(_16375_), .Y(_16376_));
NAND_g _22516_ (.A(_13409_), .B(_16376_), .Y(_16377_));
AND_g _22517_ (.A(_13724_), .B(_16373_), .Y(_16378_));
NOR_g _22518_ (.A(_13728_), .B(_16378_), .Y(_16379_));
NAND_g _22519_ (.A(_16377_), .B(_16379_), .Y(_16380_));
AND_g _22520_ (.A(_16279_), .B(_16380_), .Y(_00528_));
NAND_g _22521_ (.A(_11006_), .B(_13728_), .Y(_16381_));
NOR_g _22522_ (.A(cpuregs_16[26]), .B(_00011_[2]), .Y(_16382_));
AND_g _22523_ (.A(_11201_), .B(_00011_[2]), .Y(_16383_));
NOR_g _22524_ (.A(_16382_), .B(_16383_), .Y(_16384_));
NOR_g _22525_ (.A(cpuregs_18[26]), .B(_00011_[2]), .Y(_16385_));
AND_g _22526_ (.A(_11020_), .B(_00011_[2]), .Y(_16386_));
NOR_g _22527_ (.A(_16385_), .B(_16386_), .Y(_16387_));
NOR_g _22528_ (.A(cpuregs_17[26]), .B(_00011_[2]), .Y(_16388_));
NAND_g _22529_ (.A(_11036_), .B(_00011_[2]), .Y(_16389_));
NAND_g _22530_ (.A(_11189_), .B(_00011_[2]), .Y(_16390_));
NOR_g _22531_ (.A(cpuregs_19[26]), .B(_00011_[2]), .Y(_16391_));
NOR_g _22532_ (.A(_11217_), .B(_16391_), .Y(_16392_));
NAND_g _22533_ (.A(_16390_), .B(_16392_), .Y(_16393_));
NAND_g _22534_ (.A(_11217_), .B(_16387_), .Y(_16394_));
AND_g _22535_ (.A(_16393_), .B(_16394_), .Y(_16395_));
NAND_g _22536_ (.A(_00011_[1]), .B(_16395_), .Y(_16396_));
NOR_g _22537_ (.A(_11217_), .B(_16388_), .Y(_16397_));
NAND_g _22538_ (.A(_16389_), .B(_16397_), .Y(_16398_));
NAND_g _22539_ (.A(_11217_), .B(_16384_), .Y(_16399_));
AND_g _22540_ (.A(_16398_), .B(_16399_), .Y(_16400_));
NAND_g _22541_ (.A(_11218_), .B(_16400_), .Y(_16401_));
AND_g _22542_ (.A(_16396_), .B(_16401_), .Y(_16402_));
NAND_g _22543_ (.A(_11220_), .B(_16402_), .Y(_16403_));
NAND_g _22544_ (.A(cpuregs_27[26]), .B(_00011_[1]), .Y(_16404_));
NAND_g _22545_ (.A(cpuregs_25[26]), .B(_11218_), .Y(_16405_));
NAND_g _22546_ (.A(_16404_), .B(_16405_), .Y(_16406_));
NAND_g _22547_ (.A(_11219_), .B(_16406_), .Y(_16407_));
NAND_g _22548_ (.A(cpuregs_31[26]), .B(_00011_[1]), .Y(_16408_));
NAND_g _22549_ (.A(cpuregs_29[26]), .B(_11218_), .Y(_16409_));
NAND_g _22550_ (.A(_16408_), .B(_16409_), .Y(_16410_));
NAND_g _22551_ (.A(_00011_[2]), .B(_16410_), .Y(_16411_));
AND_g _22552_ (.A(_00011_[0]), .B(_16411_), .Y(_16412_));
NAND_g _22553_ (.A(_16407_), .B(_16412_), .Y(_16413_));
NAND_g _22554_ (.A(cpuregs_26[26]), .B(_00011_[1]), .Y(_16414_));
NAND_g _22555_ (.A(cpuregs_24[26]), .B(_11218_), .Y(_16415_));
NAND_g _22556_ (.A(_16414_), .B(_16415_), .Y(_16416_));
NAND_g _22557_ (.A(_11219_), .B(_16416_), .Y(_16417_));
NAND_g _22558_ (.A(cpuregs_30[26]), .B(_00011_[1]), .Y(_16418_));
NAND_g _22559_ (.A(cpuregs_28[26]), .B(_11218_), .Y(_16419_));
NAND_g _22560_ (.A(_16418_), .B(_16419_), .Y(_16420_));
NAND_g _22561_ (.A(_00011_[2]), .B(_16420_), .Y(_16421_));
AND_g _22562_ (.A(_11217_), .B(_16421_), .Y(_16422_));
NAND_g _22563_ (.A(_16417_), .B(_16422_), .Y(_16423_));
AND_g _22564_ (.A(_00011_[3]), .B(_16423_), .Y(_16424_));
NAND_g _22565_ (.A(_16413_), .B(_16424_), .Y(_16425_));
AND_g _22566_ (.A(_16403_), .B(_16425_), .Y(_16426_));
NAND_g _22567_ (.A(cpuregs_1[26]), .B(_11219_), .Y(_16427_));
NAND_g _22568_ (.A(cpuregs_5[26]), .B(_00011_[2]), .Y(_16428_));
AND_g _22569_ (.A(_00011_[0]), .B(_16428_), .Y(_16429_));
NAND_g _22570_ (.A(_16427_), .B(_16429_), .Y(_16430_));
NAND_g _22571_ (.A(cpuregs_0[26]), .B(_11219_), .Y(_16431_));
NAND_g _22572_ (.A(cpuregs_4[26]), .B(_00011_[2]), .Y(_16432_));
AND_g _22573_ (.A(_11217_), .B(_16432_), .Y(_16433_));
NAND_g _22574_ (.A(_16431_), .B(_16433_), .Y(_16434_));
AND_g _22575_ (.A(_11218_), .B(_16434_), .Y(_16435_));
NAND_g _22576_ (.A(_16430_), .B(_16435_), .Y(_16436_));
NAND_g _22577_ (.A(cpuregs_3[26]), .B(_11219_), .Y(_16437_));
NAND_g _22578_ (.A(cpuregs_7[26]), .B(_00011_[2]), .Y(_16438_));
AND_g _22579_ (.A(_00011_[0]), .B(_16438_), .Y(_16439_));
NAND_g _22580_ (.A(_16437_), .B(_16439_), .Y(_16440_));
NAND_g _22581_ (.A(cpuregs_2[26]), .B(_11219_), .Y(_16441_));
NAND_g _22582_ (.A(cpuregs_6[26]), .B(_00011_[2]), .Y(_16442_));
AND_g _22583_ (.A(_11217_), .B(_16442_), .Y(_16443_));
NAND_g _22584_ (.A(_16441_), .B(_16443_), .Y(_16444_));
AND_g _22585_ (.A(_00011_[1]), .B(_16444_), .Y(_16445_));
NAND_g _22586_ (.A(_16440_), .B(_16445_), .Y(_16446_));
NAND_g _22587_ (.A(_16436_), .B(_16446_), .Y(_16447_));
NAND_g _22588_ (.A(_11220_), .B(_16447_), .Y(_16448_));
NAND_g _22589_ (.A(cpuregs_14[26]), .B(_11217_), .Y(_16449_));
NAND_g _22590_ (.A(cpuregs_15[26]), .B(_00011_[0]), .Y(_16450_));
NAND_g _22591_ (.A(_16449_), .B(_16450_), .Y(_16451_));
NAND_g _22592_ (.A(_00011_[2]), .B(_16451_), .Y(_16452_));
NAND_g _22593_ (.A(cpuregs_10[26]), .B(_11217_), .Y(_16453_));
NAND_g _22594_ (.A(cpuregs_11[26]), .B(_00011_[0]), .Y(_16454_));
NAND_g _22595_ (.A(_16453_), .B(_16454_), .Y(_16455_));
NAND_g _22596_ (.A(_11219_), .B(_16455_), .Y(_16456_));
AND_g _22597_ (.A(_16452_), .B(_16456_), .Y(_16457_));
NAND_g _22598_ (.A(cpuregs_12[26]), .B(_11217_), .Y(_16458_));
NAND_g _22599_ (.A(cpuregs_13[26]), .B(_00011_[0]), .Y(_16459_));
NAND_g _22600_ (.A(_16458_), .B(_16459_), .Y(_01699_));
NAND_g _22601_ (.A(_00011_[2]), .B(_01699_), .Y(_01700_));
NAND_g _22602_ (.A(cpuregs_8[26]), .B(_11217_), .Y(_01701_));
NAND_g _22603_ (.A(cpuregs_9[26]), .B(_00011_[0]), .Y(_01702_));
NAND_g _22604_ (.A(_01701_), .B(_01702_), .Y(_01703_));
NAND_g _22605_ (.A(_11219_), .B(_01703_), .Y(_01704_));
AND_g _22606_ (.A(_01700_), .B(_01704_), .Y(_01705_));
NAND_g _22607_ (.A(_11218_), .B(_01705_), .Y(_01706_));
NAND_g _22608_ (.A(_00011_[1]), .B(_16457_), .Y(_01707_));
AND_g _22609_ (.A(_00011_[3]), .B(_01706_), .Y(_01708_));
NAND_g _22610_ (.A(_01707_), .B(_01708_), .Y(_01709_));
NAND_g _22611_ (.A(_00011_[4]), .B(_16426_), .Y(_01710_));
AND_g _22612_ (.A(_11221_), .B(_16448_), .Y(_01711_));
NAND_g _22613_ (.A(_01709_), .B(_01711_), .Y(_01712_));
AND_g _22614_ (.A(_13734_), .B(_01712_), .Y(_01713_));
AND_g _22615_ (.A(_01710_), .B(_01713_), .Y(_01714_));
NAND_g _22616_ (.A(_14358_), .B(_01714_), .Y(_01715_));
AND_g _22617_ (.A(decoded_imm[26]), .B(_13830_), .Y(_01716_));
NAND_g _22618_ (.A(_13409_), .B(_01716_), .Y(_01717_));
AND_g _22619_ (.A(_13727_), .B(_01717_), .Y(_01718_));
NAND_g _22620_ (.A(_01715_), .B(_01718_), .Y(_01719_));
AND_g _22621_ (.A(_16381_), .B(_01719_), .Y(_00529_));
NAND_g _22622_ (.A(_11007_), .B(_13728_), .Y(_01720_));
NAND_g _22623_ (.A(cpuregs_19[27]), .B(_11219_), .Y(_01721_));
NAND_g _22624_ (.A(cpuregs_23[27]), .B(_00011_[2]), .Y(_01722_));
AND_g _22625_ (.A(_00011_[0]), .B(_01722_), .Y(_01723_));
NAND_g _22626_ (.A(_01721_), .B(_01723_), .Y(_01724_));
NAND_g _22627_ (.A(cpuregs_18[27]), .B(_11219_), .Y(_01725_));
NAND_g _22628_ (.A(cpuregs_22[27]), .B(_00011_[2]), .Y(_01726_));
AND_g _22629_ (.A(_11217_), .B(_01726_), .Y(_01727_));
NAND_g _22630_ (.A(_01725_), .B(_01727_), .Y(_01728_));
AND_g _22631_ (.A(_11220_), .B(_01728_), .Y(_01729_));
NAND_g _22632_ (.A(_01724_), .B(_01729_), .Y(_01730_));
NAND_g _22633_ (.A(cpuregs_27[27]), .B(_11219_), .Y(_01731_));
NAND_g _22634_ (.A(cpuregs_31[27]), .B(_00011_[2]), .Y(_01732_));
AND_g _22635_ (.A(_00011_[0]), .B(_01732_), .Y(_01733_));
NAND_g _22636_ (.A(_01731_), .B(_01733_), .Y(_01734_));
NAND_g _22637_ (.A(cpuregs_26[27]), .B(_11219_), .Y(_01735_));
NAND_g _22638_ (.A(cpuregs_30[27]), .B(_00011_[2]), .Y(_01736_));
AND_g _22639_ (.A(_11217_), .B(_01736_), .Y(_01737_));
NAND_g _22640_ (.A(_01735_), .B(_01737_), .Y(_01738_));
AND_g _22641_ (.A(_00011_[3]), .B(_01738_), .Y(_01739_));
NAND_g _22642_ (.A(_01734_), .B(_01739_), .Y(_01740_));
NAND_g _22643_ (.A(_01730_), .B(_01740_), .Y(_01741_));
NAND_g _22644_ (.A(_00011_[1]), .B(_01741_), .Y(_01742_));
NAND_g _22645_ (.A(cpuregs_21[27]), .B(_00011_[2]), .Y(_01743_));
NAND_g _22646_ (.A(cpuregs_17[27]), .B(_11219_), .Y(_01744_));
AND_g _22647_ (.A(_00011_[0]), .B(_01744_), .Y(_01745_));
NAND_g _22648_ (.A(_01743_), .B(_01745_), .Y(_01746_));
NAND_g _22649_ (.A(cpuregs_20[27]), .B(_00011_[2]), .Y(_01747_));
NAND_g _22650_ (.A(cpuregs_16[27]), .B(_11219_), .Y(_01748_));
AND_g _22651_ (.A(_11217_), .B(_01748_), .Y(_01749_));
NAND_g _22652_ (.A(_01747_), .B(_01749_), .Y(_01750_));
AND_g _22653_ (.A(_11220_), .B(_01750_), .Y(_01751_));
NAND_g _22654_ (.A(_01746_), .B(_01751_), .Y(_01752_));
NAND_g _22655_ (.A(cpuregs_25[27]), .B(_11219_), .Y(_01753_));
NAND_g _22656_ (.A(cpuregs_29[27]), .B(_00011_[2]), .Y(_01754_));
AND_g _22657_ (.A(_00011_[0]), .B(_01754_), .Y(_01755_));
NAND_g _22658_ (.A(_01753_), .B(_01755_), .Y(_01756_));
NAND_g _22659_ (.A(cpuregs_24[27]), .B(_11219_), .Y(_01757_));
NAND_g _22660_ (.A(cpuregs_28[27]), .B(_00011_[2]), .Y(_01758_));
AND_g _22661_ (.A(_11217_), .B(_01758_), .Y(_01759_));
NAND_g _22662_ (.A(_01757_), .B(_01759_), .Y(_01760_));
AND_g _22663_ (.A(_00011_[3]), .B(_01760_), .Y(_01761_));
NAND_g _22664_ (.A(_01756_), .B(_01761_), .Y(_01762_));
NAND_g _22665_ (.A(_01752_), .B(_01762_), .Y(_01763_));
NAND_g _22666_ (.A(_11218_), .B(_01763_), .Y(_01764_));
NAND_g _22667_ (.A(_01742_), .B(_01764_), .Y(_01765_));
NAND_g _22668_ (.A(_00011_[4]), .B(_01765_), .Y(_01766_));
NAND_g _22669_ (.A(cpuregs_6[27]), .B(_00011_[2]), .Y(_01767_));
NAND_g _22670_ (.A(cpuregs_2[27]), .B(_11219_), .Y(_01768_));
AND_g _22671_ (.A(_01767_), .B(_01768_), .Y(_01769_));
NAND_g _22672_ (.A(_11217_), .B(_01769_), .Y(_01770_));
NAND_g _22673_ (.A(cpuregs_7[27]), .B(_00011_[2]), .Y(_01771_));
NAND_g _22674_ (.A(cpuregs_3[27]), .B(_11219_), .Y(_01772_));
AND_g _22675_ (.A(_00011_[0]), .B(_01772_), .Y(_01773_));
NAND_g _22676_ (.A(_01771_), .B(_01773_), .Y(_01774_));
AND_g _22677_ (.A(_11220_), .B(_01774_), .Y(_01775_));
NAND_g _22678_ (.A(_01770_), .B(_01775_), .Y(_01776_));
NOR_g _22679_ (.A(cpuregs_10[27]), .B(_00011_[2]), .Y(_01777_));
AND_g _22680_ (.A(_11106_), .B(_00011_[2]), .Y(_01778_));
NOR_g _22681_ (.A(_01777_), .B(_01778_), .Y(_01779_));
NOR_g _22682_ (.A(cpuregs_11[27]), .B(_00011_[2]), .Y(_01780_));
NOT_g _22683_ (.A(_01780_), .Y(_01781_));
NAND_g _22684_ (.A(_11170_), .B(_00011_[2]), .Y(_01782_));
AND_g _22685_ (.A(_00011_[0]), .B(_01782_), .Y(_01783_));
NAND_g _22686_ (.A(_01781_), .B(_01783_), .Y(_01784_));
NAND_g _22687_ (.A(_11217_), .B(_01779_), .Y(_01785_));
NAND_g _22688_ (.A(_01784_), .B(_01785_), .Y(_01786_));
NAND_g _22689_ (.A(_00011_[3]), .B(_01786_), .Y(_01787_));
AND_g _22690_ (.A(_01776_), .B(_01787_), .Y(_01788_));
NAND_g _22691_ (.A(cpuregs_4[27]), .B(_00011_[2]), .Y(_01789_));
NAND_g _22692_ (.A(cpuregs_0[27]), .B(_11219_), .Y(_01790_));
AND_g _22693_ (.A(_01789_), .B(_01790_), .Y(_01791_));
NAND_g _22694_ (.A(_11217_), .B(_01791_), .Y(_01792_));
NAND_g _22695_ (.A(cpuregs_5[27]), .B(_00011_[2]), .Y(_01793_));
NAND_g _22696_ (.A(cpuregs_1[27]), .B(_11219_), .Y(_01794_));
AND_g _22697_ (.A(_00011_[0]), .B(_01794_), .Y(_01795_));
NAND_g _22698_ (.A(_01793_), .B(_01795_), .Y(_01796_));
AND_g _22699_ (.A(_11220_), .B(_01796_), .Y(_01797_));
AND_g _22700_ (.A(_01792_), .B(_01797_), .Y(_01798_));
NAND_g _22701_ (.A(_10936_), .B(_11219_), .Y(_01799_));
NAND_g _22702_ (.A(_11154_), .B(_00011_[2]), .Y(_01800_));
NOR_g _22703_ (.A(cpuregs_8[27]), .B(_00011_[2]), .Y(_01801_));
AND_g _22704_ (.A(_11122_), .B(_00011_[2]), .Y(_01802_));
NOR_g _22705_ (.A(_01801_), .B(_01802_), .Y(_01803_));
AND_g _22706_ (.A(_00011_[0]), .B(_01800_), .Y(_01804_));
NAND_g _22707_ (.A(_01799_), .B(_01804_), .Y(_01805_));
NAND_g _22708_ (.A(_11217_), .B(_01803_), .Y(_01806_));
NAND_g _22709_ (.A(_01805_), .B(_01806_), .Y(_01807_));
AND_g _22710_ (.A(_00011_[3]), .B(_01807_), .Y(_01808_));
NOR_g _22711_ (.A(_01798_), .B(_01808_), .Y(_01809_));
NAND_g _22712_ (.A(_11218_), .B(_01809_), .Y(_01810_));
NAND_g _22713_ (.A(_00011_[1]), .B(_01788_), .Y(_01811_));
AND_g _22714_ (.A(_01810_), .B(_01811_), .Y(_01812_));
NAND_g _22715_ (.A(_11221_), .B(_01812_), .Y(_01813_));
NAND_g _22716_ (.A(_01766_), .B(_01813_), .Y(_01814_));
AND_g _22717_ (.A(_13734_), .B(_01814_), .Y(_01815_));
NAND_g _22718_ (.A(_14358_), .B(_01815_), .Y(_01816_));
AND_g _22719_ (.A(decoded_imm[27]), .B(_13830_), .Y(_01817_));
NAND_g _22720_ (.A(_13409_), .B(_01817_), .Y(_01818_));
AND_g _22721_ (.A(_13727_), .B(_01818_), .Y(_01819_));
NAND_g _22722_ (.A(_01816_), .B(_01819_), .Y(_01820_));
AND_g _22723_ (.A(_01720_), .B(_01820_), .Y(_00530_));
NAND_g _22724_ (.A(_11008_), .B(_13728_), .Y(_01821_));
NAND_g _22725_ (.A(cpuregs_25[28]), .B(_11219_), .Y(_01822_));
NAND_g _22726_ (.A(cpuregs_29[28]), .B(_00011_[2]), .Y(_01823_));
AND_g _22727_ (.A(_00011_[0]), .B(_01823_), .Y(_01824_));
NAND_g _22728_ (.A(_01822_), .B(_01824_), .Y(_01825_));
NAND_g _22729_ (.A(cpuregs_24[28]), .B(_11219_), .Y(_01826_));
NAND_g _22730_ (.A(cpuregs_28[28]), .B(_00011_[2]), .Y(_01827_));
AND_g _22731_ (.A(_11217_), .B(_01827_), .Y(_01828_));
NAND_g _22732_ (.A(_01826_), .B(_01828_), .Y(_01829_));
AND_g _22733_ (.A(_11218_), .B(_01829_), .Y(_01830_));
NAND_g _22734_ (.A(_01825_), .B(_01830_), .Y(_01831_));
NAND_g _22735_ (.A(cpuregs_31[28]), .B(_00011_[2]), .Y(_01832_));
NAND_g _22736_ (.A(cpuregs_27[28]), .B(_11219_), .Y(_01833_));
AND_g _22737_ (.A(_00011_[0]), .B(_01833_), .Y(_01834_));
NAND_g _22738_ (.A(_01832_), .B(_01834_), .Y(_01835_));
NAND_g _22739_ (.A(cpuregs_26[28]), .B(_11219_), .Y(_01836_));
NAND_g _22740_ (.A(cpuregs_30[28]), .B(_00011_[2]), .Y(_01837_));
AND_g _22741_ (.A(_11217_), .B(_01837_), .Y(_01838_));
NAND_g _22742_ (.A(_01836_), .B(_01838_), .Y(_01839_));
AND_g _22743_ (.A(_00011_[1]), .B(_01839_), .Y(_01840_));
NAND_g _22744_ (.A(_01835_), .B(_01840_), .Y(_01841_));
NAND_g _22745_ (.A(_01831_), .B(_01841_), .Y(_01842_));
NAND_g _22746_ (.A(_00011_[3]), .B(_01842_), .Y(_01843_));
NAND_g _22747_ (.A(cpuregs_23[28]), .B(_00011_[2]), .Y(_01844_));
NAND_g _22748_ (.A(cpuregs_19[28]), .B(_11219_), .Y(_01845_));
AND_g _22749_ (.A(_00011_[0]), .B(_01845_), .Y(_01846_));
NAND_g _22750_ (.A(_01844_), .B(_01846_), .Y(_01847_));
NAND_g _22751_ (.A(cpuregs_22[28]), .B(_00011_[2]), .Y(_01848_));
NAND_g _22752_ (.A(cpuregs_18[28]), .B(_11219_), .Y(_01849_));
AND_g _22753_ (.A(_01848_), .B(_01849_), .Y(_01850_));
NAND_g _22754_ (.A(_11217_), .B(_01850_), .Y(_01851_));
AND_g _22755_ (.A(_00011_[1]), .B(_01847_), .Y(_01852_));
NAND_g _22756_ (.A(_01851_), .B(_01852_), .Y(_01853_));
NAND_g _22757_ (.A(cpuregs_21[28]), .B(_00011_[0]), .Y(_01854_));
NAND_g _22758_ (.A(cpuregs_20[28]), .B(_11217_), .Y(_01855_));
NAND_g _22759_ (.A(_01854_), .B(_01855_), .Y(_01856_));
NAND_g _22760_ (.A(_00011_[2]), .B(_01856_), .Y(_01857_));
NAND_g _22761_ (.A(cpuregs_17[28]), .B(_00011_[0]), .Y(_01858_));
NAND_g _22762_ (.A(cpuregs_16[28]), .B(_11217_), .Y(_01859_));
NAND_g _22763_ (.A(_01858_), .B(_01859_), .Y(_01860_));
NAND_g _22764_ (.A(_11219_), .B(_01860_), .Y(_01861_));
NAND_g _22765_ (.A(_01857_), .B(_01861_), .Y(_01862_));
NAND_g _22766_ (.A(_11218_), .B(_01862_), .Y(_01863_));
NAND_g _22767_ (.A(_01853_), .B(_01863_), .Y(_01864_));
NAND_g _22768_ (.A(_11220_), .B(_01864_), .Y(_01865_));
AND_g _22769_ (.A(_01843_), .B(_01865_), .Y(_01866_));
NAND_g _22770_ (.A(cpuregs_1[28]), .B(_11219_), .Y(_01867_));
NAND_g _22771_ (.A(cpuregs_5[28]), .B(_00011_[2]), .Y(_01868_));
AND_g _22772_ (.A(_00011_[0]), .B(_01868_), .Y(_01869_));
NAND_g _22773_ (.A(_01867_), .B(_01869_), .Y(_01870_));
NAND_g _22774_ (.A(cpuregs_0[28]), .B(_11219_), .Y(_01871_));
NAND_g _22775_ (.A(cpuregs_4[28]), .B(_00011_[2]), .Y(_01872_));
AND_g _22776_ (.A(_11217_), .B(_01872_), .Y(_01873_));
NAND_g _22777_ (.A(_01871_), .B(_01873_), .Y(_01874_));
AND_g _22778_ (.A(_11218_), .B(_01874_), .Y(_01875_));
NAND_g _22779_ (.A(_01870_), .B(_01875_), .Y(_01876_));
NAND_g _22780_ (.A(cpuregs_3[28]), .B(_11219_), .Y(_01877_));
NAND_g _22781_ (.A(cpuregs_7[28]), .B(_00011_[2]), .Y(_01878_));
AND_g _22782_ (.A(_00011_[0]), .B(_01878_), .Y(_01879_));
NAND_g _22783_ (.A(_01877_), .B(_01879_), .Y(_01880_));
NAND_g _22784_ (.A(cpuregs_2[28]), .B(_11219_), .Y(_01881_));
NAND_g _22785_ (.A(cpuregs_6[28]), .B(_00011_[2]), .Y(_01882_));
AND_g _22786_ (.A(_11217_), .B(_01882_), .Y(_01883_));
NAND_g _22787_ (.A(_01881_), .B(_01883_), .Y(_01884_));
AND_g _22788_ (.A(_00011_[1]), .B(_01884_), .Y(_01885_));
NAND_g _22789_ (.A(_01880_), .B(_01885_), .Y(_01886_));
NAND_g _22790_ (.A(_01876_), .B(_01886_), .Y(_01887_));
NAND_g _22791_ (.A(_11220_), .B(_01887_), .Y(_01888_));
NAND_g _22792_ (.A(cpuregs_14[28]), .B(_11217_), .Y(_01889_));
NAND_g _22793_ (.A(cpuregs_15[28]), .B(_00011_[0]), .Y(_01890_));
NAND_g _22794_ (.A(_01889_), .B(_01890_), .Y(_01891_));
NAND_g _22795_ (.A(_00011_[2]), .B(_01891_), .Y(_01892_));
NAND_g _22796_ (.A(cpuregs_10[28]), .B(_11217_), .Y(_01893_));
NAND_g _22797_ (.A(cpuregs_11[28]), .B(_00011_[0]), .Y(_01894_));
NAND_g _22798_ (.A(_01893_), .B(_01894_), .Y(_01895_));
NAND_g _22799_ (.A(_11219_), .B(_01895_), .Y(_01896_));
AND_g _22800_ (.A(_01892_), .B(_01896_), .Y(_01897_));
NAND_g _22801_ (.A(cpuregs_12[28]), .B(_11217_), .Y(_01898_));
NAND_g _22802_ (.A(cpuregs_13[28]), .B(_00011_[0]), .Y(_01899_));
NAND_g _22803_ (.A(_01898_), .B(_01899_), .Y(_01900_));
NAND_g _22804_ (.A(_00011_[2]), .B(_01900_), .Y(_01901_));
NAND_g _22805_ (.A(cpuregs_8[28]), .B(_11217_), .Y(_01902_));
NAND_g _22806_ (.A(cpuregs_9[28]), .B(_00011_[0]), .Y(_01903_));
NAND_g _22807_ (.A(_01902_), .B(_01903_), .Y(_01904_));
NAND_g _22808_ (.A(_11219_), .B(_01904_), .Y(_01905_));
AND_g _22809_ (.A(_01901_), .B(_01905_), .Y(_01906_));
NAND_g _22810_ (.A(_11218_), .B(_01906_), .Y(_01907_));
NAND_g _22811_ (.A(_00011_[1]), .B(_01897_), .Y(_01908_));
AND_g _22812_ (.A(_00011_[3]), .B(_01907_), .Y(_01909_));
NAND_g _22813_ (.A(_01908_), .B(_01909_), .Y(_01910_));
NAND_g _22814_ (.A(_00011_[4]), .B(_01866_), .Y(_01911_));
AND_g _22815_ (.A(_11221_), .B(_01888_), .Y(_01912_));
NAND_g _22816_ (.A(_01910_), .B(_01912_), .Y(_01913_));
AND_g _22817_ (.A(_13734_), .B(_01913_), .Y(_01914_));
AND_g _22818_ (.A(_01911_), .B(_01914_), .Y(_01915_));
NAND_g _22819_ (.A(_14358_), .B(_01915_), .Y(_01916_));
AND_g _22820_ (.A(decoded_imm[28]), .B(_13830_), .Y(_01917_));
NAND_g _22821_ (.A(_13409_), .B(_01917_), .Y(_01918_));
AND_g _22822_ (.A(_13727_), .B(_01918_), .Y(_01919_));
NAND_g _22823_ (.A(_01916_), .B(_01919_), .Y(_01920_));
AND_g _22824_ (.A(_01821_), .B(_01920_), .Y(_00531_));
NAND_g _22825_ (.A(_11009_), .B(_13728_), .Y(_01921_));
NAND_g _22826_ (.A(cpuregs_19[29]), .B(_11219_), .Y(_01922_));
NAND_g _22827_ (.A(cpuregs_23[29]), .B(_00011_[2]), .Y(_01923_));
AND_g _22828_ (.A(_00011_[0]), .B(_01923_), .Y(_01924_));
NAND_g _22829_ (.A(_01922_), .B(_01924_), .Y(_01925_));
NAND_g _22830_ (.A(cpuregs_18[29]), .B(_11219_), .Y(_01926_));
NAND_g _22831_ (.A(cpuregs_22[29]), .B(_00011_[2]), .Y(_01927_));
AND_g _22832_ (.A(_11217_), .B(_01927_), .Y(_01928_));
NAND_g _22833_ (.A(_01926_), .B(_01928_), .Y(_01929_));
AND_g _22834_ (.A(_11220_), .B(_01929_), .Y(_01930_));
NAND_g _22835_ (.A(_01925_), .B(_01930_), .Y(_01931_));
NAND_g _22836_ (.A(cpuregs_27[29]), .B(_11219_), .Y(_01932_));
NAND_g _22837_ (.A(cpuregs_31[29]), .B(_00011_[2]), .Y(_01933_));
AND_g _22838_ (.A(_00011_[0]), .B(_01933_), .Y(_01934_));
NAND_g _22839_ (.A(_01932_), .B(_01934_), .Y(_01935_));
NAND_g _22840_ (.A(cpuregs_26[29]), .B(_11219_), .Y(_01936_));
NAND_g _22841_ (.A(cpuregs_30[29]), .B(_00011_[2]), .Y(_01937_));
AND_g _22842_ (.A(_11217_), .B(_01937_), .Y(_01938_));
NAND_g _22843_ (.A(_01936_), .B(_01938_), .Y(_01939_));
AND_g _22844_ (.A(_00011_[3]), .B(_01939_), .Y(_01940_));
NAND_g _22845_ (.A(_01935_), .B(_01940_), .Y(_01941_));
NAND_g _22846_ (.A(_01931_), .B(_01941_), .Y(_01942_));
NAND_g _22847_ (.A(_00011_[1]), .B(_01942_), .Y(_01943_));
NOR_g _22848_ (.A(cpuregs_16[29]), .B(_00011_[2]), .Y(_01944_));
AND_g _22849_ (.A(_11202_), .B(_00011_[2]), .Y(_01945_));
NOR_g _22850_ (.A(_01944_), .B(_01945_), .Y(_01946_));
NOR_g _22851_ (.A(cpuregs_17[29]), .B(_00011_[2]), .Y(_01947_));
NAND_g _22852_ (.A(_11037_), .B(_00011_[2]), .Y(_01948_));
NOR_g _22853_ (.A(cpuregs_24[29]), .B(_00011_[2]), .Y(_01949_));
AND_g _22854_ (.A(_11101_), .B(_00011_[2]), .Y(_01950_));
NOR_g _22855_ (.A(_01949_), .B(_01950_), .Y(_01951_));
NOR_g _22856_ (.A(cpuregs_25[29]), .B(_00011_[2]), .Y(_01952_));
NAND_g _22857_ (.A(_10933_), .B(_00011_[2]), .Y(_01953_));
NAND_g _22858_ (.A(_11217_), .B(_01946_), .Y(_01954_));
NOR_g _22859_ (.A(_11217_), .B(_01947_), .Y(_01955_));
NAND_g _22860_ (.A(_01948_), .B(_01955_), .Y(_01956_));
AND_g _22861_ (.A(_01954_), .B(_01956_), .Y(_01957_));
NAND_g _22862_ (.A(_11220_), .B(_01957_), .Y(_01958_));
NOR_g _22863_ (.A(_11217_), .B(_01952_), .Y(_01959_));
NAND_g _22864_ (.A(_01953_), .B(_01959_), .Y(_01960_));
NAND_g _22865_ (.A(_11217_), .B(_01951_), .Y(_01961_));
AND_g _22866_ (.A(_01960_), .B(_01961_), .Y(_01962_));
NAND_g _22867_ (.A(_00011_[3]), .B(_01962_), .Y(_01963_));
AND_g _22868_ (.A(_01958_), .B(_01963_), .Y(_01964_));
NAND_g _22869_ (.A(_11218_), .B(_01964_), .Y(_01965_));
NAND_g _22870_ (.A(cpuregs_1[29]), .B(_11219_), .Y(_01966_));
NAND_g _22871_ (.A(cpuregs_5[29]), .B(_00011_[2]), .Y(_01967_));
AND_g _22872_ (.A(_00011_[0]), .B(_01967_), .Y(_01968_));
NAND_g _22873_ (.A(_01966_), .B(_01968_), .Y(_01969_));
NAND_g _22874_ (.A(cpuregs_0[29]), .B(_11219_), .Y(_01970_));
NAND_g _22875_ (.A(cpuregs_4[29]), .B(_00011_[2]), .Y(_01971_));
AND_g _22876_ (.A(_11217_), .B(_01971_), .Y(_01972_));
NAND_g _22877_ (.A(_01970_), .B(_01972_), .Y(_01973_));
AND_g _22878_ (.A(_11220_), .B(_01973_), .Y(_01974_));
NAND_g _22879_ (.A(_01969_), .B(_01974_), .Y(_01975_));
NAND_g _22880_ (.A(cpuregs_13[29]), .B(_00011_[2]), .Y(_01976_));
NAND_g _22881_ (.A(cpuregs_9[29]), .B(_11219_), .Y(_01977_));
AND_g _22882_ (.A(_00011_[0]), .B(_01977_), .Y(_01978_));
NAND_g _22883_ (.A(_01976_), .B(_01978_), .Y(_01979_));
NAND_g _22884_ (.A(cpuregs_12[29]), .B(_00011_[2]), .Y(_01980_));
NAND_g _22885_ (.A(cpuregs_8[29]), .B(_11219_), .Y(_01981_));
AND_g _22886_ (.A(_11217_), .B(_01981_), .Y(_01982_));
NAND_g _22887_ (.A(_01980_), .B(_01982_), .Y(_01983_));
AND_g _22888_ (.A(_00011_[3]), .B(_01983_), .Y(_01984_));
NAND_g _22889_ (.A(_01979_), .B(_01984_), .Y(_01985_));
NAND_g _22890_ (.A(_01975_), .B(_01985_), .Y(_01986_));
NAND_g _22891_ (.A(_11218_), .B(_01986_), .Y(_01987_));
NAND_g _22892_ (.A(cpuregs_14[29]), .B(_11217_), .Y(_01988_));
NAND_g _22893_ (.A(cpuregs_15[29]), .B(_00011_[0]), .Y(_01989_));
NAND_g _22894_ (.A(_01988_), .B(_01989_), .Y(_01990_));
NAND_g _22895_ (.A(_00011_[2]), .B(_01990_), .Y(_01991_));
NAND_g _22896_ (.A(cpuregs_10[29]), .B(_11217_), .Y(_01992_));
NAND_g _22897_ (.A(cpuregs_11[29]), .B(_00011_[0]), .Y(_01993_));
NAND_g _22898_ (.A(_01992_), .B(_01993_), .Y(_01994_));
NAND_g _22899_ (.A(_11219_), .B(_01994_), .Y(_01995_));
NAND_g _22900_ (.A(_01991_), .B(_01995_), .Y(_01996_));
NAND_g _22901_ (.A(_00011_[3]), .B(_01996_), .Y(_01997_));
NAND_g _22902_ (.A(cpuregs_6[29]), .B(_11217_), .Y(_01998_));
NAND_g _22903_ (.A(cpuregs_7[29]), .B(_00011_[0]), .Y(_01999_));
NAND_g _22904_ (.A(_01998_), .B(_01999_), .Y(_02000_));
NAND_g _22905_ (.A(_00011_[2]), .B(_02000_), .Y(_02001_));
NAND_g _22906_ (.A(cpuregs_2[29]), .B(_11217_), .Y(_02002_));
NAND_g _22907_ (.A(cpuregs_3[29]), .B(_00011_[0]), .Y(_02003_));
NAND_g _22908_ (.A(_02002_), .B(_02003_), .Y(_02004_));
NAND_g _22909_ (.A(_11219_), .B(_02004_), .Y(_02005_));
NAND_g _22910_ (.A(_02001_), .B(_02005_), .Y(_02006_));
NAND_g _22911_ (.A(_11220_), .B(_02006_), .Y(_02007_));
NAND_g _22912_ (.A(_01997_), .B(_02007_), .Y(_02008_));
NAND_g _22913_ (.A(_00011_[1]), .B(_02008_), .Y(_02009_));
AND_g _22914_ (.A(_01987_), .B(_02009_), .Y(_02010_));
AND_g _22915_ (.A(_00011_[4]), .B(_01943_), .Y(_02011_));
NAND_g _22916_ (.A(_01965_), .B(_02011_), .Y(_02012_));
NAND_g _22917_ (.A(_11221_), .B(_02010_), .Y(_02013_));
AND_g _22918_ (.A(_02012_), .B(_02013_), .Y(_02014_));
AND_g _22919_ (.A(_13734_), .B(_02014_), .Y(_02015_));
NAND_g _22920_ (.A(_13833_), .B(_02015_), .Y(_02016_));
NAND_g _22921_ (.A(decoded_imm[29]), .B(_13830_), .Y(_02017_));
NAND_g _22922_ (.A(_02016_), .B(_02017_), .Y(_02018_));
NAND_g _22923_ (.A(_13409_), .B(_02018_), .Y(_02019_));
AND_g _22924_ (.A(_13724_), .B(_02015_), .Y(_02020_));
NOR_g _22925_ (.A(_13728_), .B(_02020_), .Y(_02021_));
NAND_g _22926_ (.A(_02019_), .B(_02021_), .Y(_02022_));
AND_g _22927_ (.A(_01921_), .B(_02022_), .Y(_00532_));
NAND_g _22928_ (.A(_11010_), .B(_13728_), .Y(_02023_));
NAND_g _22929_ (.A(cpuregs_31[30]), .B(_00011_[1]), .Y(_02024_));
NAND_g _22930_ (.A(cpuregs_29[30]), .B(_11218_), .Y(_02025_));
NAND_g _22931_ (.A(_02024_), .B(_02025_), .Y(_02026_));
NAND_g _22932_ (.A(_00011_[2]), .B(_02026_), .Y(_02027_));
NAND_g _22933_ (.A(cpuregs_27[30]), .B(_00011_[1]), .Y(_02028_));
NAND_g _22934_ (.A(cpuregs_25[30]), .B(_11218_), .Y(_02029_));
NAND_g _22935_ (.A(_02028_), .B(_02029_), .Y(_02030_));
NAND_g _22936_ (.A(_11219_), .B(_02030_), .Y(_02031_));
NAND_g _22937_ (.A(_02027_), .B(_02031_), .Y(_02032_));
NAND_g _22938_ (.A(_00011_[0]), .B(_02032_), .Y(_02033_));
NAND_g _22939_ (.A(cpuregs_30[30]), .B(_00011_[1]), .Y(_02034_));
NAND_g _22940_ (.A(cpuregs_28[30]), .B(_11218_), .Y(_02035_));
NAND_g _22941_ (.A(_02034_), .B(_02035_), .Y(_02036_));
NAND_g _22942_ (.A(_00011_[2]), .B(_02036_), .Y(_02037_));
NAND_g _22943_ (.A(cpuregs_26[30]), .B(_00011_[1]), .Y(_02038_));
NAND_g _22944_ (.A(cpuregs_24[30]), .B(_11218_), .Y(_02039_));
NAND_g _22945_ (.A(_02038_), .B(_02039_), .Y(_02040_));
NAND_g _22946_ (.A(_11219_), .B(_02040_), .Y(_02041_));
NAND_g _22947_ (.A(_02037_), .B(_02041_), .Y(_02042_));
NAND_g _22948_ (.A(_11217_), .B(_02042_), .Y(_02043_));
NAND_g _22949_ (.A(_02033_), .B(_02043_), .Y(_02044_));
NAND_g _22950_ (.A(_00011_[3]), .B(_02044_), .Y(_02045_));
NOR_g _22951_ (.A(cpuregs_18[30]), .B(_00011_[2]), .Y(_02046_));
NOR_g _22952_ (.A(cpuregs_22[30]), .B(_11219_), .Y(_02047_));
NOR_g _22953_ (.A(_02046_), .B(_02047_), .Y(_02048_));
NOR_g _22954_ (.A(cpuregs_16[30]), .B(_00011_[2]), .Y(_02049_));
NOR_g _22955_ (.A(cpuregs_20[30]), .B(_11219_), .Y(_02050_));
NOR_g _22956_ (.A(_02049_), .B(_02050_), .Y(_02051_));
NAND_g _22957_ (.A(_11191_), .B(_00011_[2]), .Y(_02052_));
NOR_g _22958_ (.A(cpuregs_19[30]), .B(_00011_[2]), .Y(_02053_));
NOR_g _22959_ (.A(cpuregs_17[30]), .B(_00011_[2]), .Y(_02054_));
NAND_g _22960_ (.A(_11038_), .B(_00011_[2]), .Y(_02055_));
NOR_g _22961_ (.A(_11217_), .B(_02053_), .Y(_02056_));
NAND_g _22962_ (.A(_02052_), .B(_02056_), .Y(_02057_));
NAND_g _22963_ (.A(_11217_), .B(_02048_), .Y(_02058_));
AND_g _22964_ (.A(_02057_), .B(_02058_), .Y(_02059_));
NAND_g _22965_ (.A(_00011_[1]), .B(_02059_), .Y(_02060_));
NOR_g _22966_ (.A(_11217_), .B(_02054_), .Y(_02061_));
NAND_g _22967_ (.A(_02055_), .B(_02061_), .Y(_02062_));
NAND_g _22968_ (.A(_11217_), .B(_02051_), .Y(_02063_));
AND_g _22969_ (.A(_02062_), .B(_02063_), .Y(_02064_));
NAND_g _22970_ (.A(_11218_), .B(_02064_), .Y(_02065_));
AND_g _22971_ (.A(_11220_), .B(_02065_), .Y(_02066_));
NAND_g _22972_ (.A(_02060_), .B(_02066_), .Y(_02067_));
AND_g _22973_ (.A(_02045_), .B(_02067_), .Y(_02068_));
NAND_g _22974_ (.A(cpuregs_13[30]), .B(_11218_), .Y(_02069_));
NAND_g _22975_ (.A(cpuregs_15[30]), .B(_00011_[1]), .Y(_02070_));
AND_g _22976_ (.A(_00011_[2]), .B(_02070_), .Y(_02071_));
NAND_g _22977_ (.A(_02069_), .B(_02071_), .Y(_02072_));
NAND_g _22978_ (.A(cpuregs_9[30]), .B(_11218_), .Y(_02073_));
NAND_g _22979_ (.A(cpuregs_11[30]), .B(_00011_[1]), .Y(_02074_));
AND_g _22980_ (.A(_11219_), .B(_02074_), .Y(_02075_));
NAND_g _22981_ (.A(_02073_), .B(_02075_), .Y(_02076_));
AND_g _22982_ (.A(_00011_[0]), .B(_02076_), .Y(_02077_));
NAND_g _22983_ (.A(_02072_), .B(_02077_), .Y(_02078_));
NAND_g _22984_ (.A(cpuregs_12[30]), .B(_11218_), .Y(_02079_));
NAND_g _22985_ (.A(cpuregs_14[30]), .B(_00011_[1]), .Y(_02080_));
AND_g _22986_ (.A(_00011_[2]), .B(_02080_), .Y(_02081_));
NAND_g _22987_ (.A(_02079_), .B(_02081_), .Y(_02082_));
NAND_g _22988_ (.A(cpuregs_8[30]), .B(_11218_), .Y(_02083_));
NAND_g _22989_ (.A(cpuregs_10[30]), .B(_00011_[1]), .Y(_02084_));
AND_g _22990_ (.A(_11219_), .B(_02084_), .Y(_02085_));
NAND_g _22991_ (.A(_02083_), .B(_02085_), .Y(_02086_));
AND_g _22992_ (.A(_11217_), .B(_02086_), .Y(_02087_));
NAND_g _22993_ (.A(_02082_), .B(_02087_), .Y(_02088_));
NAND_g _22994_ (.A(_02078_), .B(_02088_), .Y(_02089_));
NAND_g _22995_ (.A(_00011_[3]), .B(_02089_), .Y(_02090_));
NAND_g _22996_ (.A(_10948_), .B(_00011_[2]), .Y(_02091_));
NOR_g _22997_ (.A(cpuregs_2[30]), .B(_00011_[2]), .Y(_02092_));
NOR_g _22998_ (.A(_00011_[0]), .B(_02092_), .Y(_02093_));
NAND_g _22999_ (.A(_02091_), .B(_02093_), .Y(_02094_));
NAND_g _23000_ (.A(_11134_), .B(_00011_[2]), .Y(_02095_));
NOR_g _23001_ (.A(cpuregs_3[30]), .B(_00011_[2]), .Y(_02096_));
NOR_g _23002_ (.A(_11217_), .B(_02096_), .Y(_02097_));
NAND_g _23003_ (.A(_02095_), .B(_02097_), .Y(_02098_));
AND_g _23004_ (.A(_02094_), .B(_02098_), .Y(_02099_));
NAND_g _23005_ (.A(_10960_), .B(_00011_[2]), .Y(_02100_));
NOR_g _23006_ (.A(cpuregs_0[30]), .B(_00011_[2]), .Y(_02101_));
NOR_g _23007_ (.A(_00011_[0]), .B(_02101_), .Y(_02102_));
NAND_g _23008_ (.A(_02100_), .B(_02102_), .Y(_02103_));
NAND_g _23009_ (.A(_11118_), .B(_00011_[2]), .Y(_02104_));
NOR_g _23010_ (.A(cpuregs_1[30]), .B(_00011_[2]), .Y(_02105_));
NOR_g _23011_ (.A(_11217_), .B(_02105_), .Y(_02106_));
NAND_g _23012_ (.A(_02104_), .B(_02106_), .Y(_02107_));
NAND_g _23013_ (.A(_00011_[1]), .B(_02099_), .Y(_02108_));
AND_g _23014_ (.A(_11218_), .B(_02103_), .Y(_02109_));
NAND_g _23015_ (.A(_02107_), .B(_02109_), .Y(_02110_));
AND_g _23016_ (.A(_02108_), .B(_02110_), .Y(_02111_));
NAND_g _23017_ (.A(_11220_), .B(_02111_), .Y(_02112_));
NAND_g _23018_ (.A(_02090_), .B(_02112_), .Y(_02113_));
NAND_g _23019_ (.A(_00011_[4]), .B(_02068_), .Y(_02114_));
NOR_g _23020_ (.A(_00011_[4]), .B(_02113_), .Y(_02115_));
NOR_g _23021_ (.A(_13733_), .B(_02115_), .Y(_02116_));
AND_g _23022_ (.A(_02114_), .B(_02116_), .Y(_02117_));
NAND_g _23023_ (.A(_13833_), .B(_02117_), .Y(_02118_));
NAND_g _23024_ (.A(decoded_imm[30]), .B(_13830_), .Y(_02119_));
NAND_g _23025_ (.A(_02118_), .B(_02119_), .Y(_02120_));
NAND_g _23026_ (.A(_13409_), .B(_02120_), .Y(_02121_));
NAND_g _23027_ (.A(_13724_), .B(_02117_), .Y(_02122_));
AND_g _23028_ (.A(_13727_), .B(_02122_), .Y(_02123_));
NAND_g _23029_ (.A(_02121_), .B(_02123_), .Y(_02124_));
AND_g _23030_ (.A(_02023_), .B(_02124_), .Y(_00533_));
NAND_g _23031_ (.A(_11011_), .B(_13728_), .Y(_02125_));
NOR_g _23032_ (.A(cpuregs_16[31]), .B(_00011_[2]), .Y(_02126_));
NOR_g _23033_ (.A(cpuregs_20[31]), .B(_11219_), .Y(_02127_));
NOR_g _23034_ (.A(_02126_), .B(_02127_), .Y(_02128_));
NOR_g _23035_ (.A(cpuregs_18[31]), .B(_00011_[2]), .Y(_02129_));
NOR_g _23036_ (.A(cpuregs_22[31]), .B(_11219_), .Y(_02130_));
NOR_g _23037_ (.A(_02129_), .B(_02130_), .Y(_02131_));
NOR_g _23038_ (.A(cpuregs_17[31]), .B(_00011_[2]), .Y(_02132_));
NAND_g _23039_ (.A(_11039_), .B(_00011_[2]), .Y(_02133_));
NAND_g _23040_ (.A(_11192_), .B(_00011_[2]), .Y(_02134_));
NOR_g _23041_ (.A(cpuregs_19[31]), .B(_00011_[2]), .Y(_02135_));
NOR_g _23042_ (.A(_11217_), .B(_02135_), .Y(_02136_));
NAND_g _23043_ (.A(_02134_), .B(_02136_), .Y(_02137_));
NAND_g _23044_ (.A(_11217_), .B(_02131_), .Y(_02138_));
AND_g _23045_ (.A(_02137_), .B(_02138_), .Y(_02139_));
NAND_g _23046_ (.A(_00011_[1]), .B(_02139_), .Y(_02140_));
NOR_g _23047_ (.A(_11217_), .B(_02132_), .Y(_02141_));
NAND_g _23048_ (.A(_02133_), .B(_02141_), .Y(_02142_));
NAND_g _23049_ (.A(_11217_), .B(_02128_), .Y(_02143_));
AND_g _23050_ (.A(_02142_), .B(_02143_), .Y(_02144_));
NAND_g _23051_ (.A(_11218_), .B(_02144_), .Y(_02145_));
AND_g _23052_ (.A(_02140_), .B(_02145_), .Y(_02146_));
NAND_g _23053_ (.A(_11220_), .B(_02146_), .Y(_02147_));
NAND_g _23054_ (.A(cpuregs_27[31]), .B(_00011_[1]), .Y(_02148_));
NAND_g _23055_ (.A(cpuregs_25[31]), .B(_11218_), .Y(_02149_));
NAND_g _23056_ (.A(_02148_), .B(_02149_), .Y(_02150_));
NAND_g _23057_ (.A(_11219_), .B(_02150_), .Y(_02151_));
NAND_g _23058_ (.A(cpuregs_31[31]), .B(_00011_[1]), .Y(_02152_));
NAND_g _23059_ (.A(cpuregs_29[31]), .B(_11218_), .Y(_02153_));
NAND_g _23060_ (.A(_02152_), .B(_02153_), .Y(_02154_));
NAND_g _23061_ (.A(_00011_[2]), .B(_02154_), .Y(_02155_));
AND_g _23062_ (.A(_00011_[0]), .B(_02155_), .Y(_02156_));
NAND_g _23063_ (.A(_02151_), .B(_02156_), .Y(_02157_));
NAND_g _23064_ (.A(cpuregs_26[31]), .B(_00011_[1]), .Y(_02158_));
NAND_g _23065_ (.A(cpuregs_24[31]), .B(_11218_), .Y(_02159_));
NAND_g _23066_ (.A(_02158_), .B(_02159_), .Y(_02160_));
NAND_g _23067_ (.A(_11219_), .B(_02160_), .Y(_02161_));
NAND_g _23068_ (.A(cpuregs_30[31]), .B(_00011_[1]), .Y(_02162_));
NAND_g _23069_ (.A(cpuregs_28[31]), .B(_11218_), .Y(_02163_));
NAND_g _23070_ (.A(_02162_), .B(_02163_), .Y(_02164_));
NAND_g _23071_ (.A(_00011_[2]), .B(_02164_), .Y(_02165_));
AND_g _23072_ (.A(_11217_), .B(_02165_), .Y(_02166_));
NAND_g _23073_ (.A(_02161_), .B(_02166_), .Y(_02167_));
AND_g _23074_ (.A(_00011_[3]), .B(_02167_), .Y(_02168_));
NAND_g _23075_ (.A(_02157_), .B(_02168_), .Y(_02169_));
AND_g _23076_ (.A(_02147_), .B(_02169_), .Y(_02170_));
NAND_g _23077_ (.A(cpuregs_1[31]), .B(_11219_), .Y(_02171_));
NAND_g _23078_ (.A(cpuregs_5[31]), .B(_00011_[2]), .Y(_02172_));
AND_g _23079_ (.A(_00011_[0]), .B(_02172_), .Y(_02173_));
NAND_g _23080_ (.A(_02171_), .B(_02173_), .Y(_02174_));
NAND_g _23081_ (.A(cpuregs_0[31]), .B(_11219_), .Y(_02175_));
NAND_g _23082_ (.A(cpuregs_4[31]), .B(_00011_[2]), .Y(_02176_));
AND_g _23083_ (.A(_11217_), .B(_02176_), .Y(_02177_));
NAND_g _23084_ (.A(_02175_), .B(_02177_), .Y(_02178_));
AND_g _23085_ (.A(_11218_), .B(_02178_), .Y(_02179_));
NAND_g _23086_ (.A(_02174_), .B(_02179_), .Y(_02180_));
NAND_g _23087_ (.A(cpuregs_3[31]), .B(_11219_), .Y(_02181_));
NAND_g _23088_ (.A(cpuregs_7[31]), .B(_00011_[2]), .Y(_02182_));
AND_g _23089_ (.A(_00011_[0]), .B(_02182_), .Y(_02183_));
NAND_g _23090_ (.A(_02181_), .B(_02183_), .Y(_02184_));
NAND_g _23091_ (.A(cpuregs_2[31]), .B(_11219_), .Y(_02185_));
NAND_g _23092_ (.A(cpuregs_6[31]), .B(_00011_[2]), .Y(_02186_));
AND_g _23093_ (.A(_11217_), .B(_02186_), .Y(_02187_));
NAND_g _23094_ (.A(_02185_), .B(_02187_), .Y(_02188_));
AND_g _23095_ (.A(_00011_[1]), .B(_02188_), .Y(_02189_));
NAND_g _23096_ (.A(_02184_), .B(_02189_), .Y(_02190_));
NAND_g _23097_ (.A(_02180_), .B(_02190_), .Y(_02191_));
NAND_g _23098_ (.A(_11220_), .B(_02191_), .Y(_02192_));
NAND_g _23099_ (.A(cpuregs_14[31]), .B(_11217_), .Y(_02193_));
NAND_g _23100_ (.A(cpuregs_15[31]), .B(_00011_[0]), .Y(_02194_));
NAND_g _23101_ (.A(_02193_), .B(_02194_), .Y(_02195_));
NAND_g _23102_ (.A(_00011_[2]), .B(_02195_), .Y(_02196_));
NAND_g _23103_ (.A(cpuregs_10[31]), .B(_11217_), .Y(_02197_));
NAND_g _23104_ (.A(cpuregs_11[31]), .B(_00011_[0]), .Y(_02198_));
NAND_g _23105_ (.A(_02197_), .B(_02198_), .Y(_02199_));
NAND_g _23106_ (.A(_11219_), .B(_02199_), .Y(_02200_));
AND_g _23107_ (.A(_02196_), .B(_02200_), .Y(_02201_));
NAND_g _23108_ (.A(cpuregs_12[31]), .B(_11217_), .Y(_02202_));
NAND_g _23109_ (.A(cpuregs_13[31]), .B(_00011_[0]), .Y(_02203_));
NAND_g _23110_ (.A(_02202_), .B(_02203_), .Y(_02204_));
NAND_g _23111_ (.A(_00011_[2]), .B(_02204_), .Y(_02205_));
NAND_g _23112_ (.A(cpuregs_8[31]), .B(_11217_), .Y(_02206_));
NAND_g _23113_ (.A(cpuregs_9[31]), .B(_00011_[0]), .Y(_02207_));
NAND_g _23114_ (.A(_02206_), .B(_02207_), .Y(_02208_));
NAND_g _23115_ (.A(_11219_), .B(_02208_), .Y(_02209_));
AND_g _23116_ (.A(_02205_), .B(_02209_), .Y(_02210_));
NAND_g _23117_ (.A(_11218_), .B(_02210_), .Y(_02211_));
NAND_g _23118_ (.A(_00011_[1]), .B(_02201_), .Y(_02212_));
AND_g _23119_ (.A(_00011_[3]), .B(_02211_), .Y(_02213_));
NAND_g _23120_ (.A(_02212_), .B(_02213_), .Y(_02214_));
NAND_g _23121_ (.A(_00011_[4]), .B(_02170_), .Y(_02215_));
AND_g _23122_ (.A(_11221_), .B(_02192_), .Y(_02216_));
NAND_g _23123_ (.A(_02214_), .B(_02216_), .Y(_02217_));
AND_g _23124_ (.A(_13734_), .B(_02217_), .Y(_02218_));
AND_g _23125_ (.A(_02215_), .B(_02218_), .Y(_02219_));
NAND_g _23126_ (.A(_14358_), .B(_02219_), .Y(_02220_));
AND_g _23127_ (.A(decoded_imm[31]), .B(_13830_), .Y(_02221_));
NAND_g _23128_ (.A(_13409_), .B(_02221_), .Y(_02222_));
AND_g _23129_ (.A(_13727_), .B(_02222_), .Y(_02223_));
NAND_g _23130_ (.A(_02220_), .B(_02223_), .Y(_02224_));
AND_g _23131_ (.A(_02125_), .B(_02224_), .Y(_00534_));
NOR_g _23132_ (.A(mem_do_prefetch), .B(_11916_), .Y(_02225_));
NAND_g _23133_ (.A(_13414_), .B(_02225_), .Y(_02226_));
NOT_g _23134_ (.A(_02226_), .Y(_00535_));
NAND_g _23135_ (.A(_13409_), .B(_13831_), .Y(_02227_));
AND_g _23136_ (.A(_13388_), .B(_13726_), .Y(_02228_));
NOT_g _23137_ (.A(_02228_), .Y(dbg_ascii_state[27]));
NAND_g _23138_ (.A(_11263_), .B(_02228_), .Y(dbg_ascii_state[9]));
AND_g _23139_ (.A(_13390_), .B(dbg_ascii_state[9]), .Y(_02229_));
AND_g _23140_ (.A(_02227_), .B(_02229_), .Y(_02230_));
NOR_g _23141_ (.A(mem_do_rinst), .B(_02230_), .Y(_02231_));
NOR_g _23142_ (.A(_12535_), .B(_02231_), .Y(_02232_));
NAND_g _23143_ (.A(_10901_), .B(_10964_), .Y(_02233_));
NAND_g _23144_ (.A(_10898_), .B(is_sll_srl_sra), .Y(_02234_));
NAND_g _23145_ (.A(_02233_), .B(_02234_), .Y(_02235_));
NAND_g _23146_ (.A(_10980_), .B(_02235_), .Y(_02236_));
NAND_g _23147_ (.A(_13833_), .B(_02236_), .Y(_02237_));
NOR_g _23148_ (.A(_10901_), .B(_13829_), .Y(_02238_));
AND_g _23149_ (.A(is_lb_lh_lw_lbu_lhu), .B(_13610_), .Y(_02239_));
NOR_g _23150_ (.A(_02238_), .B(_02239_), .Y(_02240_));
NAND_g _23151_ (.A(_02237_), .B(_02240_), .Y(_02241_));
NAND_g _23152_ (.A(_13409_), .B(_02241_), .Y(_02242_));
NAND_g _23153_ (.A(mem_do_prefetch), .B(_13416_), .Y(_02243_));
NAND_g _23154_ (.A(_11262_), .B(_12536_), .Y(_02244_));
NAND_g _23155_ (.A(_13724_), .B(_02236_), .Y(_02245_));
AND_g _23156_ (.A(_02243_), .B(_02245_), .Y(_02246_));
AND_g _23157_ (.A(_02230_), .B(_02246_), .Y(_02247_));
AND_g _23158_ (.A(_02244_), .B(_02247_), .Y(_02248_));
NAND_g _23159_ (.A(_02242_), .B(_02248_), .Y(_02249_));
NAND_g _23160_ (.A(_02232_), .B(_02249_), .Y(_02250_));
NOR_g _23161_ (.A(pcpi_rs1[31]), .B(pcpi_rs2[31]), .Y(_02251_));
NAND_g _23162_ (.A(pcpi_rs1[31]), .B(pcpi_rs2[31]), .Y(_02252_));
XOR_g _23163_ (.A(pcpi_rs1[31]), .B(pcpi_rs2[31]), .Y(_02253_));
XNOR_g _23164_ (.A(pcpi_rs1[31]), .B(pcpi_rs2[31]), .Y(_02254_));
NAND_g _23165_ (.A(_11010_), .B(pcpi_rs1[30]), .Y(_02255_));
NOR_g _23166_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_02256_));
NAND_g _23167_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_02257_));
XOR_g _23168_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_02258_));
XNOR_g _23169_ (.A(pcpi_rs2[30]), .B(pcpi_rs1[30]), .Y(_02259_));
NAND_g _23170_ (.A(_11009_), .B(pcpi_rs1[29]), .Y(_02260_));
NOR_g _23171_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_02261_));
AND_g _23172_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_02262_));
NAND_g _23173_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_02263_));
XOR_g _23174_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_02264_));
XNOR_g _23175_ (.A(pcpi_rs2[29]), .B(pcpi_rs1[29]), .Y(_02265_));
AND_g _23176_ (.A(_11008_), .B(pcpi_rs1[28]), .Y(_02266_));
NAND_g _23177_ (.A(_02265_), .B(_02266_), .Y(_02267_));
AND_g _23178_ (.A(_02260_), .B(_02267_), .Y(_02268_));
NAND_g _23179_ (.A(_02260_), .B(_02267_), .Y(_02269_));
NOR_g _23180_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_02270_));
NAND_g _23181_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_02271_));
XOR_g _23182_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_02272_));
XNOR_g _23183_ (.A(pcpi_rs2[28]), .B(pcpi_rs1[28]), .Y(_02273_));
NOR_g _23184_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_02274_));
NOT_g _23185_ (.A(_02274_), .Y(_02275_));
NAND_g _23186_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_02276_));
XOR_g _23187_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_02277_));
XNOR_g _23188_ (.A(pcpi_rs2[27]), .B(pcpi_rs1[27]), .Y(_02278_));
AND_g _23189_ (.A(_11006_), .B(pcpi_rs1[26]), .Y(_02279_));
NAND_g _23190_ (.A(_11006_), .B(pcpi_rs1[26]), .Y(_02280_));
NAND_g _23191_ (.A(_02278_), .B(_02279_), .Y(_02281_));
NAND_g _23192_ (.A(_11007_), .B(pcpi_rs1[27]), .Y(_02282_));
AND_g _23193_ (.A(_02281_), .B(_02282_), .Y(_02283_));
NAND_g _23194_ (.A(_11005_), .B(pcpi_rs1[25]), .Y(_02284_));
NOR_g _23195_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_02285_));
NAND_g _23196_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_02286_));
XOR_g _23197_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_02287_));
XNOR_g _23198_ (.A(pcpi_rs2[25]), .B(pcpi_rs1[25]), .Y(_02288_));
AND_g _23199_ (.A(_11004_), .B(pcpi_rs1[24]), .Y(_02289_));
NAND_g _23200_ (.A(_11004_), .B(pcpi_rs1[24]), .Y(_02290_));
NAND_g _23201_ (.A(_02288_), .B(_02289_), .Y(_02291_));
AND_g _23202_ (.A(_02284_), .B(_02291_), .Y(_02292_));
NAND_g _23203_ (.A(_02284_), .B(_02291_), .Y(_02293_));
NOR_g _23204_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_02294_));
NAND_g _23205_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_02295_));
XOR_g _23206_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_02296_));
XNOR_g _23207_ (.A(pcpi_rs2[24]), .B(pcpi_rs1[24]), .Y(_02297_));
NAND_g _23208_ (.A(_11003_), .B(pcpi_rs1[23]), .Y(_02298_));
NOR_g _23209_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_02299_));
NAND_g _23210_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_02300_));
XOR_g _23211_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_02301_));
XNOR_g _23212_ (.A(pcpi_rs2[23]), .B(pcpi_rs1[23]), .Y(_02302_));
NAND_g _23213_ (.A(_11002_), .B(pcpi_rs1[22]), .Y(_02303_));
NOR_g _23214_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_02304_));
NAND_g _23215_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_02305_));
XOR_g _23216_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_02306_));
XNOR_g _23217_ (.A(pcpi_rs2[22]), .B(pcpi_rs1[22]), .Y(_02307_));
NAND_g _23218_ (.A(_11001_), .B(pcpi_rs1[21]), .Y(_02308_));
NOR_g _23219_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_02309_));
NAND_g _23220_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_02310_));
XOR_g _23221_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_02311_));
XNOR_g _23222_ (.A(pcpi_rs2[21]), .B(pcpi_rs1[21]), .Y(_02312_));
AND_g _23223_ (.A(_11000_), .B(pcpi_rs1[20]), .Y(_02313_));
NAND_g _23224_ (.A(_11000_), .B(pcpi_rs1[20]), .Y(_02314_));
NAND_g _23225_ (.A(_02312_), .B(_02313_), .Y(_02315_));
NAND_g _23226_ (.A(_02308_), .B(_02315_), .Y(_02316_));
NAND_g _23227_ (.A(_02307_), .B(_02316_), .Y(_02317_));
NAND_g _23228_ (.A(_02303_), .B(_02317_), .Y(_02318_));
NAND_g _23229_ (.A(_02302_), .B(_02318_), .Y(_02319_));
AND_g _23230_ (.A(_02298_), .B(_02319_), .Y(_02320_));
AND_g _23231_ (.A(_02302_), .B(_02307_), .Y(_02321_));
NOR_g _23232_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_02322_));
NAND_g _23233_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_02323_));
XOR_g _23234_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_02324_));
XNOR_g _23235_ (.A(pcpi_rs2[20]), .B(pcpi_rs1[20]), .Y(_02325_));
AND_g _23236_ (.A(_02312_), .B(_02325_), .Y(_02326_));
AND_g _23237_ (.A(_02321_), .B(_02326_), .Y(_02327_));
NAND_g _23238_ (.A(_10999_), .B(pcpi_rs1[19]), .Y(_02328_));
NOR_g _23239_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_02329_));
NAND_g _23240_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_02330_));
XOR_g _23241_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_02331_));
XNOR_g _23242_ (.A(pcpi_rs2[19]), .B(pcpi_rs1[19]), .Y(_02332_));
NAND_g _23243_ (.A(_10998_), .B(pcpi_rs1[18]), .Y(_02333_));
NOR_g _23244_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_02334_));
NAND_g _23245_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_02335_));
XOR_g _23246_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_02336_));
XNOR_g _23247_ (.A(pcpi_rs2[18]), .B(pcpi_rs1[18]), .Y(_02337_));
NAND_g _23248_ (.A(_10997_), .B(pcpi_rs1[17]), .Y(_02338_));
NOR_g _23249_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_02339_));
NOT_g _23250_ (.A(_02339_), .Y(_02340_));
NAND_g _23251_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_02341_));
XOR_g _23252_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_02342_));
XNOR_g _23253_ (.A(pcpi_rs2[17]), .B(pcpi_rs1[17]), .Y(_02343_));
AND_g _23254_ (.A(_10996_), .B(pcpi_rs1[16]), .Y(_02344_));
NAND_g _23255_ (.A(_10996_), .B(pcpi_rs1[16]), .Y(_02345_));
NAND_g _23256_ (.A(_02343_), .B(_02344_), .Y(_02346_));
AND_g _23257_ (.A(_02338_), .B(_02346_), .Y(_02347_));
NAND_g _23258_ (.A(_02338_), .B(_02346_), .Y(_02348_));
NAND_g _23259_ (.A(_02337_), .B(_02348_), .Y(_02349_));
NAND_g _23260_ (.A(_02333_), .B(_02349_), .Y(_02350_));
NAND_g _23261_ (.A(_02332_), .B(_02350_), .Y(_02351_));
AND_g _23262_ (.A(_02328_), .B(_02351_), .Y(_02352_));
NOT_g _23263_ (.A(_02352_), .Y(_02353_));
AND_g _23264_ (.A(_02332_), .B(_02337_), .Y(_02354_));
NOR_g _23265_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_02355_));
NAND_g _23266_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_02356_));
XOR_g _23267_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_02357_));
XNOR_g _23268_ (.A(pcpi_rs2[16]), .B(pcpi_rs1[16]), .Y(_02358_));
AND_g _23269_ (.A(_02343_), .B(_02358_), .Y(_02359_));
AND_g _23270_ (.A(_02354_), .B(_02359_), .Y(_02360_));
NOR_g _23271_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_02361_));
NAND_g _23272_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_02362_));
XOR_g _23273_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_02363_));
XNOR_g _23274_ (.A(pcpi_rs2[15]), .B(pcpi_rs1[15]), .Y(_02364_));
NOR_g _23275_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_02365_));
NAND_g _23276_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_02366_));
XOR_g _23277_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_02367_));
XNOR_g _23278_ (.A(pcpi_rs2[14]), .B(pcpi_rs1[14]), .Y(_02368_));
AND_g _23279_ (.A(_02364_), .B(_02368_), .Y(_02369_));
NOR_g _23280_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_02370_));
NAND_g _23281_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_02371_));
XOR_g _23282_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_02372_));
XNOR_g _23283_ (.A(pcpi_rs2[13]), .B(pcpi_rs1[13]), .Y(_02373_));
NOR_g _23284_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_02374_));
NAND_g _23285_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_02375_));
XOR_g _23286_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_02376_));
XNOR_g _23287_ (.A(pcpi_rs2[12]), .B(pcpi_rs1[12]), .Y(_02377_));
AND_g _23288_ (.A(_02373_), .B(_02377_), .Y(_02378_));
NOR_g _23289_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_02379_));
NAND_g _23290_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_02380_));
XOR_g _23291_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_02381_));
XNOR_g _23292_ (.A(pcpi_rs2[11]), .B(pcpi_rs1[11]), .Y(_02382_));
NOR_g _23293_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_02383_));
NAND_g _23294_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_02384_));
XOR_g _23295_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_02385_));
XNOR_g _23296_ (.A(pcpi_rs2[10]), .B(pcpi_rs1[10]), .Y(_02386_));
AND_g _23297_ (.A(_02382_), .B(_02386_), .Y(_02387_));
NOR_g _23298_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_02388_));
NAND_g _23299_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_02389_));
XOR_g _23300_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_02390_));
XNOR_g _23301_ (.A(pcpi_rs2[9]), .B(pcpi_rs1[9]), .Y(_02391_));
NOR_g _23302_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_02392_));
NAND_g _23303_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_02393_));
XOR_g _23304_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_02394_));
XNOR_g _23305_ (.A(pcpi_rs2[7]), .B(pcpi_rs1[7]), .Y(_02395_));
NOR_g _23306_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_02396_));
NOT_g _23307_ (.A(_02396_), .Y(_02397_));
NAND_g _23308_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_02398_));
XOR_g _23309_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_02399_));
XNOR_g _23310_ (.A(pcpi_rs2[6]), .B(pcpi_rs1[6]), .Y(_02400_));
AND_g _23311_ (.A(_02395_), .B(_02400_), .Y(_02401_));
NAND_g _23312_ (.A(_10985_), .B(pcpi_rs1[5]), .Y(_02402_));
NOR_g _23313_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_02403_));
NAND_g _23314_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_02404_));
XOR_g _23315_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_02405_));
XNOR_g _23316_ (.A(pcpi_rs2[5]), .B(pcpi_rs1[5]), .Y(_02406_));
NOR_g _23317_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_02407_));
AND_g _23318_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_02408_));
NAND_g _23319_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_02409_));
XOR_g _23320_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_02410_));
XNOR_g _23321_ (.A(pcpi_rs2[4]), .B(pcpi_rs1[4]), .Y(_02411_));
NAND_g _23322_ (.A(_10983_), .B(pcpi_rs1[2]), .Y(_02412_));
NOR_g _23323_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_02413_));
AND_g _23324_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_02414_));
NAND_g _23325_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_02415_));
XOR_g _23326_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_02416_));
XNOR_g _23327_ (.A(pcpi_rs2[2]), .B(pcpi_rs1[2]), .Y(_02417_));
NAND_g _23328_ (.A(_10982_), .B(pcpi_rs1[1]), .Y(_02418_));
NOR_g _23329_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_02419_));
AND_g _23330_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_02420_));
NAND_g _23331_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_02421_));
XOR_g _23332_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_02422_));
XNOR_g _23333_ (.A(pcpi_rs2[1]), .B(pcpi_rs1[1]), .Y(_02423_));
NOR_g _23334_ (.A(pcpi_rs2[0]), .B(pcpi_rs1[0]), .Y(_02424_));
NAND_g _23335_ (.A(pcpi_rs2[0]), .B(pcpi_rs1[0]), .Y(_02425_));
XNOR_g _23336_ (.A(pcpi_rs2[0]), .B(pcpi_rs1[0]), .Y(_02426_));
NAND_g _23337_ (.A(pcpi_rs2[0]), .B(_11135_), .Y(_02427_));
NAND_g _23338_ (.A(_02423_), .B(_02427_), .Y(_02428_));
NAND_g _23339_ (.A(_02418_), .B(_02428_), .Y(_02429_));
NAND_g _23340_ (.A(_02417_), .B(_02429_), .Y(_02430_));
NAND_g _23341_ (.A(_02412_), .B(_02430_), .Y(_02431_));
NAND_g _23342_ (.A(pcpi_rs1[3]), .B(_02431_), .Y(_02432_));
AND_g _23343_ (.A(pcpi_rs2[3]), .B(_02432_), .Y(_02433_));
NOR_g _23344_ (.A(pcpi_rs1[3]), .B(_02431_), .Y(_02434_));
NOR_g _23345_ (.A(_02433_), .B(_02434_), .Y(_02435_));
NAND_g _23346_ (.A(_02411_), .B(_02435_), .Y(_02436_));
NAND_g _23347_ (.A(_10984_), .B(pcpi_rs1[4]), .Y(_02437_));
NAND_g _23348_ (.A(_02436_), .B(_02437_), .Y(_02438_));
NAND_g _23349_ (.A(_02406_), .B(_02438_), .Y(_02439_));
NAND_g _23350_ (.A(_02402_), .B(_02439_), .Y(_02440_));
NAND_g _23351_ (.A(_02401_), .B(_02440_), .Y(_02441_));
NAND_g _23352_ (.A(_10987_), .B(pcpi_rs1[7]), .Y(_02442_));
AND_g _23353_ (.A(_10986_), .B(pcpi_rs1[6]), .Y(_02443_));
NAND_g _23354_ (.A(_02395_), .B(_02443_), .Y(_02444_));
AND_g _23355_ (.A(_02442_), .B(_02444_), .Y(_02445_));
NAND_g _23356_ (.A(_02441_), .B(_02445_), .Y(_02446_));
NOR_g _23357_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_02447_));
NAND_g _23358_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_02448_));
XOR_g _23359_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_02449_));
XNOR_g _23360_ (.A(pcpi_rs2[8]), .B(pcpi_rs1[8]), .Y(_02450_));
NAND_g _23361_ (.A(_02446_), .B(_02450_), .Y(_02451_));
AND_g _23362_ (.A(_02391_), .B(_02450_), .Y(_02452_));
AND_g _23363_ (.A(_02446_), .B(_02452_), .Y(_02453_));
NAND_g _23364_ (.A(_02446_), .B(_02452_), .Y(_02454_));
NAND_g _23365_ (.A(_02387_), .B(_02453_), .Y(_02455_));
NAND_g _23366_ (.A(_10990_), .B(pcpi_rs1[10]), .Y(_02456_));
NAND_g _23367_ (.A(_10989_), .B(pcpi_rs1[9]), .Y(_02457_));
AND_g _23368_ (.A(_10988_), .B(pcpi_rs1[8]), .Y(_02458_));
NAND_g _23369_ (.A(_02391_), .B(_02458_), .Y(_02459_));
AND_g _23370_ (.A(_02457_), .B(_02459_), .Y(_02460_));
NAND_g _23371_ (.A(_02457_), .B(_02459_), .Y(_02461_));
NAND_g _23372_ (.A(_02386_), .B(_02461_), .Y(_02462_));
NAND_g _23373_ (.A(_02456_), .B(_02462_), .Y(_02463_));
NAND_g _23374_ (.A(_02382_), .B(_02463_), .Y(_02464_));
NAND_g _23375_ (.A(_10991_), .B(pcpi_rs1[11]), .Y(_02465_));
AND_g _23376_ (.A(_02464_), .B(_02465_), .Y(_02466_));
NAND_g _23377_ (.A(_02455_), .B(_02466_), .Y(_02467_));
NAND_g _23378_ (.A(_02377_), .B(_02467_), .Y(_02468_));
NAND_g _23379_ (.A(_02378_), .B(_02467_), .Y(_02469_));
AND_g _23380_ (.A(_02369_), .B(_02378_), .Y(_02470_));
NAND_g _23381_ (.A(_02467_), .B(_02470_), .Y(_02471_));
NAND_g _23382_ (.A(_10993_), .B(pcpi_rs1[13]), .Y(_02472_));
AND_g _23383_ (.A(_10992_), .B(pcpi_rs1[12]), .Y(_02473_));
NAND_g _23384_ (.A(_10992_), .B(pcpi_rs1[12]), .Y(_02474_));
NAND_g _23385_ (.A(_02373_), .B(_02473_), .Y(_02475_));
AND_g _23386_ (.A(_02472_), .B(_02475_), .Y(_02476_));
NAND_g _23387_ (.A(_02472_), .B(_02475_), .Y(_02477_));
NAND_g _23388_ (.A(_02369_), .B(_02477_), .Y(_02478_));
AND_g _23389_ (.A(_10994_), .B(pcpi_rs1[14]), .Y(_02479_));
NAND_g _23390_ (.A(_10994_), .B(pcpi_rs1[14]), .Y(_02480_));
NAND_g _23391_ (.A(_02364_), .B(_02479_), .Y(_02481_));
NAND_g _23392_ (.A(_10995_), .B(pcpi_rs1[15]), .Y(_02482_));
AND_g _23393_ (.A(_02481_), .B(_02482_), .Y(_02483_));
AND_g _23394_ (.A(_02478_), .B(_02483_), .Y(_02484_));
NAND_g _23395_ (.A(_02471_), .B(_02484_), .Y(_02485_));
NAND_g _23396_ (.A(_02360_), .B(_02485_), .Y(_02486_));
NAND_g _23397_ (.A(_02352_), .B(_02486_), .Y(_02487_));
NAND_g _23398_ (.A(_02327_), .B(_02487_), .Y(_02488_));
NAND_g _23399_ (.A(_02320_), .B(_02488_), .Y(_02489_));
AND_g _23400_ (.A(_02297_), .B(_02489_), .Y(_02490_));
NAND_g _23401_ (.A(_02297_), .B(_02489_), .Y(_02491_));
NAND_g _23402_ (.A(_02288_), .B(_02490_), .Y(_02492_));
NAND_g _23403_ (.A(_02292_), .B(_02492_), .Y(_02493_));
NOR_g _23404_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_02494_));
NAND_g _23405_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_02495_));
XOR_g _23406_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_02496_));
XNOR_g _23407_ (.A(pcpi_rs2[26]), .B(pcpi_rs1[26]), .Y(_02497_));
NAND_g _23408_ (.A(_02493_), .B(_02497_), .Y(_02498_));
AND_g _23409_ (.A(_02278_), .B(_02497_), .Y(_02499_));
NAND_g _23410_ (.A(_02493_), .B(_02499_), .Y(_02500_));
NAND_g _23411_ (.A(_02283_), .B(_02500_), .Y(_02501_));
AND_g _23412_ (.A(_02273_), .B(_02501_), .Y(_02502_));
NAND_g _23413_ (.A(_02273_), .B(_02501_), .Y(_02503_));
NAND_g _23414_ (.A(_02265_), .B(_02502_), .Y(_02504_));
NAND_g _23415_ (.A(_02268_), .B(_02504_), .Y(_02505_));
NAND_g _23416_ (.A(_02259_), .B(_02505_), .Y(_02506_));
AND_g _23417_ (.A(_02255_), .B(_02506_), .Y(_02507_));
NAND_g _23418_ (.A(_02255_), .B(_02506_), .Y(_02508_));
AND_g _23419_ (.A(_02254_), .B(_02259_), .Y(_02509_));
AND_g _23420_ (.A(_02265_), .B(_02273_), .Y(_02510_));
AND_g _23421_ (.A(_02509_), .B(_02510_), .Y(_02511_));
AND_g _23422_ (.A(_02288_), .B(_02297_), .Y(_02512_));
AND_g _23423_ (.A(_02499_), .B(_02512_), .Y(_02513_));
AND_g _23424_ (.A(_02511_), .B(_02513_), .Y(_02514_));
AND_g _23425_ (.A(_02327_), .B(_02360_), .Y(_02515_));
AND_g _23426_ (.A(_02514_), .B(_02515_), .Y(_02516_));
NAND_g _23427_ (.A(_02485_), .B(_02516_), .Y(_02517_));
NAND_g _23428_ (.A(_02293_), .B(_02499_), .Y(_02518_));
NAND_g _23429_ (.A(_02283_), .B(_02518_), .Y(_02519_));
AND_g _23430_ (.A(_02511_), .B(_02519_), .Y(_02520_));
NAND_g _23431_ (.A(_02269_), .B(_02509_), .Y(_02521_));
NAND_g _23432_ (.A(pcpi_rs1[31]), .B(_11011_), .Y(_02522_));
NOR_g _23433_ (.A(_02253_), .B(_02255_), .Y(_02523_));
AND_g _23434_ (.A(_02521_), .B(_02522_), .Y(_02524_));
NOR_g _23435_ (.A(_02520_), .B(_02523_), .Y(_02525_));
NAND_g _23436_ (.A(_02327_), .B(_02353_), .Y(_02526_));
NAND_g _23437_ (.A(_02320_), .B(_02526_), .Y(_02527_));
NAND_g _23438_ (.A(_02514_), .B(_02527_), .Y(_02528_));
AND_g _23439_ (.A(_02524_), .B(_02528_), .Y(_02529_));
AND_g _23440_ (.A(_02525_), .B(_02529_), .Y(_02530_));
AND_g _23441_ (.A(_02517_), .B(_02530_), .Y(_02531_));
NAND_g _23442_ (.A(_02517_), .B(_02530_), .Y(_02532_));
NAND_g _23443_ (.A(_02254_), .B(_02507_), .Y(_02533_));
NAND_g _23444_ (.A(_02522_), .B(_02533_), .Y(_02534_));
AND_g _23445_ (.A(_02522_), .B(_02533_), .Y(_02535_));
NAND_g _23446_ (.A(is_slti_blt_slt), .B(_02534_), .Y(_02536_));
NAND_g _23447_ (.A(instr_bge), .B(_02535_), .Y(_02537_));
NAND_g _23448_ (.A(is_sltiu_bltu_sltu), .B(_02531_), .Y(_02538_));
NAND_g _23449_ (.A(instr_bgeu), .B(_02532_), .Y(_02539_));
AND_g _23450_ (.A(_02423_), .B(_02426_), .Y(_02540_));
NOR_g _23451_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_02541_));
AND_g _23452_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_02542_));
NAND_g _23453_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_02543_));
XOR_g _23454_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_02544_));
XNOR_g _23455_ (.A(pcpi_rs2[3]), .B(pcpi_rs1[3]), .Y(_02545_));
AND_g _23456_ (.A(_02417_), .B(_02540_), .Y(_02546_));
AND_g _23457_ (.A(_02545_), .B(_02546_), .Y(_02547_));
AND_g _23458_ (.A(_02387_), .B(_02401_), .Y(_02548_));
AND_g _23459_ (.A(_02406_), .B(_02411_), .Y(_02549_));
AND_g _23460_ (.A(_02452_), .B(_02549_), .Y(_02550_));
AND_g _23461_ (.A(_02548_), .B(_02550_), .Y(_02551_));
AND_g _23462_ (.A(_02470_), .B(_02551_), .Y(_02552_));
AND_g _23463_ (.A(_02516_), .B(_02552_), .Y(_02553_));
AND_g _23464_ (.A(_02547_), .B(_02553_), .Y(_02554_));
NAND_g _23465_ (.A(_02547_), .B(_02553_), .Y(_02555_));
NAND_g _23466_ (.A(instr_beq), .B(_02554_), .Y(_02556_));
NAND_g _23467_ (.A(instr_bne), .B(_02555_), .Y(_02557_));
AND_g _23468_ (.A(_02556_), .B(_02557_), .Y(_02558_));
AND_g _23469_ (.A(_02539_), .B(_02558_), .Y(_02559_));
AND_g _23470_ (.A(_02538_), .B(_02559_), .Y(_02560_));
AND_g _23471_ (.A(_02537_), .B(_02560_), .Y(_02561_));
NAND_g _23472_ (.A(_02536_), .B(_02561_), .Y(_02562_));
AND_g _23473_ (.A(resetn), .B(_11271_), .Y(_02563_));
NAND_g _23474_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(_02562_), .Y(_02564_));
AND_g _23475_ (.A(_02562_), .B(_02563_), .Y(_02565_));
NAND_g _23476_ (.A(_02562_), .B(_02563_), .Y(_02566_));
NAND_g _23477_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(_02565_), .Y(_02567_));
NAND_g _23478_ (.A(_02250_), .B(_02567_), .Y(_00536_));
AND_g _23479_ (.A(resetn), .B(_13428_), .Y(_02568_));
NOT_g _23480_ (.A(_02568_), .Y(_02569_));
NAND_g _23481_ (.A(mem_do_rdata), .B(_12534_), .Y(_02570_));
NAND_g _23482_ (.A(_02569_), .B(_02570_), .Y(_00537_));
NAND_g _23483_ (.A(resetn), .B(_13430_), .Y(_02571_));
NAND_g _23484_ (.A(mem_do_wdata), .B(_12534_), .Y(_02572_));
NAND_g _23485_ (.A(_02571_), .B(_02572_), .Y(_00538_));
NOR_g _23486_ (.A(instr_lb), .B(instr_lh), .Y(_02573_));
NOR_g _23487_ (.A(instr_lbu), .B(instr_lhu), .Y(_02574_));
AND_g _23488_ (.A(_10965_), .B(_02574_), .Y(_02575_));
NOT_g _23489_ (.A(_02575_), .Y(_00005_));
AND_g _23490_ (.A(_10965_), .B(_02573_), .Y(_02576_));
AND_g _23491_ (.A(_02574_), .B(_02576_), .Y(_02577_));
NAND_g _23492_ (.A(_13428_), .B(_02577_), .Y(_02578_));
NAND_g _23493_ (.A(_13430_), .B(_13585_), .Y(_02579_));
NAND_g _23494_ (.A(_11263_), .B(_13413_), .Y(dbg_ascii_state[18]));
AND_g _23495_ (.A(_02578_), .B(dbg_ascii_state[18]), .Y(_02580_));
AND_g _23496_ (.A(_02579_), .B(_02580_), .Y(_02581_));
AND_g _23497_ (.A(_13406_), .B(_02581_), .Y(_02582_));
NOR_g _23498_ (.A(_13429_), .B(_13579_), .Y(_02583_));
AND_g _23499_ (.A(instr_sh), .B(_13430_), .Y(_02584_));
NOR_g _23500_ (.A(_02583_), .B(_02584_), .Y(_02585_));
NOR_g _23501_ (.A(mem_wordsize[0]), .B(_02582_), .Y(_02586_));
AND_g _23502_ (.A(_02582_), .B(_02585_), .Y(_02587_));
NOR_g _23503_ (.A(_02586_), .B(_02587_), .Y(_00539_));
NOR_g _23504_ (.A(_13429_), .B(_13578_), .Y(_02588_));
AND_g _23505_ (.A(instr_sb), .B(_13430_), .Y(_02589_));
NOR_g _23506_ (.A(_02588_), .B(_02589_), .Y(_02590_));
AND_g _23507_ (.A(_02582_), .B(_02590_), .Y(_02591_));
NOR_g _23508_ (.A(mem_wordsize[1]), .B(_02582_), .Y(_02592_));
NOR_g _23509_ (.A(_02591_), .B(_02592_), .Y(_00540_));
NOR_g _23510_ (.A(mem_do_rinst), .B(mem_do_prefetch), .Y(_02593_));
NAND_g _23511_ (.A(_10898_), .B(_10901_), .Y(_02594_));
NAND_g _23512_ (.A(_10901_), .B(_11908_), .Y(_02595_));
AND_g _23513_ (.A(_11907_), .B(_02593_), .Y(_02596_));
NAND_g _23514_ (.A(_11907_), .B(_02593_), .Y(_02597_));
NOR_g _23515_ (.A(_10963_), .B(trap), .Y(_02598_));
AND_g _23516_ (.A(_11912_), .B(_02598_), .Y(_02599_));
AND_g _23517_ (.A(mem_do_wdata), .B(_11912_), .Y(_02600_));
AND_g _23518_ (.A(resetn), .B(_02600_), .Y(mem_la_write));
AND_g _23519_ (.A(_11912_), .B(_02595_), .Y(_02601_));
AND_g _23520_ (.A(resetn), .B(_02601_), .Y(mem_la_read));
AND_g _23521_ (.A(_02597_), .B(_02599_), .Y(_02602_));
NAND_g _23522_ (.A(_02597_), .B(_02599_), .Y(_02603_));
NAND_g _23523_ (.A(_02596_), .B(_02599_), .Y(_02604_));
XOR_g _23524_ (.A(mem_state[0]), .B(mem_state[1]), .Y(_02605_));
AND_g _23525_ (.A(_11911_), .B(_02598_), .Y(_02606_));
NAND_g _23526_ (.A(_02605_), .B(_02606_), .Y(_02607_));
AND_g _23527_ (.A(_02604_), .B(_02607_), .Y(_02608_));
NAND_g _23528_ (.A(resetn), .B(trap), .Y(_02609_));
NOR_g _23529_ (.A(mem_ready), .B(_02609_), .Y(_02610_));
AND_g _23530_ (.A(_11903_), .B(_02598_), .Y(_02611_));
NOR_g _23531_ (.A(_02610_), .B(_02611_), .Y(_02612_));
NAND_g _23532_ (.A(_02608_), .B(_02612_), .Y(_02613_));
NAND_g _23533_ (.A(mem_valid), .B(_02613_), .Y(_02614_));
NAND_g _23534_ (.A(_02603_), .B(_02614_), .Y(_00541_));
NAND_g _23535_ (.A(cpu_state[7]), .B(_11259_), .Y(_02615_));
NOR_g _23536_ (.A(cpu_state[6]), .B(_02615_), .Y(_02616_));
NAND_g _23537_ (.A(_11258_), .B(_02616_), .Y(_02617_));
NOR_g _23538_ (.A(_10963_), .B(_02617_), .Y(_00542_));
AND_g _23539_ (.A(_11263_), .B(_11272_), .Y(_02618_));
NAND_g _23540_ (.A(latched_store), .B(_02618_), .Y(_02619_));
NAND_g _23541_ (.A(_13409_), .B(_13566_), .Y(_02620_));
AND_g _23542_ (.A(_13388_), .B(_13403_), .Y(_02621_));
AND_g _23543_ (.A(_02620_), .B(_02621_), .Y(_02622_));
AND_g _23544_ (.A(_02619_), .B(_02622_), .Y(_02623_));
NAND_g _23545_ (.A(_11274_), .B(_02623_), .Y(_02624_));
NAND_g _23546_ (.A(resetn), .B(_02624_), .Y(_02625_));
NAND_g _23547_ (.A(_02566_), .B(_02625_), .Y(_00543_));
NOR_g _23548_ (.A(latched_stalu), .B(_11273_), .Y(_02626_));
NOT_g _23549_ (.A(_02626_), .Y(_02627_));
AND_g _23550_ (.A(_12549_), .B(_02627_), .Y(_00544_));
NAND_g _23551_ (.A(latched_branch), .B(_02618_), .Y(_02628_));
NAND_g _23552_ (.A(instr_jalr), .B(_11273_), .Y(_02629_));
NAND_g _23553_ (.A(instr_jal), .B(launch_next_insn), .Y(_02630_));
AND_g _23554_ (.A(_02628_), .B(_02629_), .Y(_02631_));
NAND_g _23555_ (.A(_02630_), .B(_02631_), .Y(_02632_));
NAND_g _23556_ (.A(resetn), .B(_02632_), .Y(_02633_));
NAND_g _23557_ (.A(_02567_), .B(_02633_), .Y(_00545_));
NOR_g _23558_ (.A(_11042_), .B(_11835_), .Y(_02634_));
AND_g _23559_ (.A(_11765_), .B(_02634_), .Y(_02635_));
NAND_g _23560_ (.A(_11765_), .B(_02634_), .Y(_02636_));
NAND_g _23561_ (.A(_11301_), .B(_02635_), .Y(_02637_));
NAND_g _23562_ (.A(cpuregs_22[0]), .B(_02636_), .Y(_02638_));
NAND_g _23563_ (.A(_02637_), .B(_02638_), .Y(_00546_));
NAND_g _23564_ (.A(_11310_), .B(_02635_), .Y(_02639_));
NAND_g _23565_ (.A(cpuregs_22[1]), .B(_02636_), .Y(_02640_));
NAND_g _23566_ (.A(_02639_), .B(_02640_), .Y(_00547_));
NAND_g _23567_ (.A(_11319_), .B(_02635_), .Y(_02641_));
NAND_g _23568_ (.A(cpuregs_22[2]), .B(_02636_), .Y(_02642_));
NAND_g _23569_ (.A(_02641_), .B(_02642_), .Y(_00548_));
NAND_g _23570_ (.A(_11332_), .B(_02635_), .Y(_02643_));
NAND_g _23571_ (.A(cpuregs_22[3]), .B(_02636_), .Y(_02644_));
NAND_g _23572_ (.A(_02643_), .B(_02644_), .Y(_00549_));
NAND_g _23573_ (.A(_11345_), .B(_02635_), .Y(_02645_));
NAND_g _23574_ (.A(cpuregs_22[4]), .B(_02636_), .Y(_02646_));
NAND_g _23575_ (.A(_02645_), .B(_02646_), .Y(_00550_));
NAND_g _23576_ (.A(_11358_), .B(_02635_), .Y(_02647_));
NAND_g _23577_ (.A(cpuregs_22[5]), .B(_02636_), .Y(_02648_));
NAND_g _23578_ (.A(_02647_), .B(_02648_), .Y(_00551_));
NAND_g _23579_ (.A(_11371_), .B(_02635_), .Y(_02649_));
NAND_g _23580_ (.A(cpuregs_22[6]), .B(_02636_), .Y(_02650_));
NAND_g _23581_ (.A(_02649_), .B(_02650_), .Y(_00552_));
NAND_g _23582_ (.A(_11384_), .B(_02635_), .Y(_02651_));
NAND_g _23583_ (.A(cpuregs_22[7]), .B(_02636_), .Y(_02652_));
NAND_g _23584_ (.A(_02651_), .B(_02652_), .Y(_00553_));
NAND_g _23585_ (.A(_11397_), .B(_02635_), .Y(_02653_));
NAND_g _23586_ (.A(cpuregs_22[8]), .B(_02636_), .Y(_02654_));
NAND_g _23587_ (.A(_02653_), .B(_02654_), .Y(_00554_));
NAND_g _23588_ (.A(_11410_), .B(_02635_), .Y(_02655_));
NAND_g _23589_ (.A(cpuregs_22[9]), .B(_02636_), .Y(_02656_));
NAND_g _23590_ (.A(_02655_), .B(_02656_), .Y(_00555_));
NAND_g _23591_ (.A(_11423_), .B(_02635_), .Y(_02657_));
NAND_g _23592_ (.A(cpuregs_22[10]), .B(_02636_), .Y(_02658_));
NAND_g _23593_ (.A(_02657_), .B(_02658_), .Y(_00556_));
NAND_g _23594_ (.A(_11436_), .B(_02635_), .Y(_02659_));
NAND_g _23595_ (.A(cpuregs_22[11]), .B(_02636_), .Y(_02660_));
NAND_g _23596_ (.A(_02659_), .B(_02660_), .Y(_00557_));
NAND_g _23597_ (.A(_11449_), .B(_02635_), .Y(_02661_));
NAND_g _23598_ (.A(cpuregs_22[12]), .B(_02636_), .Y(_02662_));
NAND_g _23599_ (.A(_02661_), .B(_02662_), .Y(_00558_));
NAND_g _23600_ (.A(_11462_), .B(_02635_), .Y(_02663_));
NAND_g _23601_ (.A(cpuregs_22[13]), .B(_02636_), .Y(_02664_));
NAND_g _23602_ (.A(_02663_), .B(_02664_), .Y(_00559_));
NAND_g _23603_ (.A(_11475_), .B(_02635_), .Y(_02665_));
NAND_g _23604_ (.A(cpuregs_22[14]), .B(_02636_), .Y(_02666_));
NAND_g _23605_ (.A(_02665_), .B(_02666_), .Y(_00560_));
NAND_g _23606_ (.A(_11488_), .B(_02635_), .Y(_02667_));
NAND_g _23607_ (.A(cpuregs_22[15]), .B(_02636_), .Y(_02668_));
NAND_g _23608_ (.A(_02667_), .B(_02668_), .Y(_00561_));
NAND_g _23609_ (.A(_11501_), .B(_02635_), .Y(_02669_));
NAND_g _23610_ (.A(cpuregs_22[16]), .B(_02636_), .Y(_02670_));
NAND_g _23611_ (.A(_02669_), .B(_02670_), .Y(_00562_));
AND_g _23612_ (.A(_11017_), .B(_02636_), .Y(_02671_));
NOR_g _23613_ (.A(_11514_), .B(_02636_), .Y(_02672_));
NOR_g _23614_ (.A(_02671_), .B(_02672_), .Y(_00563_));
NAND_g _23615_ (.A(_11527_), .B(_02635_), .Y(_02673_));
NAND_g _23616_ (.A(cpuregs_22[18]), .B(_02636_), .Y(_02674_));
NAND_g _23617_ (.A(_02673_), .B(_02674_), .Y(_00564_));
NAND_g _23618_ (.A(_11540_), .B(_02635_), .Y(_02675_));
NAND_g _23619_ (.A(cpuregs_22[19]), .B(_02636_), .Y(_02676_));
NAND_g _23620_ (.A(_02675_), .B(_02676_), .Y(_00565_));
NAND_g _23621_ (.A(_11553_), .B(_02635_), .Y(_02677_));
NAND_g _23622_ (.A(cpuregs_22[20]), .B(_02636_), .Y(_02678_));
NAND_g _23623_ (.A(_02677_), .B(_02678_), .Y(_00566_));
NAND_g _23624_ (.A(_11566_), .B(_02635_), .Y(_02679_));
NAND_g _23625_ (.A(cpuregs_22[21]), .B(_02636_), .Y(_02680_));
NAND_g _23626_ (.A(_02679_), .B(_02680_), .Y(_00567_));
NAND_g _23627_ (.A(_11579_), .B(_02635_), .Y(_02681_));
NAND_g _23628_ (.A(cpuregs_22[22]), .B(_02636_), .Y(_02682_));
NAND_g _23629_ (.A(_02681_), .B(_02682_), .Y(_00568_));
NAND_g _23630_ (.A(_11592_), .B(_02635_), .Y(_02683_));
NAND_g _23631_ (.A(cpuregs_22[23]), .B(_02636_), .Y(_02684_));
NAND_g _23632_ (.A(_02683_), .B(_02684_), .Y(_00569_));
NAND_g _23633_ (.A(_11605_), .B(_02635_), .Y(_02685_));
NAND_g _23634_ (.A(cpuregs_22[24]), .B(_02636_), .Y(_02686_));
NAND_g _23635_ (.A(_02685_), .B(_02686_), .Y(_00570_));
NAND_g _23636_ (.A(_11618_), .B(_02635_), .Y(_02687_));
NAND_g _23637_ (.A(cpuregs_22[25]), .B(_02636_), .Y(_02688_));
NAND_g _23638_ (.A(_02687_), .B(_02688_), .Y(_00571_));
NAND_g _23639_ (.A(_11631_), .B(_02635_), .Y(_02689_));
NAND_g _23640_ (.A(cpuregs_22[26]), .B(_02636_), .Y(_02690_));
NAND_g _23641_ (.A(_02689_), .B(_02690_), .Y(_00572_));
NAND_g _23642_ (.A(_11644_), .B(_02635_), .Y(_02691_));
NAND_g _23643_ (.A(cpuregs_22[27]), .B(_02636_), .Y(_02692_));
NAND_g _23644_ (.A(_02691_), .B(_02692_), .Y(_00573_));
NAND_g _23645_ (.A(_11657_), .B(_02635_), .Y(_02693_));
NAND_g _23646_ (.A(cpuregs_22[28]), .B(_02636_), .Y(_02694_));
NAND_g _23647_ (.A(_02693_), .B(_02694_), .Y(_00574_));
NAND_g _23648_ (.A(_11670_), .B(_02635_), .Y(_02695_));
NAND_g _23649_ (.A(cpuregs_22[29]), .B(_02636_), .Y(_02696_));
NAND_g _23650_ (.A(_02695_), .B(_02696_), .Y(_00575_));
NAND_g _23651_ (.A(_11683_), .B(_02635_), .Y(_02697_));
NAND_g _23652_ (.A(cpuregs_22[30]), .B(_02636_), .Y(_02698_));
NAND_g _23653_ (.A(_02697_), .B(_02698_), .Y(_00576_));
NAND_g _23654_ (.A(_11695_), .B(_02635_), .Y(_02699_));
NAND_g _23655_ (.A(cpuregs_22[31]), .B(_02636_), .Y(_02700_));
NAND_g _23656_ (.A(_02699_), .B(_02700_), .Y(_00577_));
AND_g _23657_ (.A(_11289_), .B(_02634_), .Y(_02701_));
NAND_g _23658_ (.A(_11289_), .B(_02634_), .Y(_02702_));
NAND_g _23659_ (.A(cpuregs_21[0]), .B(_02702_), .Y(_02703_));
NAND_g _23660_ (.A(_11301_), .B(_02701_), .Y(_02704_));
NAND_g _23661_ (.A(_02703_), .B(_02704_), .Y(_00578_));
NAND_g _23662_ (.A(cpuregs_21[1]), .B(_02702_), .Y(_02705_));
NAND_g _23663_ (.A(_11310_), .B(_02701_), .Y(_02706_));
NAND_g _23664_ (.A(_02705_), .B(_02706_), .Y(_00579_));
NAND_g _23665_ (.A(cpuregs_21[2]), .B(_02702_), .Y(_02707_));
NAND_g _23666_ (.A(_11319_), .B(_02701_), .Y(_02708_));
NAND_g _23667_ (.A(_02707_), .B(_02708_), .Y(_00580_));
NAND_g _23668_ (.A(cpuregs_21[3]), .B(_02702_), .Y(_02709_));
NAND_g _23669_ (.A(_11332_), .B(_02701_), .Y(_02710_));
NAND_g _23670_ (.A(_02709_), .B(_02710_), .Y(_00581_));
NAND_g _23671_ (.A(cpuregs_21[4]), .B(_02702_), .Y(_02711_));
NAND_g _23672_ (.A(_11345_), .B(_02701_), .Y(_02712_));
NAND_g _23673_ (.A(_02711_), .B(_02712_), .Y(_00582_));
NAND_g _23674_ (.A(cpuregs_21[5]), .B(_02702_), .Y(_02713_));
NAND_g _23675_ (.A(_11358_), .B(_02701_), .Y(_02714_));
NAND_g _23676_ (.A(_02713_), .B(_02714_), .Y(_00583_));
NAND_g _23677_ (.A(cpuregs_21[6]), .B(_02702_), .Y(_02715_));
NAND_g _23678_ (.A(_11371_), .B(_02701_), .Y(_02716_));
NAND_g _23679_ (.A(_02715_), .B(_02716_), .Y(_00584_));
NAND_g _23680_ (.A(cpuregs_21[7]), .B(_02702_), .Y(_02717_));
NAND_g _23681_ (.A(_11384_), .B(_02701_), .Y(_02718_));
NAND_g _23682_ (.A(_02717_), .B(_02718_), .Y(_00585_));
NAND_g _23683_ (.A(cpuregs_21[8]), .B(_02702_), .Y(_02719_));
NAND_g _23684_ (.A(_11397_), .B(_02701_), .Y(_02720_));
NAND_g _23685_ (.A(_02719_), .B(_02720_), .Y(_00586_));
NAND_g _23686_ (.A(cpuregs_21[9]), .B(_02702_), .Y(_02721_));
NAND_g _23687_ (.A(_11410_), .B(_02701_), .Y(_02722_));
NAND_g _23688_ (.A(_02721_), .B(_02722_), .Y(_00587_));
NAND_g _23689_ (.A(cpuregs_21[10]), .B(_02702_), .Y(_02723_));
NAND_g _23690_ (.A(_11423_), .B(_02701_), .Y(_02724_));
NAND_g _23691_ (.A(_02723_), .B(_02724_), .Y(_00588_));
NAND_g _23692_ (.A(cpuregs_21[11]), .B(_02702_), .Y(_02725_));
NAND_g _23693_ (.A(_11436_), .B(_02701_), .Y(_02726_));
NAND_g _23694_ (.A(_02725_), .B(_02726_), .Y(_00589_));
NAND_g _23695_ (.A(cpuregs_21[12]), .B(_02702_), .Y(_02727_));
NAND_g _23696_ (.A(_11449_), .B(_02701_), .Y(_02728_));
NAND_g _23697_ (.A(_02727_), .B(_02728_), .Y(_00590_));
NAND_g _23698_ (.A(cpuregs_21[13]), .B(_02702_), .Y(_02729_));
NAND_g _23699_ (.A(_11462_), .B(_02701_), .Y(_02730_));
NAND_g _23700_ (.A(_02729_), .B(_02730_), .Y(_00591_));
NAND_g _23701_ (.A(cpuregs_21[14]), .B(_02702_), .Y(_02731_));
NAND_g _23702_ (.A(_11475_), .B(_02701_), .Y(_02732_));
NAND_g _23703_ (.A(_02731_), .B(_02732_), .Y(_00592_));
NAND_g _23704_ (.A(cpuregs_21[15]), .B(_02702_), .Y(_02733_));
NAND_g _23705_ (.A(_11488_), .B(_02701_), .Y(_02734_));
NAND_g _23706_ (.A(_02733_), .B(_02734_), .Y(_00593_));
NAND_g _23707_ (.A(cpuregs_21[16]), .B(_02702_), .Y(_02735_));
NAND_g _23708_ (.A(_11501_), .B(_02701_), .Y(_02736_));
NAND_g _23709_ (.A(_02735_), .B(_02736_), .Y(_00594_));
AND_g _23710_ (.A(_11031_), .B(_02702_), .Y(_02737_));
NOR_g _23711_ (.A(_11514_), .B(_02702_), .Y(_02738_));
NOR_g _23712_ (.A(_02737_), .B(_02738_), .Y(_00595_));
NAND_g _23713_ (.A(cpuregs_21[18]), .B(_02702_), .Y(_02739_));
NAND_g _23714_ (.A(_11527_), .B(_02701_), .Y(_02740_));
NAND_g _23715_ (.A(_02739_), .B(_02740_), .Y(_00596_));
NAND_g _23716_ (.A(cpuregs_21[19]), .B(_02702_), .Y(_02741_));
NAND_g _23717_ (.A(_11540_), .B(_02701_), .Y(_02742_));
NAND_g _23718_ (.A(_02741_), .B(_02742_), .Y(_00597_));
NAND_g _23719_ (.A(cpuregs_21[20]), .B(_02702_), .Y(_02743_));
NAND_g _23720_ (.A(_11553_), .B(_02701_), .Y(_02744_));
NAND_g _23721_ (.A(_02743_), .B(_02744_), .Y(_00598_));
NAND_g _23722_ (.A(cpuregs_21[21]), .B(_02702_), .Y(_02745_));
NAND_g _23723_ (.A(_11566_), .B(_02701_), .Y(_02746_));
NAND_g _23724_ (.A(_02745_), .B(_02746_), .Y(_00599_));
NAND_g _23725_ (.A(cpuregs_21[22]), .B(_02702_), .Y(_02747_));
NAND_g _23726_ (.A(_11579_), .B(_02701_), .Y(_02748_));
NAND_g _23727_ (.A(_02747_), .B(_02748_), .Y(_00600_));
NAND_g _23728_ (.A(cpuregs_21[23]), .B(_02702_), .Y(_02749_));
NAND_g _23729_ (.A(_11592_), .B(_02701_), .Y(_02750_));
NAND_g _23730_ (.A(_02749_), .B(_02750_), .Y(_00601_));
NAND_g _23731_ (.A(cpuregs_21[24]), .B(_02702_), .Y(_02751_));
NAND_g _23732_ (.A(_11605_), .B(_02701_), .Y(_02752_));
NAND_g _23733_ (.A(_02751_), .B(_02752_), .Y(_00602_));
NAND_g _23734_ (.A(cpuregs_21[25]), .B(_02702_), .Y(_02753_));
NAND_g _23735_ (.A(_11618_), .B(_02701_), .Y(_02754_));
NAND_g _23736_ (.A(_02753_), .B(_02754_), .Y(_00603_));
NAND_g _23737_ (.A(cpuregs_21[26]), .B(_02702_), .Y(_02755_));
NAND_g _23738_ (.A(_11631_), .B(_02701_), .Y(_02756_));
NAND_g _23739_ (.A(_02755_), .B(_02756_), .Y(_00604_));
NAND_g _23740_ (.A(cpuregs_21[27]), .B(_02702_), .Y(_02757_));
NAND_g _23741_ (.A(_11644_), .B(_02701_), .Y(_02758_));
NAND_g _23742_ (.A(_02757_), .B(_02758_), .Y(_00605_));
NAND_g _23743_ (.A(cpuregs_21[28]), .B(_02702_), .Y(_02759_));
NAND_g _23744_ (.A(_11657_), .B(_02701_), .Y(_02760_));
NAND_g _23745_ (.A(_02759_), .B(_02760_), .Y(_00606_));
NAND_g _23746_ (.A(cpuregs_21[29]), .B(_02702_), .Y(_02761_));
NAND_g _23747_ (.A(_11670_), .B(_02701_), .Y(_02762_));
NAND_g _23748_ (.A(_02761_), .B(_02762_), .Y(_00607_));
NAND_g _23749_ (.A(cpuregs_21[30]), .B(_02702_), .Y(_02763_));
NAND_g _23750_ (.A(_11683_), .B(_02701_), .Y(_02764_));
NAND_g _23751_ (.A(_02763_), .B(_02764_), .Y(_00608_));
NAND_g _23752_ (.A(cpuregs_21[31]), .B(_02702_), .Y(_02765_));
NAND_g _23753_ (.A(_11695_), .B(_02701_), .Y(_02766_));
NAND_g _23754_ (.A(_02765_), .B(_02766_), .Y(_00609_));
NAND_g _23755_ (.A(is_lbu_lhu_lw), .B(_02568_), .Y(_02767_));
AND_g _23756_ (.A(_11263_), .B(_13403_), .Y(_02768_));
AND_g _23757_ (.A(_11263_), .B(_13429_), .Y(_02769_));
AND_g _23758_ (.A(latched_is_lu), .B(resetn), .Y(_02770_));
NAND_g _23759_ (.A(_02769_), .B(_02770_), .Y(_02771_));
NAND_g _23760_ (.A(_02767_), .B(_02771_), .Y(_00610_));
NAND_g _23761_ (.A(instr_lh), .B(_02568_), .Y(_02772_));
AND_g _23762_ (.A(latched_is_lh), .B(resetn), .Y(_02773_));
NAND_g _23763_ (.A(_02769_), .B(_02773_), .Y(_02774_));
NAND_g _23764_ (.A(_02772_), .B(_02774_), .Y(_00611_));
NAND_g _23765_ (.A(instr_lb), .B(_02568_), .Y(_02775_));
AND_g _23766_ (.A(latched_is_lb), .B(resetn), .Y(_02776_));
NAND_g _23767_ (.A(_02769_), .B(_02776_), .Y(_02777_));
NAND_g _23768_ (.A(_02775_), .B(_02777_), .Y(_00612_));
NAND_g _23769_ (.A(decoded_imm_j[11]), .B(_11223_), .Y(_02778_));
NAND_g _23770_ (.A(cached_insn_rs2[0]), .B(decoder_pseudo_trigger_q), .Y(_02779_));
NOR_g _23771_ (.A(q_insn_rs2[0]), .B(dbg_next), .Y(_02780_));
AND_g _23772_ (.A(dbg_next), .B(_02779_), .Y(_02781_));
AND_g _23773_ (.A(_02778_), .B(_02781_), .Y(_02782_));
NOR_g _23774_ (.A(_02780_), .B(_02782_), .Y(_00613_));
NAND_g _23775_ (.A(decoded_imm_j[1]), .B(_11223_), .Y(_02783_));
NAND_g _23776_ (.A(cached_insn_rs2[1]), .B(decoder_pseudo_trigger_q), .Y(_02784_));
NOR_g _23777_ (.A(dbg_next), .B(q_insn_rs2[1]), .Y(_02785_));
AND_g _23778_ (.A(dbg_next), .B(_02784_), .Y(_02786_));
AND_g _23779_ (.A(_02783_), .B(_02786_), .Y(_02787_));
NOR_g _23780_ (.A(_02785_), .B(_02787_), .Y(_00614_));
NAND_g _23781_ (.A(decoded_imm_j[2]), .B(_11223_), .Y(_02788_));
NAND_g _23782_ (.A(cached_insn_rs2[2]), .B(decoder_pseudo_trigger_q), .Y(_02789_));
NOR_g _23783_ (.A(dbg_next), .B(q_insn_rs2[2]), .Y(_02790_));
AND_g _23784_ (.A(dbg_next), .B(_02789_), .Y(_02791_));
AND_g _23785_ (.A(_02788_), .B(_02791_), .Y(_02792_));
NOR_g _23786_ (.A(_02790_), .B(_02792_), .Y(_00615_));
NAND_g _23787_ (.A(decoded_imm_j[3]), .B(_11223_), .Y(_02793_));
NAND_g _23788_ (.A(cached_insn_rs2[3]), .B(decoder_pseudo_trigger_q), .Y(_02794_));
NOR_g _23789_ (.A(dbg_next), .B(q_insn_rs2[3]), .Y(_02795_));
AND_g _23790_ (.A(dbg_next), .B(_02794_), .Y(_02796_));
AND_g _23791_ (.A(_02793_), .B(_02796_), .Y(_02797_));
NOR_g _23792_ (.A(_02795_), .B(_02797_), .Y(_00616_));
NAND_g _23793_ (.A(decoded_imm_j[4]), .B(_11223_), .Y(_02798_));
NAND_g _23794_ (.A(cached_insn_rs2[4]), .B(decoder_pseudo_trigger_q), .Y(_02799_));
NOR_g _23795_ (.A(dbg_next), .B(q_insn_rs2[4]), .Y(_02800_));
AND_g _23796_ (.A(dbg_next), .B(_02799_), .Y(_02801_));
AND_g _23797_ (.A(_02798_), .B(_02801_), .Y(_02802_));
NOR_g _23798_ (.A(_02800_), .B(_02802_), .Y(_00617_));
NOR_g _23799_ (.A(_10963_), .B(_02618_), .Y(_02803_));
NAND_g _23800_ (.A(_11274_), .B(_02803_), .Y(_02804_));
NAND_g _23801_ (.A(latched_rd[0]), .B(_02804_), .Y(_02805_));
NAND_g _23802_ (.A(decoded_rd[0]), .B(_11275_), .Y(_02806_));
NAND_g _23803_ (.A(_02805_), .B(_02806_), .Y(_00618_));
NAND_g _23804_ (.A(latched_rd[1]), .B(_02804_), .Y(_02807_));
NAND_g _23805_ (.A(decoded_rd[1]), .B(_11275_), .Y(_02808_));
NAND_g _23806_ (.A(_02807_), .B(_02808_), .Y(_00619_));
NAND_g _23807_ (.A(latched_rd[2]), .B(_02804_), .Y(_02809_));
NAND_g _23808_ (.A(decoded_rd[2]), .B(_11275_), .Y(_02810_));
NAND_g _23809_ (.A(_02809_), .B(_02810_), .Y(_00620_));
NAND_g _23810_ (.A(latched_rd[3]), .B(_02804_), .Y(_02811_));
NAND_g _23811_ (.A(decoded_rd[3]), .B(_11275_), .Y(_02812_));
NAND_g _23812_ (.A(_02811_), .B(_02812_), .Y(_00621_));
NAND_g _23813_ (.A(latched_rd[4]), .B(_02804_), .Y(_02813_));
NAND_g _23814_ (.A(decoded_rd[4]), .B(_11275_), .Y(_02814_));
NAND_g _23815_ (.A(_02813_), .B(_02814_), .Y(_00622_));
NAND_g _23816_ (.A(_11040_), .B(q_ascii_instr[0]), .Y(_02815_));
AND_g _23817_ (.A(_10907_), .B(_13418_), .Y(_02816_));
AND_g _23818_ (.A(_13575_), .B(_02816_), .Y(_02817_));
NOR_g _23819_ (.A(instr_bne), .B(instr_beq), .Y(_02818_));
NOR_g _23820_ (.A(instr_jal), .B(_12519_), .Y(_02819_));
NAND_g _23821_ (.A(_10962_), .B(_12520_), .Y(_02820_));
NAND_g _23822_ (.A(_02818_), .B(_02820_), .Y(_02821_));
NAND_g _23823_ (.A(instr_jalr), .B(_02818_), .Y(_02822_));
AND_g _23824_ (.A(_10921_), .B(_02822_), .Y(_02823_));
NAND_g _23825_ (.A(_02821_), .B(_02823_), .Y(_02824_));
NAND_g _23826_ (.A(_13569_), .B(_02824_), .Y(_02825_));
NAND_g _23827_ (.A(_02573_), .B(_02825_), .Y(_02826_));
NAND_g _23828_ (.A(_02575_), .B(_02826_), .Y(_02827_));
NAND_g _23829_ (.A(_13585_), .B(_02827_), .Y(_02828_));
AND_g _23830_ (.A(_10913_), .B(_13580_), .Y(_02829_));
NOR_g _23831_ (.A(instr_xori), .B(instr_sltiu), .Y(_02830_));
AND_g _23832_ (.A(_10915_), .B(_13598_), .Y(_02831_));
AND_g _23833_ (.A(_13580_), .B(_02831_), .Y(_02832_));
NAND_g _23834_ (.A(_13587_), .B(_02830_), .Y(_02833_));
AND_g _23835_ (.A(_13587_), .B(_02832_), .Y(_02834_));
AND_g _23836_ (.A(_13417_), .B(_02834_), .Y(_02835_));
AND_g _23837_ (.A(_10912_), .B(_13598_), .Y(_02836_));
AND_g _23838_ (.A(_13583_), .B(_13598_), .Y(_02837_));
AND_g _23839_ (.A(_10968_), .B(_02835_), .Y(_02838_));
NAND_g _23840_ (.A(_02828_), .B(_02838_), .Y(_02839_));
NAND_g _23841_ (.A(_13596_), .B(_02839_), .Y(_02840_));
NAND_g _23842_ (.A(_10908_), .B(_02840_), .Y(_02841_));
NAND_g _23843_ (.A(_02817_), .B(_02841_), .Y(_02842_));
NAND_g _23844_ (.A(instr_sra), .B(_13575_), .Y(_02843_));
AND_g _23845_ (.A(_10972_), .B(_02843_), .Y(_02844_));
NAND_g _23846_ (.A(_02842_), .B(_02844_), .Y(_02845_));
AND_g _23847_ (.A(_13564_), .B(_02845_), .Y(_02846_));
NAND_g _23848_ (.A(_13564_), .B(_02845_), .Y(_02847_));
NAND_g _23849_ (.A(_11223_), .B(_02847_), .Y(_02848_));
NAND_g _23850_ (.A(_11050_), .B(decoder_pseudo_trigger_q), .Y(_02849_));
AND_g _23851_ (.A(dbg_next), .B(_02849_), .Y(_02850_));
NAND_g _23852_ (.A(_02848_), .B(_02850_), .Y(_02851_));
NAND_g _23853_ (.A(_02815_), .B(_02851_), .Y(_00623_));
NAND_g _23854_ (.A(_11040_), .B(q_ascii_instr[1]), .Y(_02852_));
NOR_g _23855_ (.A(instr_bge), .B(instr_beq), .Y(_02853_));
AND_g _23856_ (.A(_13570_), .B(_02853_), .Y(_02854_));
NOR_g _23857_ (.A(instr_bltu), .B(instr_jalr), .Y(_02855_));
AND_g _23858_ (.A(_02854_), .B(_02855_), .Y(_02856_));
AND_g _23859_ (.A(instr_auipc), .B(_10962_), .Y(_02857_));
AND_g _23860_ (.A(_02856_), .B(_02857_), .Y(_02858_));
NAND_g _23861_ (.A(instr_jalr), .B(_02854_), .Y(_02859_));
NOR_g _23862_ (.A(instr_bltu), .B(_02859_), .Y(_02860_));
NOR_g _23863_ (.A(_02858_), .B(_02860_), .Y(_02861_));
NOR_g _23864_ (.A(instr_bgeu), .B(_02861_), .Y(_02862_));
NOR_g _23865_ (.A(instr_lb), .B(_02862_), .Y(_02863_));
NOR_g _23866_ (.A(instr_lh), .B(_02863_), .Y(_02864_));
NOR_g _23867_ (.A(instr_lw), .B(_02864_), .Y(_02865_));
NOT_g _23868_ (.A(_02865_), .Y(_02866_));
NAND_g _23869_ (.A(_02574_), .B(_02866_), .Y(_02867_));
NAND_g _23870_ (.A(_13584_), .B(_02867_), .Y(_02868_));
AND_g _23871_ (.A(_12522_), .B(_02835_), .Y(_02869_));
NAND_g _23872_ (.A(instr_sh), .B(_10968_), .Y(_02870_));
AND_g _23873_ (.A(_02869_), .B(_02870_), .Y(_02871_));
NAND_g _23874_ (.A(_02868_), .B(_02871_), .Y(_02872_));
NAND_g _23875_ (.A(_10910_), .B(_02872_), .Y(_02873_));
NAND_g _23876_ (.A(_13594_), .B(_02873_), .Y(_02874_));
NAND_g _23877_ (.A(_10907_), .B(_02874_), .Y(_02875_));
NAND_g _23878_ (.A(_13418_), .B(_02875_), .Y(_02876_));
AND_g _23879_ (.A(_10904_), .B(_02876_), .Y(_02877_));
NOT_g _23880_ (.A(_02877_), .Y(_02878_));
NOR_g _23881_ (.A(instr_and), .B(instr_rdcycle), .Y(_02879_));
AND_g _23882_ (.A(_10903_), .B(_13563_), .Y(_02880_));
NAND_g _23883_ (.A(_02878_), .B(_02880_), .Y(_02881_));
NAND_g _23884_ (.A(_10974_), .B(_02881_), .Y(_02882_));
NAND_g _23885_ (.A(_10975_), .B(_02882_), .Y(_02883_));
NAND_g _23886_ (.A(_11223_), .B(_02883_), .Y(_02884_));
NAND_g _23887_ (.A(_11051_), .B(decoder_pseudo_trigger_q), .Y(_02885_));
AND_g _23888_ (.A(dbg_next), .B(_02885_), .Y(_02886_));
NAND_g _23889_ (.A(_02884_), .B(_02886_), .Y(_02887_));
NAND_g _23890_ (.A(_02852_), .B(_02887_), .Y(_00624_));
NAND_g _23891_ (.A(_11040_), .B(q_ascii_instr[2]), .Y(_02888_));
NAND_g _23892_ (.A(instr_jal), .B(_13567_), .Y(_02889_));
NAND_g _23893_ (.A(_13571_), .B(_02889_), .Y(_02890_));
NAND_g _23894_ (.A(_02573_), .B(_02890_), .Y(_02891_));
NAND_g _23895_ (.A(_02575_), .B(_02891_), .Y(_02892_));
NAND_g _23896_ (.A(_13589_), .B(_02892_), .Y(_02893_));
NAND_g _23897_ (.A(instr_sw), .B(_13587_), .Y(_02894_));
AND_g _23898_ (.A(_10915_), .B(_02894_), .Y(_02895_));
NAND_g _23899_ (.A(_02893_), .B(_02895_), .Y(_02896_));
NAND_g _23900_ (.A(_02837_), .B(_02896_), .Y(_02897_));
NAND_g _23901_ (.A(_10911_), .B(_02897_), .Y(_02898_));
NAND_g _23902_ (.A(_10910_), .B(_02898_), .Y(_02899_));
NAND_g _23903_ (.A(_13591_), .B(_02899_), .Y(_02900_));
NAND_g _23904_ (.A(_10907_), .B(_02900_), .Y(_02901_));
AND_g _23905_ (.A(_10906_), .B(_02901_), .Y(_02902_));
NOT_g _23906_ (.A(_02902_), .Y(_02903_));
AND_g _23907_ (.A(_10905_), .B(_13575_), .Y(_02904_));
NAND_g _23908_ (.A(_02903_), .B(_02904_), .Y(_02905_));
NAND_g _23909_ (.A(_02879_), .B(_02905_), .Y(_02906_));
AND_g _23910_ (.A(_13564_), .B(_02906_), .Y(_02907_));
NAND_g _23911_ (.A(_13564_), .B(_02906_), .Y(_02908_));
NAND_g _23912_ (.A(_11223_), .B(_02908_), .Y(_02909_));
NAND_g _23913_ (.A(_11052_), .B(decoder_pseudo_trigger_q), .Y(_02910_));
AND_g _23914_ (.A(dbg_next), .B(_02910_), .Y(_02911_));
NAND_g _23915_ (.A(_02909_), .B(_02911_), .Y(_02912_));
NAND_g _23916_ (.A(_02888_), .B(_02912_), .Y(_00625_));
NAND_g _23917_ (.A(_11040_), .B(q_ascii_instr[3]), .Y(_02913_));
NAND_g _23918_ (.A(instr_rdcycleh), .B(_10974_), .Y(_02914_));
AND_g _23919_ (.A(_10975_), .B(_02914_), .Y(_02915_));
NOR_g _23920_ (.A(instr_rdinstrh), .B(decoder_pseudo_trigger_q), .Y(_02916_));
AND_g _23921_ (.A(_02914_), .B(_02916_), .Y(_02917_));
AND_g _23922_ (.A(_10961_), .B(instr_lui), .Y(_02918_));
NOR_g _23923_ (.A(instr_jal), .B(_02918_), .Y(_02919_));
NOR_g _23924_ (.A(instr_lb), .B(_02919_), .Y(_02920_));
AND_g _23925_ (.A(_13573_), .B(_02920_), .Y(_02921_));
NOR_g _23926_ (.A(instr_lh), .B(_02921_), .Y(_02922_));
NAND_g _23927_ (.A(_10966_), .B(_02575_), .Y(_02923_));
NOR_g _23928_ (.A(_02922_), .B(_02923_), .Y(_02924_));
NOR_g _23929_ (.A(instr_sh), .B(_02924_), .Y(_02925_));
NAND_g _23930_ (.A(_13587_), .B(_02925_), .Y(_02926_));
NAND_g _23931_ (.A(_02895_), .B(_02926_), .Y(_02927_));
NAND_g _23932_ (.A(_02837_), .B(_02927_), .Y(_02928_));
NAND_g _23933_ (.A(_12522_), .B(_02928_), .Y(_02929_));
NAND_g _23934_ (.A(_10909_), .B(_02929_), .Y(_02930_));
AND_g _23935_ (.A(_13593_), .B(_02930_), .Y(_02931_));
NOR_g _23936_ (.A(instr_srl), .B(_02931_), .Y(_02932_));
NOT_g _23937_ (.A(_02932_), .Y(_02933_));
NOR_g _23938_ (.A(instr_rdcycle), .B(instr_rdinstr), .Y(_02934_));
NOT_g _23939_ (.A(_02934_), .Y(_02935_));
AND_g _23940_ (.A(_10974_), .B(_13563_), .Y(_02936_));
AND_g _23941_ (.A(_02904_), .B(_02936_), .Y(_02937_));
NAND_g _23942_ (.A(_02933_), .B(_02937_), .Y(_02938_));
NAND_g _23943_ (.A(_02917_), .B(_02938_), .Y(_02939_));
NAND_g _23944_ (.A(_11053_), .B(decoder_pseudo_trigger_q), .Y(_02940_));
AND_g _23945_ (.A(dbg_next), .B(_02940_), .Y(_02941_));
NAND_g _23946_ (.A(_02939_), .B(_02941_), .Y(_02942_));
NAND_g _23947_ (.A(_02913_), .B(_02942_), .Y(_00626_));
NAND_g _23948_ (.A(_11040_), .B(q_ascii_instr[4]), .Y(_02943_));
NAND_g _23949_ (.A(_10921_), .B(instr_bne), .Y(_02944_));
AND_g _23950_ (.A(_10920_), .B(_02944_), .Y(_02945_));
NAND_g _23951_ (.A(_13572_), .B(_02945_), .Y(_02946_));
NAND_g _23952_ (.A(_13568_), .B(_02946_), .Y(_02947_));
NAND_g _23953_ (.A(_02573_), .B(_02947_), .Y(_02948_));
NAND_g _23954_ (.A(_02575_), .B(_02948_), .Y(_02949_));
NAND_g _23955_ (.A(_13589_), .B(_02949_), .Y(_02950_));
NAND_g _23956_ (.A(_02895_), .B(_02950_), .Y(_02951_));
AND_g _23957_ (.A(_13596_), .B(_02837_), .Y(_02952_));
NAND_g _23958_ (.A(_02951_), .B(_02952_), .Y(_02953_));
NAND_g _23959_ (.A(_13593_), .B(_02953_), .Y(_02954_));
NAND_g _23960_ (.A(_13418_), .B(_02954_), .Y(_02955_));
NAND_g _23961_ (.A(_10904_), .B(_02955_), .Y(_02956_));
NAND_g _23962_ (.A(_02880_), .B(_02956_), .Y(_02957_));
NAND_g _23963_ (.A(_10974_), .B(_02957_), .Y(_02958_));
NAND_g _23964_ (.A(_10975_), .B(_02958_), .Y(_02959_));
NAND_g _23965_ (.A(_11223_), .B(_02959_), .Y(_02960_));
NAND_g _23966_ (.A(_11054_), .B(decoder_pseudo_trigger_q), .Y(_02961_));
AND_g _23967_ (.A(dbg_next), .B(_02961_), .Y(_02962_));
NAND_g _23968_ (.A(_02960_), .B(_02962_), .Y(_02963_));
NAND_g _23969_ (.A(_02943_), .B(_02963_), .Y(_00627_));
NAND_g _23970_ (.A(_11040_), .B(q_ascii_instr[8]), .Y(_02964_));
AND_g _23971_ (.A(instr_rdcycleh), .B(_13562_), .Y(_02965_));
NOR_g _23972_ (.A(decoder_pseudo_trigger_q), .B(_02965_), .Y(_02966_));
NOR_g _23973_ (.A(instr_jalr), .B(_02919_), .Y(_02967_));
NOT_g _23974_ (.A(_02967_), .Y(_02968_));
NAND_g _23975_ (.A(_02853_), .B(_02968_), .Y(_02969_));
NOR_g _23976_ (.A(instr_bge), .B(_13570_), .Y(_02970_));
NOR_g _23977_ (.A(instr_bltu), .B(_02970_), .Y(_02971_));
NAND_g _23978_ (.A(_02969_), .B(_02971_), .Y(_02972_));
NAND_g _23979_ (.A(_10918_), .B(_02972_), .Y(_02973_));
NAND_g _23980_ (.A(_02577_), .B(_02973_), .Y(_02974_));
NAND_g _23981_ (.A(_13585_), .B(_02974_), .Y(_02975_));
NAND_g _23982_ (.A(_13587_), .B(_02975_), .Y(_02976_));
NAND_g _23983_ (.A(_10915_), .B(_02976_), .Y(_02977_));
NAND_g _23984_ (.A(_02837_), .B(_02977_), .Y(_02978_));
NAND_g _23985_ (.A(_10971_), .B(_02978_), .Y(_02979_));
NAND_g _23986_ (.A(_10911_), .B(_02979_), .Y(_02980_));
NAND_g _23987_ (.A(_10910_), .B(_02980_), .Y(_02981_));
NAND_g _23988_ (.A(_13591_), .B(_02981_), .Y(_02982_));
NAND_g _23989_ (.A(_10907_), .B(_02982_), .Y(_02983_));
NAND_g _23990_ (.A(_13418_), .B(_02983_), .Y(_02984_));
AND_g _23991_ (.A(_10904_), .B(_02984_), .Y(_02985_));
NOT_g _23992_ (.A(_02985_), .Y(_02986_));
AND_g _23993_ (.A(_13562_), .B(_02879_), .Y(_02987_));
AND_g _23994_ (.A(_10974_), .B(_02879_), .Y(_02988_));
NAND_g _23995_ (.A(_02986_), .B(_02987_), .Y(_02989_));
NAND_g _23996_ (.A(_02966_), .B(_02989_), .Y(_02990_));
NAND_g _23997_ (.A(_11055_), .B(decoder_pseudo_trigger_q), .Y(_02991_));
AND_g _23998_ (.A(dbg_next), .B(_02991_), .Y(_02992_));
NAND_g _23999_ (.A(_02990_), .B(_02992_), .Y(_02993_));
NAND_g _24000_ (.A(_02964_), .B(_02993_), .Y(_00628_));
NAND_g _24001_ (.A(_11040_), .B(q_ascii_instr[9]), .Y(_02994_));
AND_g _24002_ (.A(_10918_), .B(_02576_), .Y(_02995_));
NOR_g _24003_ (.A(instr_bltu), .B(_02945_), .Y(_02996_));
AND_g _24004_ (.A(_02995_), .B(_02996_), .Y(_02997_));
NOR_g _24005_ (.A(instr_lbu), .B(_02997_), .Y(_02998_));
NOR_g _24006_ (.A(instr_lhu), .B(_02998_), .Y(_02999_));
NOT_g _24007_ (.A(_02999_), .Y(_03000_));
NAND_g _24008_ (.A(_13585_), .B(_03000_), .Y(_03001_));
NAND_g _24009_ (.A(_13588_), .B(_03001_), .Y(_03002_));
NAND_g _24010_ (.A(_13598_), .B(_03002_), .Y(_03003_));
AND_g _24011_ (.A(_13583_), .B(_13597_), .Y(_03004_));
NAND_g _24012_ (.A(_03003_), .B(_03004_), .Y(_03005_));
NAND_g _24013_ (.A(_02817_), .B(_03005_), .Y(_03006_));
NAND_g _24014_ (.A(_02936_), .B(_03006_), .Y(_03007_));
NAND_g _24015_ (.A(_02916_), .B(_03007_), .Y(_03008_));
NAND_g _24016_ (.A(_11056_), .B(decoder_pseudo_trigger_q), .Y(_03009_));
AND_g _24017_ (.A(dbg_next), .B(_03009_), .Y(_03010_));
NAND_g _24018_ (.A(_03008_), .B(_03010_), .Y(_03011_));
NAND_g _24019_ (.A(_02994_), .B(_03011_), .Y(_00629_));
NAND_g _24020_ (.A(_11040_), .B(q_ascii_instr[10]), .Y(_03012_));
AND_g _24021_ (.A(_13575_), .B(_02936_), .Y(_03013_));
AND_g _24022_ (.A(_10970_), .B(_13580_), .Y(_03014_));
AND_g _24023_ (.A(_10962_), .B(_02918_), .Y(_03015_));
NAND_g _24024_ (.A(_10962_), .B(_02918_), .Y(_03016_));
AND_g _24025_ (.A(_02856_), .B(_02995_), .Y(_03017_));
NAND_g _24026_ (.A(_03016_), .B(_03017_), .Y(_03018_));
AND_g _24027_ (.A(_13586_), .B(_02574_), .Y(_03019_));
NAND_g _24028_ (.A(_03018_), .B(_03019_), .Y(_03020_));
NAND_g _24029_ (.A(_13587_), .B(_03020_), .Y(_03021_));
NAND_g _24030_ (.A(_02831_), .B(_03021_), .Y(_03022_));
NAND_g _24031_ (.A(_03014_), .B(_03022_), .Y(_03023_));
NAND_g _24032_ (.A(_10971_), .B(_03023_), .Y(_03024_));
NAND_g _24033_ (.A(_13597_), .B(_03024_), .Y(_03025_));
NAND_g _24034_ (.A(_13418_), .B(_03025_), .Y(_03026_));
NAND_g _24035_ (.A(_03013_), .B(_03026_), .Y(_03027_));
NAND_g _24036_ (.A(_10975_), .B(_03027_), .Y(_03028_));
NAND_g _24037_ (.A(_11223_), .B(_03028_), .Y(_03029_));
NAND_g _24038_ (.A(_11057_), .B(decoder_pseudo_trigger_q), .Y(_03030_));
AND_g _24039_ (.A(dbg_next), .B(_03030_), .Y(_03031_));
NAND_g _24040_ (.A(_03029_), .B(_03031_), .Y(_03032_));
NAND_g _24041_ (.A(_03012_), .B(_03032_), .Y(_00630_));
NAND_g _24042_ (.A(_11040_), .B(q_ascii_instr[11]), .Y(_03033_));
NAND_g _24043_ (.A(_13570_), .B(_02822_), .Y(_03034_));
NAND_g _24044_ (.A(_13569_), .B(_03034_), .Y(_03035_));
AND_g _24045_ (.A(_02576_), .B(_03035_), .Y(_03036_));
NOR_g _24046_ (.A(instr_lbu), .B(_03036_), .Y(_03037_));
NOR_g _24047_ (.A(instr_lhu), .B(_03037_), .Y(_03038_));
NOT_g _24048_ (.A(_03038_), .Y(_03039_));
NAND_g _24049_ (.A(_13589_), .B(_03039_), .Y(_03040_));
NAND_g _24050_ (.A(_10915_), .B(_03040_), .Y(_03041_));
NAND_g _24051_ (.A(_02836_), .B(_03041_), .Y(_03042_));
NAND_g _24052_ (.A(_13581_), .B(_03042_), .Y(_03043_));
AND_g _24053_ (.A(_10971_), .B(_12522_), .Y(_03044_));
NAND_g _24054_ (.A(_03043_), .B(_03044_), .Y(_03045_));
NAND_g _24055_ (.A(_13590_), .B(_03045_), .Y(_03046_));
NAND_g _24056_ (.A(_10908_), .B(_03046_), .Y(_03047_));
AND_g _24057_ (.A(_10907_), .B(_03047_), .Y(_03048_));
NOT_g _24058_ (.A(_03048_), .Y(_03049_));
NAND_g _24059_ (.A(_13418_), .B(_03049_), .Y(_03050_));
AND_g _24060_ (.A(_10972_), .B(_13575_), .Y(_03051_));
NAND_g _24061_ (.A(_03050_), .B(_03051_), .Y(_03052_));
AND_g _24062_ (.A(_13564_), .B(_03052_), .Y(_03053_));
NAND_g _24063_ (.A(_13564_), .B(_03052_), .Y(_03054_));
NAND_g _24064_ (.A(_11223_), .B(_03054_), .Y(_03055_));
NAND_g _24065_ (.A(_11058_), .B(decoder_pseudo_trigger_q), .Y(_03056_));
AND_g _24066_ (.A(dbg_next), .B(_03056_), .Y(_03057_));
NAND_g _24067_ (.A(_03055_), .B(_03057_), .Y(_03058_));
NAND_g _24068_ (.A(_03033_), .B(_03058_), .Y(_00631_));
NAND_g _24069_ (.A(_11040_), .B(q_ascii_instr[12]), .Y(_03059_));
AND_g _24070_ (.A(_10916_), .B(_13598_), .Y(_03060_));
NAND_g _24071_ (.A(_02819_), .B(_02856_), .Y(_03061_));
NAND_g _24072_ (.A(_10919_), .B(_03061_), .Y(_03062_));
AND_g _24073_ (.A(_10918_), .B(_02577_), .Y(_03063_));
NAND_g _24074_ (.A(_03062_), .B(_03063_), .Y(_03064_));
NAND_g _24075_ (.A(_13585_), .B(_03064_), .Y(_03065_));
NAND_g _24076_ (.A(_10917_), .B(_03065_), .Y(_03066_));
NAND_g _24077_ (.A(_03060_), .B(_03066_), .Y(_03067_));
AND_g _24078_ (.A(instr_sltiu), .B(_13598_), .Y(_03068_));
NAND_g _24079_ (.A(instr_sltiu), .B(_13598_), .Y(_03069_));
AND_g _24080_ (.A(_12522_), .B(_13583_), .Y(_03070_));
AND_g _24081_ (.A(_03069_), .B(_03070_), .Y(_03071_));
NAND_g _24082_ (.A(_03067_), .B(_03071_), .Y(_03072_));
AND_g _24083_ (.A(_10910_), .B(_03072_), .Y(_03073_));
NOT_g _24084_ (.A(_03073_), .Y(_03074_));
NAND_g _24085_ (.A(_13590_), .B(_03074_), .Y(_03075_));
NAND_g _24086_ (.A(_10908_), .B(_03075_), .Y(_03076_));
AND_g _24087_ (.A(_10907_), .B(_03076_), .Y(_03077_));
NOT_g _24088_ (.A(_03077_), .Y(_03078_));
NAND_g _24089_ (.A(_13418_), .B(_03078_), .Y(_03079_));
NAND_g _24090_ (.A(_03013_), .B(_03079_), .Y(_03080_));
AND_g _24091_ (.A(_13562_), .B(_03080_), .Y(_03081_));
NAND_g _24092_ (.A(_11223_), .B(_03081_), .Y(_03082_));
NAND_g _24093_ (.A(_11059_), .B(decoder_pseudo_trigger_q), .Y(_03083_));
AND_g _24094_ (.A(dbg_next), .B(_03083_), .Y(_03084_));
NAND_g _24095_ (.A(_03082_), .B(_03084_), .Y(_03085_));
NAND_g _24096_ (.A(_03059_), .B(_03085_), .Y(_00632_));
NOR_g _24097_ (.A(dbg_next), .B(q_ascii_instr[14]), .Y(_03086_));
NAND_g _24098_ (.A(_11223_), .B(_13610_), .Y(_03087_));
NAND_g _24099_ (.A(cached_ascii_instr[14]), .B(decoder_pseudo_trigger_q), .Y(_03088_));
AND_g _24100_ (.A(dbg_next), .B(_03088_), .Y(_03089_));
AND_g _24101_ (.A(_03087_), .B(_03089_), .Y(_03090_));
NOR_g _24102_ (.A(_03086_), .B(_03090_), .Y(_00633_));
NAND_g _24103_ (.A(_11040_), .B(q_ascii_instr[16]), .Y(_03091_));
NAND_g _24104_ (.A(_10918_), .B(_02861_), .Y(_03092_));
NAND_g _24105_ (.A(_13585_), .B(_02577_), .Y(_03093_));
AND_g _24106_ (.A(_13589_), .B(_02577_), .Y(_03094_));
NAND_g _24107_ (.A(_03092_), .B(_03094_), .Y(_03095_));
NAND_g _24108_ (.A(_13598_), .B(_03095_), .Y(_03096_));
NAND_g _24109_ (.A(_13583_), .B(_03096_), .Y(_03097_));
NAND_g _24110_ (.A(_13596_), .B(_03097_), .Y(_03098_));
NAND_g _24111_ (.A(_13592_), .B(_03098_), .Y(_03099_));
NAND_g _24112_ (.A(_13418_), .B(_03099_), .Y(_03100_));
NAND_g _24113_ (.A(_10904_), .B(_03100_), .Y(_03101_));
NAND_g _24114_ (.A(_02988_), .B(_03101_), .Y(_03102_));
NAND_g _24115_ (.A(_02915_), .B(_03102_), .Y(_03103_));
NAND_g _24116_ (.A(_11223_), .B(_03103_), .Y(_03104_));
NAND_g _24117_ (.A(_11060_), .B(decoder_pseudo_trigger_q), .Y(_03105_));
AND_g _24118_ (.A(dbg_next), .B(_03105_), .Y(_03106_));
NAND_g _24119_ (.A(_03104_), .B(_03106_), .Y(_03107_));
NAND_g _24120_ (.A(_03091_), .B(_03107_), .Y(_00634_));
NAND_g _24121_ (.A(_11040_), .B(q_ascii_instr[17]), .Y(_03108_));
NAND_g _24122_ (.A(_02854_), .B(_02889_), .Y(_03109_));
NAND_g _24123_ (.A(_10919_), .B(_03109_), .Y(_03110_));
NAND_g _24124_ (.A(_10918_), .B(_03110_), .Y(_03111_));
NAND_g _24125_ (.A(_03094_), .B(_03111_), .Y(_03112_));
NAND_g _24126_ (.A(_02836_), .B(_03112_), .Y(_03113_));
AND_g _24127_ (.A(_10969_), .B(_03113_), .Y(_03114_));
NOT_g _24128_ (.A(_03114_), .Y(_03115_));
NAND_g _24129_ (.A(_13417_), .B(_03115_), .Y(_03116_));
NAND_g _24130_ (.A(_10911_), .B(_03116_), .Y(_03117_));
NAND_g _24131_ (.A(_13595_), .B(_03117_), .Y(_03118_));
NAND_g _24132_ (.A(_13592_), .B(_03118_), .Y(_03119_));
NAND_g _24133_ (.A(_13418_), .B(_03119_), .Y(_03120_));
AND_g _24134_ (.A(_02915_), .B(_03051_), .Y(_03121_));
NAND_g _24135_ (.A(_03120_), .B(_03121_), .Y(_03122_));
AND_g _24136_ (.A(_02915_), .B(_02935_), .Y(_03123_));
NOR_g _24137_ (.A(decoder_pseudo_trigger_q), .B(_03123_), .Y(_03124_));
NAND_g _24138_ (.A(_03122_), .B(_03124_), .Y(_03125_));
NAND_g _24139_ (.A(_11061_), .B(decoder_pseudo_trigger_q), .Y(_03126_));
AND_g _24140_ (.A(dbg_next), .B(_03126_), .Y(_03127_));
NAND_g _24141_ (.A(_03125_), .B(_03127_), .Y(_03128_));
NAND_g _24142_ (.A(_03108_), .B(_03128_), .Y(_00635_));
NAND_g _24143_ (.A(_11040_), .B(q_ascii_instr[18]), .Y(_03129_));
NAND_g _24144_ (.A(_02856_), .B(_03015_), .Y(_03130_));
NAND_g _24145_ (.A(_13568_), .B(_03130_), .Y(_03131_));
NAND_g _24146_ (.A(_02576_), .B(_03131_), .Y(_03132_));
NAND_g _24147_ (.A(_02574_), .B(_03132_), .Y(_03133_));
NAND_g _24148_ (.A(_13586_), .B(_03133_), .Y(_03134_));
NAND_g _24149_ (.A(_02834_), .B(_03134_), .Y(_03135_));
AND_g _24150_ (.A(_13417_), .B(_13596_), .Y(_03136_));
NAND_g _24151_ (.A(_03135_), .B(_03136_), .Y(_03137_));
NAND_g _24152_ (.A(_10908_), .B(_03137_), .Y(_03138_));
AND_g _24153_ (.A(_13563_), .B(_02817_), .Y(_03139_));
AND_g _24154_ (.A(_02817_), .B(_03138_), .Y(_03140_));
NAND_g _24155_ (.A(_02936_), .B(_03140_), .Y(_03141_));
NAND_g _24156_ (.A(_02917_), .B(_03141_), .Y(_03142_));
NAND_g _24157_ (.A(_11062_), .B(decoder_pseudo_trigger_q), .Y(_03143_));
AND_g _24158_ (.A(dbg_next), .B(_03143_), .Y(_03144_));
NAND_g _24159_ (.A(_03142_), .B(_03144_), .Y(_03145_));
NAND_g _24160_ (.A(_03129_), .B(_03145_), .Y(_00636_));
NAND_g _24161_ (.A(_11040_), .B(q_ascii_instr[19]), .Y(_03146_));
NAND_g _24162_ (.A(_00006_), .B(_03017_), .Y(_03147_));
NAND_g _24163_ (.A(instr_bltu), .B(_02995_), .Y(_03148_));
AND_g _24164_ (.A(_02574_), .B(_03148_), .Y(_03149_));
NAND_g _24165_ (.A(_03147_), .B(_03149_), .Y(_03150_));
NAND_g _24166_ (.A(_13586_), .B(_03150_), .Y(_03151_));
NAND_g _24167_ (.A(_03060_), .B(_03151_), .Y(_03152_));
NAND_g _24168_ (.A(_03069_), .B(_03152_), .Y(_03153_));
NAND_g _24169_ (.A(_13580_), .B(_03153_), .Y(_03154_));
NAND_g _24170_ (.A(_03136_), .B(_03154_), .Y(_03155_));
NAND_g _24171_ (.A(_13592_), .B(_03155_), .Y(_03156_));
AND_g _24172_ (.A(_13418_), .B(_03051_), .Y(_03157_));
NAND_g _24173_ (.A(_13418_), .B(_03051_), .Y(_03158_));
AND_g _24174_ (.A(_13562_), .B(_03157_), .Y(_03159_));
NAND_g _24175_ (.A(_03156_), .B(_03159_), .Y(_03160_));
NAND_g _24176_ (.A(_02966_), .B(_03160_), .Y(_03161_));
NAND_g _24177_ (.A(_11063_), .B(decoder_pseudo_trigger_q), .Y(_03162_));
AND_g _24178_ (.A(dbg_next), .B(_03162_), .Y(_03163_));
NAND_g _24179_ (.A(_03161_), .B(_03163_), .Y(_03164_));
NAND_g _24180_ (.A(_03146_), .B(_03164_), .Y(_00637_));
NAND_g _24181_ (.A(_11040_), .B(q_ascii_instr[20]), .Y(_03165_));
NAND_g _24182_ (.A(_03014_), .B(_03068_), .Y(_03166_));
NAND_g _24183_ (.A(_13417_), .B(_03166_), .Y(_03167_));
NAND_g _24184_ (.A(_10911_), .B(_03167_), .Y(_03168_));
NAND_g _24185_ (.A(_13595_), .B(_03168_), .Y(_03169_));
AND_g _24186_ (.A(_10908_), .B(_03169_), .Y(_03170_));
NOT_g _24187_ (.A(_03170_), .Y(_03171_));
NAND_g _24188_ (.A(_02816_), .B(_03171_), .Y(_03172_));
NAND_g _24189_ (.A(_03013_), .B(_03172_), .Y(_03173_));
AND_g _24190_ (.A(_13562_), .B(_03173_), .Y(_03174_));
NAND_g _24191_ (.A(_11223_), .B(_03174_), .Y(_03175_));
NAND_g _24192_ (.A(_11064_), .B(decoder_pseudo_trigger_q), .Y(_03176_));
AND_g _24193_ (.A(dbg_next), .B(_03176_), .Y(_03177_));
NAND_g _24194_ (.A(_03175_), .B(_03177_), .Y(_03178_));
NAND_g _24195_ (.A(_03165_), .B(_03178_), .Y(_00638_));
NAND_g _24196_ (.A(_11040_), .B(q_ascii_instr[22]), .Y(_03179_));
NAND_g _24197_ (.A(_13574_), .B(_02576_), .Y(_03180_));
NAND_g _24198_ (.A(_02574_), .B(_03180_), .Y(_03181_));
NAND_g _24199_ (.A(_13586_), .B(_03181_), .Y(_03182_));
AND_g _24200_ (.A(_13418_), .B(_13594_), .Y(_03183_));
AND_g _24201_ (.A(_02869_), .B(_03183_), .Y(_03184_));
NAND_g _24202_ (.A(_03182_), .B(_03184_), .Y(_03185_));
NAND_g _24203_ (.A(_13575_), .B(_03185_), .Y(_03186_));
AND_g _24204_ (.A(_10903_), .B(_13565_), .Y(_03187_));
AND_g _24205_ (.A(_03186_), .B(_03187_), .Y(_03188_));
NAND_g _24206_ (.A(_11223_), .B(_03188_), .Y(_03189_));
NAND_g _24207_ (.A(_11065_), .B(decoder_pseudo_trigger_q), .Y(_03190_));
AND_g _24208_ (.A(dbg_next), .B(_03190_), .Y(_03191_));
NAND_g _24209_ (.A(_03189_), .B(_03191_), .Y(_03192_));
NAND_g _24210_ (.A(_03179_), .B(_03192_), .Y(_00639_));
NAND_g _24211_ (.A(_11040_), .B(q_ascii_instr[24]), .Y(_03193_));
AND_g _24212_ (.A(_02995_), .B(_03019_), .Y(_03194_));
NAND_g _24213_ (.A(_02858_), .B(_03194_), .Y(_03195_));
NAND_g _24214_ (.A(_13587_), .B(_03195_), .Y(_03196_));
NAND_g _24215_ (.A(_02831_), .B(_03196_), .Y(_03197_));
NAND_g _24216_ (.A(_13583_), .B(_03197_), .Y(_03198_));
NAND_g _24217_ (.A(_13596_), .B(_03198_), .Y(_03199_));
NAND_g _24218_ (.A(_10908_), .B(_03199_), .Y(_03200_));
NAND_g _24219_ (.A(_02817_), .B(_03200_), .Y(_03201_));
NAND_g _24220_ (.A(_13563_), .B(_03201_), .Y(_03202_));
NAND_g _24221_ (.A(_10974_), .B(_03202_), .Y(_03203_));
NAND_g _24222_ (.A(_02916_), .B(_03203_), .Y(_03204_));
NAND_g _24223_ (.A(_11066_), .B(decoder_pseudo_trigger_q), .Y(_03205_));
AND_g _24224_ (.A(dbg_next), .B(_03205_), .Y(_03206_));
NAND_g _24225_ (.A(_03204_), .B(_03206_), .Y(_03207_));
NAND_g _24226_ (.A(_03193_), .B(_03207_), .Y(_00640_));
NAND_g _24227_ (.A(_11040_), .B(q_ascii_instr[25]), .Y(_03208_));
AND_g _24228_ (.A(_11223_), .B(_13564_), .Y(_03209_));
NAND_g _24229_ (.A(_11223_), .B(_13564_), .Y(_03210_));
NAND_g _24230_ (.A(_13568_), .B(_02859_), .Y(_03211_));
AND_g _24231_ (.A(_13586_), .B(_02577_), .Y(_03212_));
NAND_g _24232_ (.A(_03211_), .B(_03212_), .Y(_03213_));
NAND_g _24233_ (.A(_10916_), .B(_03213_), .Y(_03214_));
NAND_g _24234_ (.A(_02832_), .B(_03214_), .Y(_03215_));
NAND_g _24235_ (.A(_13582_), .B(_03215_), .Y(_03216_));
NAND_g _24236_ (.A(_13596_), .B(_03216_), .Y(_03217_));
NAND_g _24237_ (.A(_10908_), .B(_03217_), .Y(_03218_));
NAND_g _24238_ (.A(_03139_), .B(_03218_), .Y(_03219_));
NAND_g _24239_ (.A(_03209_), .B(_03219_), .Y(_03220_));
NAND_g _24240_ (.A(_11067_), .B(decoder_pseudo_trigger_q), .Y(_03221_));
AND_g _24241_ (.A(dbg_next), .B(_03221_), .Y(_03222_));
NAND_g _24242_ (.A(_03220_), .B(_03222_), .Y(_03223_));
NAND_g _24243_ (.A(_03208_), .B(_03223_), .Y(_00641_));
NAND_g _24244_ (.A(_11040_), .B(q_ascii_instr[26]), .Y(_03224_));
NOR_g _24245_ (.A(instr_slti), .B(_03195_), .Y(_03225_));
NOR_g _24246_ (.A(instr_sltiu), .B(_03225_), .Y(_03226_));
AND_g _24247_ (.A(_13597_), .B(_02837_), .Y(_03227_));
NOR_g _24248_ (.A(_03158_), .B(_03226_), .Y(_03228_));
NAND_g _24249_ (.A(_03227_), .B(_03228_), .Y(_03229_));
NAND_g _24250_ (.A(_10974_), .B(_03229_), .Y(_03230_));
NAND_g _24251_ (.A(_02915_), .B(_03230_), .Y(_03231_));
NAND_g _24252_ (.A(_11223_), .B(_03231_), .Y(_03232_));
NAND_g _24253_ (.A(_11068_), .B(decoder_pseudo_trigger_q), .Y(_03233_));
AND_g _24254_ (.A(dbg_next), .B(_03233_), .Y(_03234_));
NAND_g _24255_ (.A(_03232_), .B(_03234_), .Y(_03235_));
NAND_g _24256_ (.A(_03224_), .B(_03235_), .Y(_00642_));
NAND_g _24257_ (.A(_11040_), .B(q_ascii_instr[27]), .Y(_03236_));
AND_g _24258_ (.A(_13589_), .B(_02860_), .Y(_03237_));
NAND_g _24259_ (.A(_03063_), .B(_03237_), .Y(_03238_));
NAND_g _24260_ (.A(_02830_), .B(_03238_), .Y(_03239_));
AND_g _24261_ (.A(_13594_), .B(_03044_), .Y(_03240_));
AND_g _24262_ (.A(_02915_), .B(_03014_), .Y(_03241_));
AND_g _24263_ (.A(_13577_), .B(_03241_), .Y(_03242_));
AND_g _24264_ (.A(_03240_), .B(_03242_), .Y(_03243_));
NAND_g _24265_ (.A(_03239_), .B(_03243_), .Y(_03244_));
NAND_g _24266_ (.A(_03124_), .B(_03244_), .Y(_03245_));
NAND_g _24267_ (.A(_11069_), .B(decoder_pseudo_trigger_q), .Y(_03246_));
AND_g _24268_ (.A(dbg_next), .B(_03246_), .Y(_03247_));
NAND_g _24269_ (.A(_03245_), .B(_03247_), .Y(_03248_));
NAND_g _24270_ (.A(_03236_), .B(_03248_), .Y(_00643_));
NAND_g _24271_ (.A(_11040_), .B(q_ascii_instr[28]), .Y(_03249_));
NAND_g _24272_ (.A(_10916_), .B(_03195_), .Y(_03250_));
NAND_g _24273_ (.A(_10915_), .B(_03250_), .Y(_03251_));
AND_g _24274_ (.A(_10914_), .B(_03251_), .Y(_03252_));
NOT_g _24275_ (.A(_03252_), .Y(_03253_));
NAND_g _24276_ (.A(_02829_), .B(_03253_), .Y(_03254_));
NAND_g _24277_ (.A(_13582_), .B(_03254_), .Y(_03255_));
NAND_g _24278_ (.A(_13596_), .B(_03255_), .Y(_03256_));
NAND_g _24279_ (.A(_10908_), .B(_03256_), .Y(_03257_));
NAND_g _24280_ (.A(_02817_), .B(_03257_), .Y(_03258_));
AND_g _24281_ (.A(_10972_), .B(_03258_), .Y(_03259_));
NOT_g _24282_ (.A(_03259_), .Y(_03260_));
NAND_g _24283_ (.A(_13564_), .B(_03260_), .Y(_03261_));
NAND_g _24284_ (.A(_02916_), .B(_03261_), .Y(_03262_));
NAND_g _24285_ (.A(_11070_), .B(decoder_pseudo_trigger_q), .Y(_03263_));
AND_g _24286_ (.A(dbg_next), .B(_03263_), .Y(_03264_));
NAND_g _24287_ (.A(_03262_), .B(_03264_), .Y(_03265_));
NAND_g _24288_ (.A(_03249_), .B(_03265_), .Y(_00644_));
NAND_g _24289_ (.A(_11040_), .B(q_ascii_instr[30]), .Y(_03266_));
NOR_g _24290_ (.A(_02858_), .B(_03211_), .Y(_03267_));
NOR_g _24291_ (.A(_03093_), .B(_03267_), .Y(_03268_));
NOR_g _24292_ (.A(_02833_), .B(_03268_), .Y(_03269_));
NOR_g _24293_ (.A(instr_ori), .B(_03269_), .Y(_03270_));
NOT_g _24294_ (.A(_03270_), .Y(_03271_));
NAND_g _24295_ (.A(_13583_), .B(_03271_), .Y(_03272_));
NAND_g _24296_ (.A(_13596_), .B(_03272_), .Y(_03273_));
NAND_g _24297_ (.A(_10908_), .B(_03273_), .Y(_03274_));
NAND_g _24298_ (.A(_02817_), .B(_03274_), .Y(_03275_));
AND_g _24299_ (.A(_13565_), .B(_03275_), .Y(_03276_));
NAND_g _24300_ (.A(_11223_), .B(_03276_), .Y(_03277_));
NAND_g _24301_ (.A(_11071_), .B(decoder_pseudo_trigger_q), .Y(_03278_));
AND_g _24302_ (.A(dbg_next), .B(_03278_), .Y(_03279_));
NAND_g _24303_ (.A(_03277_), .B(_03279_), .Y(_03280_));
NAND_g _24304_ (.A(_03266_), .B(_03280_), .Y(_00645_));
NAND_g _24305_ (.A(_11040_), .B(q_ascii_instr[32]), .Y(_03281_));
AND_g _24306_ (.A(_02936_), .B(_03229_), .Y(_03282_));
NOT_g _24307_ (.A(_03282_), .Y(_03283_));
NOR_g _24308_ (.A(instr_rdinstrh), .B(_03282_), .Y(_03284_));
NOR_g _24309_ (.A(decoder_pseudo_trigger_q), .B(_03284_), .Y(_03285_));
NOT_g _24310_ (.A(_03285_), .Y(_03286_));
NAND_g _24311_ (.A(_11072_), .B(decoder_pseudo_trigger_q), .Y(_03287_));
AND_g _24312_ (.A(dbg_next), .B(_03287_), .Y(_03288_));
NAND_g _24313_ (.A(_03286_), .B(_03288_), .Y(_03289_));
NAND_g _24314_ (.A(_03281_), .B(_03289_), .Y(_00646_));
NAND_g _24315_ (.A(_11040_), .B(q_ascii_instr[33]), .Y(_03290_));
NOR_g _24316_ (.A(_03158_), .B(_03166_), .Y(_03291_));
AND_g _24317_ (.A(_03240_), .B(_03291_), .Y(_03292_));
NAND_g _24318_ (.A(_03240_), .B(_03291_), .Y(_03293_));
NAND_g _24319_ (.A(_10972_), .B(_03293_), .Y(_03294_));
NAND_g _24320_ (.A(_13564_), .B(_03294_), .Y(_03295_));
NAND_g _24321_ (.A(_02916_), .B(_03295_), .Y(_03296_));
NAND_g _24322_ (.A(_11073_), .B(decoder_pseudo_trigger_q), .Y(_03297_));
AND_g _24323_ (.A(dbg_next), .B(_03297_), .Y(_03298_));
NAND_g _24324_ (.A(_03296_), .B(_03298_), .Y(_03299_));
NAND_g _24325_ (.A(_03290_), .B(_03299_), .Y(_00647_));
NAND_g _24326_ (.A(_11074_), .B(decoder_pseudo_trigger_q), .Y(_03300_));
NAND_g _24327_ (.A(_11040_), .B(q_ascii_instr[35]), .Y(_03301_));
AND_g _24328_ (.A(dbg_next), .B(_03300_), .Y(_03302_));
NAND_g _24329_ (.A(_03210_), .B(_03302_), .Y(_03303_));
NAND_g _24330_ (.A(_03301_), .B(_03303_), .Y(_00648_));
NAND_g _24331_ (.A(_11040_), .B(q_ascii_instr[36]), .Y(_03304_));
NAND_g _24332_ (.A(_13562_), .B(_03292_), .Y(_03305_));
NAND_g _24333_ (.A(_02966_), .B(_03305_), .Y(_03306_));
NAND_g _24334_ (.A(_11075_), .B(decoder_pseudo_trigger_q), .Y(_03307_));
AND_g _24335_ (.A(dbg_next), .B(_03307_), .Y(_03308_));
NAND_g _24336_ (.A(_03306_), .B(_03308_), .Y(_03309_));
NAND_g _24337_ (.A(_03304_), .B(_03309_), .Y(_00649_));
NAND_g _24338_ (.A(_11040_), .B(q_ascii_instr[38]), .Y(_03310_));
NAND_g _24339_ (.A(_02916_), .B(_03282_), .Y(_03311_));
NAND_g _24340_ (.A(_11076_), .B(decoder_pseudo_trigger_q), .Y(_03312_));
AND_g _24341_ (.A(dbg_next), .B(_03312_), .Y(_03313_));
NAND_g _24342_ (.A(_03311_), .B(_03313_), .Y(_03314_));
NAND_g _24343_ (.A(_03310_), .B(_03314_), .Y(_00650_));
NOR_g _24344_ (.A(cached_ascii_instr[41]), .B(_11223_), .Y(_03315_));
NOR_g _24345_ (.A(_02966_), .B(_03315_), .Y(_03316_));
NOR_g _24346_ (.A(_11040_), .B(_03316_), .Y(_03317_));
NOR_g _24347_ (.A(dbg_next), .B(q_ascii_instr[41]), .Y(_03318_));
NOR_g _24348_ (.A(_03317_), .B(_03318_), .Y(_00651_));
NOR_g _24349_ (.A(cached_ascii_instr[43]), .B(_11223_), .Y(_03319_));
NOR_g _24350_ (.A(_02916_), .B(_03319_), .Y(_03320_));
NAND_g _24351_ (.A(_11040_), .B(q_ascii_instr[43]), .Y(_03321_));
NAND_g _24352_ (.A(dbg_next), .B(_03320_), .Y(_03322_));
NAND_g _24353_ (.A(_03321_), .B(_03322_), .Y(_00652_));
NOR_g _24354_ (.A(cached_ascii_instr[52]), .B(_11223_), .Y(_03323_));
NOR_g _24355_ (.A(_03124_), .B(_03323_), .Y(_03324_));
NOR_g _24356_ (.A(_11040_), .B(_03324_), .Y(_03325_));
NOR_g _24357_ (.A(dbg_next), .B(q_ascii_instr[52]), .Y(_03326_));
NOR_g _24358_ (.A(_03325_), .B(_03326_), .Y(_00653_));
NAND_g _24359_ (.A(cached_ascii_instr[54]), .B(decoder_pseudo_trigger_q), .Y(_03327_));
NAND_g _24360_ (.A(_11223_), .B(_13566_), .Y(_03328_));
NOR_g _24361_ (.A(dbg_next), .B(q_ascii_instr[54]), .Y(_03329_));
AND_g _24362_ (.A(dbg_next), .B(_03327_), .Y(_03330_));
AND_g _24363_ (.A(_03328_), .B(_03330_), .Y(_03331_));
NOR_g _24364_ (.A(_03329_), .B(_03331_), .Y(_00654_));
NOR_g _24365_ (.A(cached_ascii_instr[62]), .B(_11223_), .Y(_03332_));
NOR_g _24366_ (.A(_02917_), .B(_03332_), .Y(_03333_));
NOR_g _24367_ (.A(_11040_), .B(_03333_), .Y(_03334_));
NOR_g _24368_ (.A(dbg_next), .B(q_ascii_instr[62]), .Y(_03335_));
NOR_g _24369_ (.A(_03334_), .B(_03335_), .Y(_00655_));
NAND_g _24370_ (.A(decoded_imm[0]), .B(_11223_), .Y(_03336_));
NAND_g _24371_ (.A(cached_insn_imm[0]), .B(decoder_pseudo_trigger_q), .Y(_03337_));
NOR_g _24372_ (.A(dbg_next), .B(q_insn_imm[0]), .Y(_03338_));
AND_g _24373_ (.A(dbg_next), .B(_03337_), .Y(_03339_));
AND_g _24374_ (.A(_03336_), .B(_03339_), .Y(_03340_));
NOR_g _24375_ (.A(_03338_), .B(_03340_), .Y(_00656_));
NAND_g _24376_ (.A(decoded_imm[1]), .B(_11223_), .Y(_03341_));
NAND_g _24377_ (.A(cached_insn_imm[1]), .B(decoder_pseudo_trigger_q), .Y(_03342_));
NOR_g _24378_ (.A(dbg_next), .B(q_insn_imm[1]), .Y(_03343_));
AND_g _24379_ (.A(dbg_next), .B(_03342_), .Y(_03344_));
AND_g _24380_ (.A(_03341_), .B(_03344_), .Y(_03345_));
NOR_g _24381_ (.A(_03343_), .B(_03345_), .Y(_00657_));
NAND_g _24382_ (.A(decoded_imm[2]), .B(_11223_), .Y(_03346_));
NAND_g _24383_ (.A(cached_insn_imm[2]), .B(decoder_pseudo_trigger_q), .Y(_03347_));
NOR_g _24384_ (.A(dbg_next), .B(q_insn_imm[2]), .Y(_03348_));
AND_g _24385_ (.A(dbg_next), .B(_03347_), .Y(_03349_));
AND_g _24386_ (.A(_03346_), .B(_03349_), .Y(_03350_));
NOR_g _24387_ (.A(_03348_), .B(_03350_), .Y(_00658_));
NAND_g _24388_ (.A(decoded_imm[3]), .B(_11223_), .Y(_03351_));
NAND_g _24389_ (.A(cached_insn_imm[3]), .B(decoder_pseudo_trigger_q), .Y(_03352_));
NOR_g _24390_ (.A(dbg_next), .B(q_insn_imm[3]), .Y(_03353_));
AND_g _24391_ (.A(dbg_next), .B(_03352_), .Y(_03354_));
AND_g _24392_ (.A(_03351_), .B(_03354_), .Y(_03355_));
NOR_g _24393_ (.A(_03353_), .B(_03355_), .Y(_00659_));
NAND_g _24394_ (.A(decoded_imm[4]), .B(_11223_), .Y(_03356_));
NAND_g _24395_ (.A(cached_insn_imm[4]), .B(decoder_pseudo_trigger_q), .Y(_03357_));
NOR_g _24396_ (.A(dbg_next), .B(q_insn_imm[4]), .Y(_03358_));
AND_g _24397_ (.A(dbg_next), .B(_03357_), .Y(_03359_));
AND_g _24398_ (.A(_03356_), .B(_03359_), .Y(_03360_));
NOR_g _24399_ (.A(_03358_), .B(_03360_), .Y(_00660_));
NAND_g _24400_ (.A(decoded_imm[5]), .B(_11223_), .Y(_03361_));
NAND_g _24401_ (.A(cached_insn_imm[5]), .B(decoder_pseudo_trigger_q), .Y(_03362_));
NOR_g _24402_ (.A(dbg_next), .B(q_insn_imm[5]), .Y(_03363_));
AND_g _24403_ (.A(dbg_next), .B(_03362_), .Y(_03364_));
AND_g _24404_ (.A(_03361_), .B(_03364_), .Y(_03365_));
NOR_g _24405_ (.A(_03363_), .B(_03365_), .Y(_00661_));
NAND_g _24406_ (.A(decoded_imm[6]), .B(_11223_), .Y(_03366_));
NAND_g _24407_ (.A(cached_insn_imm[6]), .B(decoder_pseudo_trigger_q), .Y(_03367_));
NOR_g _24408_ (.A(dbg_next), .B(q_insn_imm[6]), .Y(_03368_));
AND_g _24409_ (.A(dbg_next), .B(_03367_), .Y(_03369_));
AND_g _24410_ (.A(_03366_), .B(_03369_), .Y(_03370_));
NOR_g _24411_ (.A(_03368_), .B(_03370_), .Y(_00662_));
NAND_g _24412_ (.A(decoded_imm[7]), .B(_11223_), .Y(_03371_));
NAND_g _24413_ (.A(cached_insn_imm[7]), .B(decoder_pseudo_trigger_q), .Y(_03372_));
NOR_g _24414_ (.A(dbg_next), .B(q_insn_imm[7]), .Y(_03373_));
AND_g _24415_ (.A(dbg_next), .B(_03372_), .Y(_03374_));
AND_g _24416_ (.A(_03371_), .B(_03374_), .Y(_03375_));
NOR_g _24417_ (.A(_03373_), .B(_03375_), .Y(_00663_));
NAND_g _24418_ (.A(decoded_imm[8]), .B(_11223_), .Y(_03376_));
NAND_g _24419_ (.A(cached_insn_imm[8]), .B(decoder_pseudo_trigger_q), .Y(_03377_));
NOR_g _24420_ (.A(dbg_next), .B(q_insn_imm[8]), .Y(_03378_));
AND_g _24421_ (.A(dbg_next), .B(_03377_), .Y(_03379_));
AND_g _24422_ (.A(_03376_), .B(_03379_), .Y(_03380_));
NOR_g _24423_ (.A(_03378_), .B(_03380_), .Y(_00664_));
NAND_g _24424_ (.A(decoded_imm[9]), .B(_11223_), .Y(_03381_));
NAND_g _24425_ (.A(cached_insn_imm[9]), .B(decoder_pseudo_trigger_q), .Y(_03382_));
NOR_g _24426_ (.A(dbg_next), .B(q_insn_imm[9]), .Y(_03383_));
AND_g _24427_ (.A(dbg_next), .B(_03382_), .Y(_03384_));
AND_g _24428_ (.A(_03381_), .B(_03384_), .Y(_03385_));
NOR_g _24429_ (.A(_03383_), .B(_03385_), .Y(_00665_));
NAND_g _24430_ (.A(decoded_imm[10]), .B(_11223_), .Y(_03386_));
NAND_g _24431_ (.A(cached_insn_imm[10]), .B(decoder_pseudo_trigger_q), .Y(_03387_));
NOR_g _24432_ (.A(dbg_next), .B(q_insn_imm[10]), .Y(_03388_));
AND_g _24433_ (.A(dbg_next), .B(_03387_), .Y(_03389_));
AND_g _24434_ (.A(_03386_), .B(_03389_), .Y(_03390_));
NOR_g _24435_ (.A(_03388_), .B(_03390_), .Y(_00666_));
NAND_g _24436_ (.A(decoded_imm[11]), .B(_11223_), .Y(_03391_));
NAND_g _24437_ (.A(cached_insn_imm[11]), .B(decoder_pseudo_trigger_q), .Y(_03392_));
NOR_g _24438_ (.A(dbg_next), .B(q_insn_imm[11]), .Y(_03393_));
AND_g _24439_ (.A(dbg_next), .B(_03392_), .Y(_03394_));
AND_g _24440_ (.A(_03391_), .B(_03394_), .Y(_03395_));
NOR_g _24441_ (.A(_03393_), .B(_03395_), .Y(_00667_));
NAND_g _24442_ (.A(decoded_imm[12]), .B(_11223_), .Y(_03396_));
NAND_g _24443_ (.A(cached_insn_imm[12]), .B(decoder_pseudo_trigger_q), .Y(_03397_));
NOR_g _24444_ (.A(dbg_next), .B(q_insn_imm[12]), .Y(_03398_));
AND_g _24445_ (.A(dbg_next), .B(_03397_), .Y(_03399_));
AND_g _24446_ (.A(_03396_), .B(_03399_), .Y(_03400_));
NOR_g _24447_ (.A(_03398_), .B(_03400_), .Y(_00668_));
NAND_g _24448_ (.A(decoded_imm[13]), .B(_11223_), .Y(_03401_));
NAND_g _24449_ (.A(cached_insn_imm[13]), .B(decoder_pseudo_trigger_q), .Y(_03402_));
NOR_g _24450_ (.A(dbg_next), .B(q_insn_imm[13]), .Y(_03403_));
AND_g _24451_ (.A(dbg_next), .B(_03402_), .Y(_03404_));
AND_g _24452_ (.A(_03401_), .B(_03404_), .Y(_03405_));
NOR_g _24453_ (.A(_03403_), .B(_03405_), .Y(_00669_));
NAND_g _24454_ (.A(decoded_imm[14]), .B(_11223_), .Y(_03406_));
NAND_g _24455_ (.A(cached_insn_imm[14]), .B(decoder_pseudo_trigger_q), .Y(_03407_));
NOR_g _24456_ (.A(dbg_next), .B(q_insn_imm[14]), .Y(_03408_));
AND_g _24457_ (.A(dbg_next), .B(_03407_), .Y(_03409_));
AND_g _24458_ (.A(_03406_), .B(_03409_), .Y(_03410_));
NOR_g _24459_ (.A(_03408_), .B(_03410_), .Y(_00670_));
NAND_g _24460_ (.A(decoded_imm[15]), .B(_11223_), .Y(_03411_));
NAND_g _24461_ (.A(cached_insn_imm[15]), .B(decoder_pseudo_trigger_q), .Y(_03412_));
NOR_g _24462_ (.A(dbg_next), .B(q_insn_imm[15]), .Y(_03413_));
AND_g _24463_ (.A(dbg_next), .B(_03412_), .Y(_03414_));
AND_g _24464_ (.A(_03411_), .B(_03414_), .Y(_03415_));
NOR_g _24465_ (.A(_03413_), .B(_03415_), .Y(_00671_));
NAND_g _24466_ (.A(decoded_imm[16]), .B(_11223_), .Y(_03416_));
NAND_g _24467_ (.A(cached_insn_imm[16]), .B(decoder_pseudo_trigger_q), .Y(_03417_));
NOR_g _24468_ (.A(dbg_next), .B(q_insn_imm[16]), .Y(_03418_));
AND_g _24469_ (.A(dbg_next), .B(_03417_), .Y(_03419_));
AND_g _24470_ (.A(_03416_), .B(_03419_), .Y(_03420_));
NOR_g _24471_ (.A(_03418_), .B(_03420_), .Y(_00672_));
NAND_g _24472_ (.A(decoded_imm[17]), .B(_11223_), .Y(_03421_));
NAND_g _24473_ (.A(cached_insn_imm[17]), .B(decoder_pseudo_trigger_q), .Y(_03422_));
NOR_g _24474_ (.A(dbg_next), .B(q_insn_imm[17]), .Y(_03423_));
AND_g _24475_ (.A(dbg_next), .B(_03422_), .Y(_03424_));
AND_g _24476_ (.A(_03421_), .B(_03424_), .Y(_03425_));
NOR_g _24477_ (.A(_03423_), .B(_03425_), .Y(_00673_));
NAND_g _24478_ (.A(decoded_imm[18]), .B(_11223_), .Y(_03426_));
NAND_g _24479_ (.A(cached_insn_imm[18]), .B(decoder_pseudo_trigger_q), .Y(_03427_));
NOR_g _24480_ (.A(dbg_next), .B(q_insn_imm[18]), .Y(_03428_));
AND_g _24481_ (.A(dbg_next), .B(_03427_), .Y(_03429_));
AND_g _24482_ (.A(_03426_), .B(_03429_), .Y(_03430_));
NOR_g _24483_ (.A(_03428_), .B(_03430_), .Y(_00674_));
NAND_g _24484_ (.A(decoded_imm[19]), .B(_11223_), .Y(_03431_));
NAND_g _24485_ (.A(cached_insn_imm[19]), .B(decoder_pseudo_trigger_q), .Y(_03432_));
NOR_g _24486_ (.A(dbg_next), .B(q_insn_imm[19]), .Y(_03433_));
AND_g _24487_ (.A(dbg_next), .B(_03432_), .Y(_03434_));
AND_g _24488_ (.A(_03431_), .B(_03434_), .Y(_03435_));
NOR_g _24489_ (.A(_03433_), .B(_03435_), .Y(_00675_));
NAND_g _24490_ (.A(decoded_imm[20]), .B(_11223_), .Y(_03436_));
NAND_g _24491_ (.A(cached_insn_imm[20]), .B(decoder_pseudo_trigger_q), .Y(_03437_));
NOR_g _24492_ (.A(dbg_next), .B(q_insn_imm[20]), .Y(_03438_));
AND_g _24493_ (.A(dbg_next), .B(_03437_), .Y(_03439_));
AND_g _24494_ (.A(_03436_), .B(_03439_), .Y(_03440_));
NOR_g _24495_ (.A(_03438_), .B(_03440_), .Y(_00676_));
NAND_g _24496_ (.A(decoded_imm[21]), .B(_11223_), .Y(_03441_));
NAND_g _24497_ (.A(cached_insn_imm[21]), .B(decoder_pseudo_trigger_q), .Y(_03442_));
NOR_g _24498_ (.A(dbg_next), .B(q_insn_imm[21]), .Y(_03443_));
AND_g _24499_ (.A(dbg_next), .B(_03442_), .Y(_03444_));
AND_g _24500_ (.A(_03441_), .B(_03444_), .Y(_03445_));
NOR_g _24501_ (.A(_03443_), .B(_03445_), .Y(_00677_));
NAND_g _24502_ (.A(decoded_imm[22]), .B(_11223_), .Y(_03446_));
NAND_g _24503_ (.A(cached_insn_imm[22]), .B(decoder_pseudo_trigger_q), .Y(_03447_));
NOR_g _24504_ (.A(dbg_next), .B(q_insn_imm[22]), .Y(_03448_));
AND_g _24505_ (.A(dbg_next), .B(_03447_), .Y(_03449_));
AND_g _24506_ (.A(_03446_), .B(_03449_), .Y(_03450_));
NOR_g _24507_ (.A(_03448_), .B(_03450_), .Y(_00678_));
NAND_g _24508_ (.A(decoded_imm[23]), .B(_11223_), .Y(_03451_));
NAND_g _24509_ (.A(cached_insn_imm[23]), .B(decoder_pseudo_trigger_q), .Y(_03452_));
NOR_g _24510_ (.A(dbg_next), .B(q_insn_imm[23]), .Y(_03453_));
AND_g _24511_ (.A(dbg_next), .B(_03452_), .Y(_03454_));
AND_g _24512_ (.A(_03451_), .B(_03454_), .Y(_03455_));
NOR_g _24513_ (.A(_03453_), .B(_03455_), .Y(_00679_));
NAND_g _24514_ (.A(decoded_imm[24]), .B(_11223_), .Y(_03456_));
NAND_g _24515_ (.A(cached_insn_imm[24]), .B(decoder_pseudo_trigger_q), .Y(_03457_));
NOR_g _24516_ (.A(dbg_next), .B(q_insn_imm[24]), .Y(_03458_));
AND_g _24517_ (.A(dbg_next), .B(_03457_), .Y(_03459_));
AND_g _24518_ (.A(_03456_), .B(_03459_), .Y(_03460_));
NOR_g _24519_ (.A(_03458_), .B(_03460_), .Y(_00680_));
NAND_g _24520_ (.A(decoded_imm[25]), .B(_11223_), .Y(_03461_));
NAND_g _24521_ (.A(cached_insn_imm[25]), .B(decoder_pseudo_trigger_q), .Y(_03462_));
NOR_g _24522_ (.A(dbg_next), .B(q_insn_imm[25]), .Y(_03463_));
AND_g _24523_ (.A(dbg_next), .B(_03462_), .Y(_03464_));
AND_g _24524_ (.A(_03461_), .B(_03464_), .Y(_03465_));
NOR_g _24525_ (.A(_03463_), .B(_03465_), .Y(_00681_));
NAND_g _24526_ (.A(decoded_imm[26]), .B(_11223_), .Y(_03466_));
NAND_g _24527_ (.A(cached_insn_imm[26]), .B(decoder_pseudo_trigger_q), .Y(_03467_));
NOR_g _24528_ (.A(dbg_next), .B(q_insn_imm[26]), .Y(_03468_));
AND_g _24529_ (.A(dbg_next), .B(_03467_), .Y(_03469_));
AND_g _24530_ (.A(_03466_), .B(_03469_), .Y(_03470_));
NOR_g _24531_ (.A(_03468_), .B(_03470_), .Y(_00682_));
NAND_g _24532_ (.A(decoded_imm[27]), .B(_11223_), .Y(_03471_));
NAND_g _24533_ (.A(cached_insn_imm[27]), .B(decoder_pseudo_trigger_q), .Y(_03472_));
NOR_g _24534_ (.A(dbg_next), .B(q_insn_imm[27]), .Y(_03473_));
AND_g _24535_ (.A(dbg_next), .B(_03472_), .Y(_03474_));
AND_g _24536_ (.A(_03471_), .B(_03474_), .Y(_03475_));
NOR_g _24537_ (.A(_03473_), .B(_03475_), .Y(_00683_));
NAND_g _24538_ (.A(decoded_imm[28]), .B(_11223_), .Y(_03476_));
NAND_g _24539_ (.A(cached_insn_imm[28]), .B(decoder_pseudo_trigger_q), .Y(_03477_));
NOR_g _24540_ (.A(dbg_next), .B(q_insn_imm[28]), .Y(_03478_));
AND_g _24541_ (.A(dbg_next), .B(_03477_), .Y(_03479_));
AND_g _24542_ (.A(_03476_), .B(_03479_), .Y(_03480_));
NOR_g _24543_ (.A(_03478_), .B(_03480_), .Y(_00684_));
NAND_g _24544_ (.A(decoded_imm[29]), .B(_11223_), .Y(_03481_));
NAND_g _24545_ (.A(cached_insn_imm[29]), .B(decoder_pseudo_trigger_q), .Y(_03482_));
NOR_g _24546_ (.A(dbg_next), .B(q_insn_imm[29]), .Y(_03483_));
AND_g _24547_ (.A(dbg_next), .B(_03482_), .Y(_03484_));
AND_g _24548_ (.A(_03481_), .B(_03484_), .Y(_03485_));
NOR_g _24549_ (.A(_03483_), .B(_03485_), .Y(_00685_));
NAND_g _24550_ (.A(decoded_imm[30]), .B(_11223_), .Y(_03486_));
NAND_g _24551_ (.A(cached_insn_imm[30]), .B(decoder_pseudo_trigger_q), .Y(_03487_));
NOR_g _24552_ (.A(dbg_next), .B(q_insn_imm[30]), .Y(_03488_));
AND_g _24553_ (.A(dbg_next), .B(_03487_), .Y(_03489_));
AND_g _24554_ (.A(_03486_), .B(_03489_), .Y(_03490_));
NOR_g _24555_ (.A(_03488_), .B(_03490_), .Y(_00686_));
NAND_g _24556_ (.A(decoded_imm[31]), .B(_11223_), .Y(_03491_));
NAND_g _24557_ (.A(cached_insn_imm[31]), .B(decoder_pseudo_trigger_q), .Y(_03492_));
NOR_g _24558_ (.A(dbg_next), .B(q_insn_imm[31]), .Y(_03493_));
AND_g _24559_ (.A(dbg_next), .B(_03492_), .Y(_03494_));
AND_g _24560_ (.A(_03491_), .B(_03494_), .Y(_03495_));
NOR_g _24561_ (.A(_03493_), .B(_03495_), .Y(_00687_));
NAND_g _24562_ (.A(decoded_rd[0]), .B(_11223_), .Y(_03496_));
NAND_g _24563_ (.A(cached_insn_rd[0]), .B(decoder_pseudo_trigger_q), .Y(_03497_));
NOR_g _24564_ (.A(dbg_next), .B(q_insn_rd[0]), .Y(_03498_));
AND_g _24565_ (.A(dbg_next), .B(_03497_), .Y(_03499_));
AND_g _24566_ (.A(_03496_), .B(_03499_), .Y(_03500_));
NOR_g _24567_ (.A(_03498_), .B(_03500_), .Y(_00688_));
NAND_g _24568_ (.A(decoded_rd[1]), .B(_11223_), .Y(_03501_));
NAND_g _24569_ (.A(cached_insn_rd[1]), .B(decoder_pseudo_trigger_q), .Y(_03502_));
NOR_g _24570_ (.A(dbg_next), .B(q_insn_rd[1]), .Y(_03503_));
AND_g _24571_ (.A(dbg_next), .B(_03502_), .Y(_03504_));
AND_g _24572_ (.A(_03501_), .B(_03504_), .Y(_03505_));
NOR_g _24573_ (.A(_03503_), .B(_03505_), .Y(_00689_));
NAND_g _24574_ (.A(decoded_rd[2]), .B(_11223_), .Y(_03506_));
NAND_g _24575_ (.A(cached_insn_rd[2]), .B(decoder_pseudo_trigger_q), .Y(_03507_));
NOR_g _24576_ (.A(dbg_next), .B(q_insn_rd[2]), .Y(_03508_));
AND_g _24577_ (.A(dbg_next), .B(_03507_), .Y(_03509_));
AND_g _24578_ (.A(_03506_), .B(_03509_), .Y(_03510_));
NOR_g _24579_ (.A(_03508_), .B(_03510_), .Y(_00690_));
NAND_g _24580_ (.A(decoded_rd[3]), .B(_11223_), .Y(_03511_));
NAND_g _24581_ (.A(cached_insn_rd[3]), .B(decoder_pseudo_trigger_q), .Y(_03512_));
NOR_g _24582_ (.A(dbg_next), .B(q_insn_rd[3]), .Y(_03513_));
AND_g _24583_ (.A(dbg_next), .B(_03512_), .Y(_03514_));
AND_g _24584_ (.A(_03511_), .B(_03514_), .Y(_03515_));
NOR_g _24585_ (.A(_03513_), .B(_03515_), .Y(_00691_));
NAND_g _24586_ (.A(decoded_rd[4]), .B(_11223_), .Y(_03516_));
NAND_g _24587_ (.A(cached_insn_rd[4]), .B(decoder_pseudo_trigger_q), .Y(_03517_));
NOR_g _24588_ (.A(dbg_next), .B(q_insn_rd[4]), .Y(_03518_));
AND_g _24589_ (.A(dbg_next), .B(_03517_), .Y(_03519_));
AND_g _24590_ (.A(_03516_), .B(_03519_), .Y(_03520_));
NOR_g _24591_ (.A(_03518_), .B(_03520_), .Y(_00692_));
NAND_g _24592_ (.A(decoded_imm_j[15]), .B(_11223_), .Y(_03521_));
NAND_g _24593_ (.A(cached_insn_rs1[0]), .B(decoder_pseudo_trigger_q), .Y(_03522_));
NOR_g _24594_ (.A(dbg_next), .B(q_insn_rs1[0]), .Y(_03523_));
AND_g _24595_ (.A(dbg_next), .B(_03522_), .Y(_03524_));
AND_g _24596_ (.A(_03521_), .B(_03524_), .Y(_03525_));
NOR_g _24597_ (.A(_03523_), .B(_03525_), .Y(_00693_));
NAND_g _24598_ (.A(decoded_imm_j[16]), .B(_11223_), .Y(_03526_));
NAND_g _24599_ (.A(cached_insn_rs1[1]), .B(decoder_pseudo_trigger_q), .Y(_03527_));
NOR_g _24600_ (.A(dbg_next), .B(q_insn_rs1[1]), .Y(_03528_));
AND_g _24601_ (.A(dbg_next), .B(_03527_), .Y(_03529_));
AND_g _24602_ (.A(_03526_), .B(_03529_), .Y(_03530_));
NOR_g _24603_ (.A(_03528_), .B(_03530_), .Y(_00694_));
NAND_g _24604_ (.A(decoded_imm_j[17]), .B(_11223_), .Y(_03531_));
NAND_g _24605_ (.A(cached_insn_rs1[2]), .B(decoder_pseudo_trigger_q), .Y(_03532_));
NOR_g _24606_ (.A(dbg_next), .B(q_insn_rs1[2]), .Y(_03533_));
AND_g _24607_ (.A(dbg_next), .B(_03532_), .Y(_03534_));
AND_g _24608_ (.A(_03531_), .B(_03534_), .Y(_03535_));
NOR_g _24609_ (.A(_03533_), .B(_03535_), .Y(_00695_));
NAND_g _24610_ (.A(decoded_imm_j[18]), .B(_11223_), .Y(_03536_));
NAND_g _24611_ (.A(cached_insn_rs1[3]), .B(decoder_pseudo_trigger_q), .Y(_03537_));
NOR_g _24612_ (.A(dbg_next), .B(q_insn_rs1[3]), .Y(_03538_));
AND_g _24613_ (.A(dbg_next), .B(_03537_), .Y(_03539_));
AND_g _24614_ (.A(_03536_), .B(_03539_), .Y(_03540_));
NOR_g _24615_ (.A(_03538_), .B(_03540_), .Y(_00696_));
NAND_g _24616_ (.A(decoded_imm_j[19]), .B(_11223_), .Y(_03541_));
NAND_g _24617_ (.A(cached_insn_rs1[4]), .B(decoder_pseudo_trigger_q), .Y(_03542_));
NOR_g _24618_ (.A(dbg_next), .B(q_insn_rs1[4]), .Y(_03543_));
AND_g _24619_ (.A(dbg_next), .B(_03542_), .Y(_03544_));
AND_g _24620_ (.A(_03541_), .B(_03544_), .Y(_03545_));
NOR_g _24621_ (.A(_03543_), .B(_03545_), .Y(_00697_));
NAND_g _24622_ (.A(decoded_rd[0]), .B(decoder_trigger_q), .Y(_03546_));
NAND_g _24623_ (.A(cached_insn_rd[0]), .B(_11045_), .Y(_03547_));
NAND_g _24624_ (.A(_03546_), .B(_03547_), .Y(_00698_));
NAND_g _24625_ (.A(decoded_rd[1]), .B(decoder_trigger_q), .Y(_03548_));
NAND_g _24626_ (.A(_11045_), .B(cached_insn_rd[1]), .Y(_03549_));
NAND_g _24627_ (.A(_03548_), .B(_03549_), .Y(_00699_));
NAND_g _24628_ (.A(decoded_rd[2]), .B(decoder_trigger_q), .Y(_03550_));
NAND_g _24629_ (.A(_11045_), .B(cached_insn_rd[2]), .Y(_03551_));
NAND_g _24630_ (.A(_03550_), .B(_03551_), .Y(_00700_));
NAND_g _24631_ (.A(decoded_rd[3]), .B(decoder_trigger_q), .Y(_03552_));
NAND_g _24632_ (.A(_11045_), .B(cached_insn_rd[3]), .Y(_03553_));
NAND_g _24633_ (.A(_03552_), .B(_03553_), .Y(_00701_));
NAND_g _24634_ (.A(decoded_rd[4]), .B(decoder_trigger_q), .Y(_03554_));
NAND_g _24635_ (.A(_11045_), .B(cached_insn_rd[4]), .Y(_03555_));
NAND_g _24636_ (.A(_03554_), .B(_03555_), .Y(_00702_));
NAND_g _24637_ (.A(decoded_imm[0]), .B(decoder_trigger_q), .Y(_03556_));
NAND_g _24638_ (.A(_11045_), .B(cached_insn_imm[0]), .Y(_03557_));
NAND_g _24639_ (.A(_03556_), .B(_03557_), .Y(_00703_));
NAND_g _24640_ (.A(decoder_trigger_q), .B(decoded_imm[1]), .Y(_03558_));
NAND_g _24641_ (.A(_11045_), .B(cached_insn_imm[1]), .Y(_03559_));
NAND_g _24642_ (.A(_03558_), .B(_03559_), .Y(_00704_));
NAND_g _24643_ (.A(decoder_trigger_q), .B(decoded_imm[2]), .Y(_03560_));
NAND_g _24644_ (.A(_11045_), .B(cached_insn_imm[2]), .Y(_03561_));
NAND_g _24645_ (.A(_03560_), .B(_03561_), .Y(_00705_));
NAND_g _24646_ (.A(decoder_trigger_q), .B(decoded_imm[3]), .Y(_03562_));
NAND_g _24647_ (.A(_11045_), .B(cached_insn_imm[3]), .Y(_03563_));
NAND_g _24648_ (.A(_03562_), .B(_03563_), .Y(_00706_));
NAND_g _24649_ (.A(decoder_trigger_q), .B(decoded_imm[4]), .Y(_03564_));
NAND_g _24650_ (.A(_11045_), .B(cached_insn_imm[4]), .Y(_03565_));
NAND_g _24651_ (.A(_03564_), .B(_03565_), .Y(_00707_));
NAND_g _24652_ (.A(decoder_trigger_q), .B(decoded_imm[5]), .Y(_03566_));
NAND_g _24653_ (.A(_11045_), .B(cached_insn_imm[5]), .Y(_03567_));
NAND_g _24654_ (.A(_03566_), .B(_03567_), .Y(_00708_));
NAND_g _24655_ (.A(decoder_trigger_q), .B(decoded_imm[6]), .Y(_03568_));
NAND_g _24656_ (.A(_11045_), .B(cached_insn_imm[6]), .Y(_03569_));
NAND_g _24657_ (.A(_03568_), .B(_03569_), .Y(_00709_));
NAND_g _24658_ (.A(decoder_trigger_q), .B(decoded_imm[7]), .Y(_03570_));
NAND_g _24659_ (.A(_11045_), .B(cached_insn_imm[7]), .Y(_03571_));
NAND_g _24660_ (.A(_03570_), .B(_03571_), .Y(_00710_));
NAND_g _24661_ (.A(decoder_trigger_q), .B(decoded_imm[8]), .Y(_03572_));
NAND_g _24662_ (.A(_11045_), .B(cached_insn_imm[8]), .Y(_03573_));
NAND_g _24663_ (.A(_03572_), .B(_03573_), .Y(_00711_));
NAND_g _24664_ (.A(decoder_trigger_q), .B(decoded_imm[9]), .Y(_03574_));
NAND_g _24665_ (.A(_11045_), .B(cached_insn_imm[9]), .Y(_03575_));
NAND_g _24666_ (.A(_03574_), .B(_03575_), .Y(_00712_));
NAND_g _24667_ (.A(decoder_trigger_q), .B(decoded_imm[10]), .Y(_03576_));
NAND_g _24668_ (.A(_11045_), .B(cached_insn_imm[10]), .Y(_03577_));
NAND_g _24669_ (.A(_03576_), .B(_03577_), .Y(_00713_));
NAND_g _24670_ (.A(decoder_trigger_q), .B(decoded_imm[11]), .Y(_03578_));
NAND_g _24671_ (.A(_11045_), .B(cached_insn_imm[11]), .Y(_03579_));
NAND_g _24672_ (.A(_03578_), .B(_03579_), .Y(_00714_));
NAND_g _24673_ (.A(decoder_trigger_q), .B(decoded_imm[12]), .Y(_03580_));
NAND_g _24674_ (.A(_11045_), .B(cached_insn_imm[12]), .Y(_03581_));
NAND_g _24675_ (.A(_03580_), .B(_03581_), .Y(_00715_));
NAND_g _24676_ (.A(decoder_trigger_q), .B(decoded_imm[13]), .Y(_03582_));
NAND_g _24677_ (.A(_11045_), .B(cached_insn_imm[13]), .Y(_03583_));
NAND_g _24678_ (.A(_03582_), .B(_03583_), .Y(_00716_));
NAND_g _24679_ (.A(decoder_trigger_q), .B(decoded_imm[14]), .Y(_03584_));
NAND_g _24680_ (.A(_11045_), .B(cached_insn_imm[14]), .Y(_03585_));
NAND_g _24681_ (.A(_03584_), .B(_03585_), .Y(_00717_));
NAND_g _24682_ (.A(decoder_trigger_q), .B(decoded_imm[15]), .Y(_03586_));
NAND_g _24683_ (.A(_11045_), .B(cached_insn_imm[15]), .Y(_03587_));
NAND_g _24684_ (.A(_03586_), .B(_03587_), .Y(_00718_));
NAND_g _24685_ (.A(decoder_trigger_q), .B(decoded_imm[16]), .Y(_03588_));
NAND_g _24686_ (.A(_11045_), .B(cached_insn_imm[16]), .Y(_03589_));
NAND_g _24687_ (.A(_03588_), .B(_03589_), .Y(_00719_));
NAND_g _24688_ (.A(decoder_trigger_q), .B(decoded_imm[17]), .Y(_03590_));
NAND_g _24689_ (.A(_11045_), .B(cached_insn_imm[17]), .Y(_03591_));
NAND_g _24690_ (.A(_03590_), .B(_03591_), .Y(_00720_));
NAND_g _24691_ (.A(decoder_trigger_q), .B(decoded_imm[18]), .Y(_03592_));
NAND_g _24692_ (.A(_11045_), .B(cached_insn_imm[18]), .Y(_03593_));
NAND_g _24693_ (.A(_03592_), .B(_03593_), .Y(_00721_));
NAND_g _24694_ (.A(decoder_trigger_q), .B(decoded_imm[19]), .Y(_03594_));
NAND_g _24695_ (.A(_11045_), .B(cached_insn_imm[19]), .Y(_03595_));
NAND_g _24696_ (.A(_03594_), .B(_03595_), .Y(_00722_));
NAND_g _24697_ (.A(decoder_trigger_q), .B(decoded_imm[20]), .Y(_03596_));
NAND_g _24698_ (.A(_11045_), .B(cached_insn_imm[20]), .Y(_03597_));
NAND_g _24699_ (.A(_03596_), .B(_03597_), .Y(_00723_));
NAND_g _24700_ (.A(decoder_trigger_q), .B(decoded_imm[21]), .Y(_03598_));
NAND_g _24701_ (.A(_11045_), .B(cached_insn_imm[21]), .Y(_03599_));
NAND_g _24702_ (.A(_03598_), .B(_03599_), .Y(_00724_));
NAND_g _24703_ (.A(decoder_trigger_q), .B(decoded_imm[22]), .Y(_03600_));
NAND_g _24704_ (.A(_11045_), .B(cached_insn_imm[22]), .Y(_03601_));
NAND_g _24705_ (.A(_03600_), .B(_03601_), .Y(_00725_));
NAND_g _24706_ (.A(decoder_trigger_q), .B(decoded_imm[23]), .Y(_03602_));
NAND_g _24707_ (.A(_11045_), .B(cached_insn_imm[23]), .Y(_03603_));
NAND_g _24708_ (.A(_03602_), .B(_03603_), .Y(_00726_));
NAND_g _24709_ (.A(decoder_trigger_q), .B(decoded_imm[24]), .Y(_03604_));
NAND_g _24710_ (.A(_11045_), .B(cached_insn_imm[24]), .Y(_03605_));
NAND_g _24711_ (.A(_03604_), .B(_03605_), .Y(_00727_));
NAND_g _24712_ (.A(decoder_trigger_q), .B(decoded_imm[25]), .Y(_03606_));
NAND_g _24713_ (.A(_11045_), .B(cached_insn_imm[25]), .Y(_03607_));
NAND_g _24714_ (.A(_03606_), .B(_03607_), .Y(_00728_));
NAND_g _24715_ (.A(decoder_trigger_q), .B(decoded_imm[26]), .Y(_03608_));
NAND_g _24716_ (.A(_11045_), .B(cached_insn_imm[26]), .Y(_03609_));
NAND_g _24717_ (.A(_03608_), .B(_03609_), .Y(_00729_));
NAND_g _24718_ (.A(decoder_trigger_q), .B(decoded_imm[27]), .Y(_03610_));
NAND_g _24719_ (.A(_11045_), .B(cached_insn_imm[27]), .Y(_03611_));
NAND_g _24720_ (.A(_03610_), .B(_03611_), .Y(_00730_));
NAND_g _24721_ (.A(decoder_trigger_q), .B(decoded_imm[28]), .Y(_03612_));
NAND_g _24722_ (.A(_11045_), .B(cached_insn_imm[28]), .Y(_03613_));
NAND_g _24723_ (.A(_03612_), .B(_03613_), .Y(_00731_));
NAND_g _24724_ (.A(decoder_trigger_q), .B(decoded_imm[29]), .Y(_03614_));
NAND_g _24725_ (.A(_11045_), .B(cached_insn_imm[29]), .Y(_03615_));
NAND_g _24726_ (.A(_03614_), .B(_03615_), .Y(_00732_));
NAND_g _24727_ (.A(decoder_trigger_q), .B(decoded_imm[30]), .Y(_03616_));
NAND_g _24728_ (.A(_11045_), .B(cached_insn_imm[30]), .Y(_03617_));
NAND_g _24729_ (.A(_03616_), .B(_03617_), .Y(_00733_));
NAND_g _24730_ (.A(decoder_trigger_q), .B(decoded_imm[31]), .Y(_03618_));
NAND_g _24731_ (.A(_11045_), .B(cached_insn_imm[31]), .Y(_03619_));
NAND_g _24732_ (.A(_03618_), .B(_03619_), .Y(_00734_));
NAND_g _24733_ (.A(decoder_trigger_q), .B(decoded_imm_j[15]), .Y(_03620_));
NAND_g _24734_ (.A(_11045_), .B(cached_insn_rs1[0]), .Y(_03621_));
NAND_g _24735_ (.A(_03620_), .B(_03621_), .Y(_00735_));
NAND_g _24736_ (.A(decoder_trigger_q), .B(decoded_imm_j[16]), .Y(_03622_));
NAND_g _24737_ (.A(_11045_), .B(cached_insn_rs1[1]), .Y(_03623_));
NAND_g _24738_ (.A(_03622_), .B(_03623_), .Y(_00736_));
NAND_g _24739_ (.A(decoder_trigger_q), .B(decoded_imm_j[17]), .Y(_03624_));
NAND_g _24740_ (.A(_11045_), .B(cached_insn_rs1[2]), .Y(_03625_));
NAND_g _24741_ (.A(_03624_), .B(_03625_), .Y(_00737_));
NAND_g _24742_ (.A(decoder_trigger_q), .B(decoded_imm_j[18]), .Y(_03626_));
NAND_g _24743_ (.A(_11045_), .B(cached_insn_rs1[3]), .Y(_03627_));
NAND_g _24744_ (.A(_03626_), .B(_03627_), .Y(_00738_));
NAND_g _24745_ (.A(decoder_trigger_q), .B(decoded_imm_j[19]), .Y(_03628_));
NAND_g _24746_ (.A(_11045_), .B(cached_insn_rs1[4]), .Y(_03629_));
NAND_g _24747_ (.A(_03628_), .B(_03629_), .Y(_00739_));
NAND_g _24748_ (.A(decoded_imm_j[11]), .B(decoder_trigger_q), .Y(_03630_));
NAND_g _24749_ (.A(_11045_), .B(cached_insn_rs2[0]), .Y(_03631_));
NAND_g _24750_ (.A(_03630_), .B(_03631_), .Y(_00740_));
NAND_g _24751_ (.A(decoded_imm_j[1]), .B(decoder_trigger_q), .Y(_03632_));
NAND_g _24752_ (.A(_11045_), .B(cached_insn_rs2[1]), .Y(_03633_));
NAND_g _24753_ (.A(_03632_), .B(_03633_), .Y(_00741_));
NAND_g _24754_ (.A(decoded_imm_j[2]), .B(decoder_trigger_q), .Y(_03634_));
NAND_g _24755_ (.A(_11045_), .B(cached_insn_rs2[2]), .Y(_03635_));
NAND_g _24756_ (.A(_03634_), .B(_03635_), .Y(_00742_));
NAND_g _24757_ (.A(decoded_imm_j[3]), .B(decoder_trigger_q), .Y(_03636_));
NAND_g _24758_ (.A(_11045_), .B(cached_insn_rs2[3]), .Y(_03637_));
NAND_g _24759_ (.A(_03636_), .B(_03637_), .Y(_00743_));
NAND_g _24760_ (.A(decoder_trigger_q), .B(decoded_imm_j[4]), .Y(_03638_));
NAND_g _24761_ (.A(_11045_), .B(cached_insn_rs2[4]), .Y(_03639_));
NAND_g _24762_ (.A(_03638_), .B(_03639_), .Y(_00744_));
NAND_g _24763_ (.A(_11045_), .B(cached_ascii_instr[0]), .Y(_03640_));
NAND_g _24764_ (.A(decoder_trigger_q), .B(_02846_), .Y(_03641_));
NAND_g _24765_ (.A(_03640_), .B(_03641_), .Y(_00745_));
NAND_g _24766_ (.A(_11045_), .B(cached_ascii_instr[1]), .Y(_03642_));
AND_g _24767_ (.A(_10975_), .B(decoder_trigger_q), .Y(_03643_));
NAND_g _24768_ (.A(_02882_), .B(_03643_), .Y(_03644_));
NAND_g _24769_ (.A(_03642_), .B(_03644_), .Y(_00746_));
NAND_g _24770_ (.A(_11045_), .B(cached_ascii_instr[2]), .Y(_03645_));
NAND_g _24771_ (.A(decoder_trigger_q), .B(_02907_), .Y(_03646_));
NAND_g _24772_ (.A(_03645_), .B(_03646_), .Y(_00747_));
AND_g _24773_ (.A(_02914_), .B(_03643_), .Y(_03647_));
NAND_g _24774_ (.A(_02938_), .B(_03647_), .Y(_03648_));
NAND_g _24775_ (.A(_11045_), .B(_11053_), .Y(_03649_));
AND_g _24776_ (.A(_03648_), .B(_03649_), .Y(_00748_));
NAND_g _24777_ (.A(_11045_), .B(cached_ascii_instr[4]), .Y(_03650_));
NAND_g _24778_ (.A(_02958_), .B(_03643_), .Y(_03651_));
NAND_g _24779_ (.A(_03650_), .B(_03651_), .Y(_00749_));
NAND_g _24780_ (.A(_11045_), .B(_11055_), .Y(_03652_));
NOR_g _24781_ (.A(_11045_), .B(_02965_), .Y(_03653_));
NAND_g _24782_ (.A(_02989_), .B(_03653_), .Y(_03654_));
AND_g _24783_ (.A(_03652_), .B(_03654_), .Y(_00750_));
NAND_g _24784_ (.A(_03007_), .B(_03643_), .Y(_03655_));
NAND_g _24785_ (.A(_11045_), .B(_11056_), .Y(_03656_));
AND_g _24786_ (.A(_03655_), .B(_03656_), .Y(_00751_));
NAND_g _24787_ (.A(_11045_), .B(cached_ascii_instr[10]), .Y(_03657_));
NAND_g _24788_ (.A(_03027_), .B(_03643_), .Y(_03658_));
NAND_g _24789_ (.A(_03657_), .B(_03658_), .Y(_00752_));
NAND_g _24790_ (.A(_11045_), .B(cached_ascii_instr[11]), .Y(_03659_));
NAND_g _24791_ (.A(decoder_trigger_q), .B(_03053_), .Y(_03660_));
NAND_g _24792_ (.A(_03659_), .B(_03660_), .Y(_00753_));
NAND_g _24793_ (.A(decoder_trigger_q), .B(_03081_), .Y(_03661_));
NAND_g _24794_ (.A(_11045_), .B(_11059_), .Y(_03662_));
AND_g _24795_ (.A(_03661_), .B(_03662_), .Y(_00754_));
NAND_g _24796_ (.A(_11045_), .B(cached_ascii_instr[14]), .Y(_03663_));
NAND_g _24797_ (.A(decoder_trigger_q), .B(_13610_), .Y(_03664_));
NAND_g _24798_ (.A(_03663_), .B(_03664_), .Y(_00755_));
NAND_g _24799_ (.A(_11045_), .B(cached_ascii_instr[16]), .Y(_03665_));
NAND_g _24800_ (.A(_03102_), .B(_03647_), .Y(_03666_));
NAND_g _24801_ (.A(_03665_), .B(_03666_), .Y(_00756_));
NAND_g _24802_ (.A(_11045_), .B(_11061_), .Y(_03667_));
NOR_g _24803_ (.A(_11045_), .B(_03123_), .Y(_03668_));
NAND_g _24804_ (.A(_03122_), .B(_03668_), .Y(_03669_));
AND_g _24805_ (.A(_03667_), .B(_03669_), .Y(_00757_));
NAND_g _24806_ (.A(_03141_), .B(_03647_), .Y(_03670_));
NAND_g _24807_ (.A(_11045_), .B(_11062_), .Y(_03671_));
AND_g _24808_ (.A(_03670_), .B(_03671_), .Y(_00758_));
NAND_g _24809_ (.A(_11045_), .B(_11063_), .Y(_03672_));
NAND_g _24810_ (.A(_03160_), .B(_03653_), .Y(_03673_));
AND_g _24811_ (.A(_03672_), .B(_03673_), .Y(_00759_));
NAND_g _24812_ (.A(decoder_trigger_q), .B(_03174_), .Y(_03674_));
NAND_g _24813_ (.A(_11045_), .B(_11064_), .Y(_03675_));
AND_g _24814_ (.A(_03674_), .B(_03675_), .Y(_00760_));
NAND_g _24815_ (.A(decoder_trigger_q), .B(_03188_), .Y(_03676_));
NAND_g _24816_ (.A(_11045_), .B(_11065_), .Y(_03677_));
AND_g _24817_ (.A(_03676_), .B(_03677_), .Y(_00761_));
NAND_g _24818_ (.A(_03203_), .B(_03643_), .Y(_03678_));
NAND_g _24819_ (.A(_11045_), .B(_11066_), .Y(_03679_));
AND_g _24820_ (.A(_03678_), .B(_03679_), .Y(_00762_));
NAND_g _24821_ (.A(_11045_), .B(_11067_), .Y(_03680_));
AND_g _24822_ (.A(decoder_trigger_q), .B(_13564_), .Y(_03681_));
NAND_g _24823_ (.A(_03219_), .B(_03681_), .Y(_03682_));
AND_g _24824_ (.A(_03680_), .B(_03682_), .Y(_00763_));
NAND_g _24825_ (.A(_11045_), .B(cached_ascii_instr[26]), .Y(_03683_));
NAND_g _24826_ (.A(_03230_), .B(_03647_), .Y(_03684_));
NAND_g _24827_ (.A(_03683_), .B(_03684_), .Y(_00764_));
NAND_g _24828_ (.A(_11045_), .B(_11069_), .Y(_03685_));
NAND_g _24829_ (.A(_03244_), .B(_03668_), .Y(_03686_));
AND_g _24830_ (.A(_03685_), .B(_03686_), .Y(_00765_));
NAND_g _24831_ (.A(_03261_), .B(_03643_), .Y(_03687_));
NAND_g _24832_ (.A(_11045_), .B(_11070_), .Y(_03688_));
AND_g _24833_ (.A(_03687_), .B(_03688_), .Y(_00766_));
NAND_g _24834_ (.A(_11045_), .B(_11071_), .Y(_03689_));
NAND_g _24835_ (.A(decoder_trigger_q), .B(_03276_), .Y(_03690_));
AND_g _24836_ (.A(_03689_), .B(_03690_), .Y(_00767_));
NAND_g _24837_ (.A(_11045_), .B(cached_ascii_instr[32]), .Y(_03691_));
NAND_g _24838_ (.A(_03283_), .B(_03643_), .Y(_03692_));
NAND_g _24839_ (.A(_03691_), .B(_03692_), .Y(_00768_));
NAND_g _24840_ (.A(_03295_), .B(_03643_), .Y(_03693_));
NAND_g _24841_ (.A(_11045_), .B(_11073_), .Y(_03694_));
AND_g _24842_ (.A(_03693_), .B(_03694_), .Y(_00769_));
NOR_g _24843_ (.A(decoder_trigger_q), .B(cached_ascii_instr[35]), .Y(_03695_));
NOR_g _24844_ (.A(_03681_), .B(_03695_), .Y(_00770_));
NAND_g _24845_ (.A(_11045_), .B(_11075_), .Y(_03696_));
NAND_g _24846_ (.A(_03305_), .B(_03653_), .Y(_03697_));
AND_g _24847_ (.A(_03696_), .B(_03697_), .Y(_00771_));
NAND_g _24848_ (.A(_03282_), .B(_03643_), .Y(_03698_));
NAND_g _24849_ (.A(_11045_), .B(_11076_), .Y(_03699_));
AND_g _24850_ (.A(_03698_), .B(_03699_), .Y(_00772_));
NOR_g _24851_ (.A(decoder_trigger_q), .B(cached_ascii_instr[41]), .Y(_03700_));
NOR_g _24852_ (.A(_03653_), .B(_03700_), .Y(_00773_));
NOR_g _24853_ (.A(decoder_trigger_q), .B(cached_ascii_instr[43]), .Y(_03701_));
NOR_g _24854_ (.A(_03643_), .B(_03701_), .Y(_00774_));
NOR_g _24855_ (.A(decoder_trigger_q), .B(cached_ascii_instr[52]), .Y(_03702_));
NOR_g _24856_ (.A(_03668_), .B(_03702_), .Y(_00775_));
AND_g _24857_ (.A(decoder_trigger_q), .B(_13565_), .Y(_03703_));
NOR_g _24858_ (.A(decoder_trigger_q), .B(cached_ascii_instr[54]), .Y(_03704_));
NOR_g _24859_ (.A(_03703_), .B(_03704_), .Y(_00776_));
NOR_g _24860_ (.A(decoder_trigger_q), .B(cached_ascii_instr[62]), .Y(_03705_));
NOR_g _24861_ (.A(_03647_), .B(_03705_), .Y(_00777_));
NAND_g _24862_ (.A(mem_instr), .B(_02603_), .Y(_03706_));
AND_g _24863_ (.A(_10893_), .B(_02599_), .Y(_03707_));
NAND_g _24864_ (.A(_02594_), .B(_03707_), .Y(_03708_));
NAND_g _24865_ (.A(_03706_), .B(_03708_), .Y(_00778_));
NAND_g _24866_ (.A(mem_rdata[15]), .B(_11910_), .Y(_03709_));
NAND_g _24867_ (.A(mem_rdata_q[15]), .B(_11911_), .Y(_03710_));
NAND_g _24868_ (.A(_03709_), .B(_03710_), .Y(_00787_));
NAND_g _24869_ (.A(mem_rdata[16]), .B(_11910_), .Y(_03711_));
NAND_g _24870_ (.A(mem_rdata_q[16]), .B(_11911_), .Y(_03712_));
NAND_g _24871_ (.A(_03711_), .B(_03712_), .Y(_00788_));
NAND_g _24872_ (.A(mem_rdata[17]), .B(_11910_), .Y(_03713_));
NAND_g _24873_ (.A(mem_rdata_q[17]), .B(_11911_), .Y(_03714_));
NAND_g _24874_ (.A(_03713_), .B(_03714_), .Y(_00789_));
NAND_g _24875_ (.A(mem_rdata[18]), .B(_11910_), .Y(_03715_));
NAND_g _24876_ (.A(mem_rdata_q[18]), .B(_11911_), .Y(_03716_));
NAND_g _24877_ (.A(_03715_), .B(_03716_), .Y(_00790_));
NAND_g _24878_ (.A(mem_rdata[19]), .B(_11910_), .Y(_03717_));
NAND_g _24879_ (.A(mem_rdata_q[19]), .B(_11911_), .Y(_03718_));
NAND_g _24880_ (.A(_03717_), .B(_03718_), .Y(_00791_));
NAND_g _24881_ (.A(mem_rdata[24]), .B(_11910_), .Y(_03719_));
NAND_g _24882_ (.A(mem_rdata_q[24]), .B(_11911_), .Y(_03720_));
NAND_g _24883_ (.A(_03719_), .B(_03720_), .Y(_00796_));
NAND_g _24884_ (.A(mem_rdata[26]), .B(_11910_), .Y(_03721_));
NAND_g _24885_ (.A(mem_rdata_q[26]), .B(_11911_), .Y(_03722_));
NAND_g _24886_ (.A(_03721_), .B(_03722_), .Y(_00798_));
NAND_g _24887_ (.A(mem_rdata[27]), .B(_11910_), .Y(_03723_));
NAND_g _24888_ (.A(mem_rdata_q[27]), .B(_11911_), .Y(_03724_));
NAND_g _24889_ (.A(_03723_), .B(_03724_), .Y(_00799_));
NAND_g _24890_ (.A(mem_rdata[30]), .B(_11910_), .Y(_03725_));
NAND_g _24891_ (.A(mem_rdata_q[30]), .B(_11911_), .Y(_03726_));
NAND_g _24892_ (.A(_03725_), .B(_03726_), .Y(_00802_));
NAND_g _24893_ (.A(mem_rdata[31]), .B(_11910_), .Y(_03727_));
NAND_g _24894_ (.A(mem_rdata_q[31]), .B(_11911_), .Y(_03728_));
NAND_g _24895_ (.A(_03727_), .B(_03728_), .Y(_00803_));
NAND_g _24896_ (.A(reg_out[2]), .B(_12542_), .Y(_03729_));
NAND_g _24897_ (.A(_12551_), .B(_03729_), .Y(_03730_));
NAND_g _24898_ (.A(_02594_), .B(_03730_), .Y(_03731_));
NAND_g _24899_ (.A(pcpi_rs1[2]), .B(_02593_), .Y(_03732_));
NAND_g _24900_ (.A(_03731_), .B(_03732_), .Y(mem_la_addr[2]));
NAND_g _24901_ (.A(_02602_), .B(mem_la_addr[2]), .Y(_03733_));
NAND_g _24902_ (.A(mem_addr[2]), .B(_02603_), .Y(_03734_));
NAND_g _24903_ (.A(_03733_), .B(_03734_), .Y(_00804_));
NAND_g _24904_ (.A(reg_out[3]), .B(_12542_), .Y(_03735_));
NAND_g _24905_ (.A(_12557_), .B(_03735_), .Y(_03736_));
NAND_g _24906_ (.A(_02594_), .B(_03736_), .Y(_03737_));
NAND_g _24907_ (.A(pcpi_rs1[3]), .B(_02593_), .Y(_03738_));
NAND_g _24908_ (.A(_03737_), .B(_03738_), .Y(mem_la_addr[3]));
NAND_g _24909_ (.A(_02602_), .B(mem_la_addr[3]), .Y(_03739_));
NAND_g _24910_ (.A(mem_addr[3]), .B(_02603_), .Y(_03740_));
NAND_g _24911_ (.A(_03739_), .B(_03740_), .Y(_00805_));
NAND_g _24912_ (.A(reg_out[4]), .B(_12542_), .Y(_03741_));
NAND_g _24913_ (.A(_12563_), .B(_03741_), .Y(_03742_));
NAND_g _24914_ (.A(_02594_), .B(_03742_), .Y(_03743_));
NAND_g _24915_ (.A(pcpi_rs1[4]), .B(_02593_), .Y(_03744_));
NAND_g _24916_ (.A(_03743_), .B(_03744_), .Y(mem_la_addr[4]));
NAND_g _24917_ (.A(mem_addr[4]), .B(_02603_), .Y(_03745_));
NAND_g _24918_ (.A(_02602_), .B(mem_la_addr[4]), .Y(_03746_));
NAND_g _24919_ (.A(_03745_), .B(_03746_), .Y(_00806_));
NAND_g _24920_ (.A(reg_out[5]), .B(_12542_), .Y(_03747_));
NAND_g _24921_ (.A(_12569_), .B(_03747_), .Y(_03748_));
NAND_g _24922_ (.A(_02594_), .B(_03748_), .Y(_03749_));
NAND_g _24923_ (.A(pcpi_rs1[5]), .B(_02593_), .Y(_03750_));
NAND_g _24924_ (.A(_03749_), .B(_03750_), .Y(mem_la_addr[5]));
NAND_g _24925_ (.A(_02602_), .B(mem_la_addr[5]), .Y(_03751_));
NAND_g _24926_ (.A(mem_addr[5]), .B(_02603_), .Y(_03752_));
NAND_g _24927_ (.A(_03751_), .B(_03752_), .Y(_00807_));
NAND_g _24928_ (.A(reg_out[6]), .B(_12542_), .Y(_03753_));
NAND_g _24929_ (.A(_12575_), .B(_03753_), .Y(_03754_));
NAND_g _24930_ (.A(_02594_), .B(_03754_), .Y(_03755_));
NAND_g _24931_ (.A(pcpi_rs1[6]), .B(_02593_), .Y(_03756_));
NAND_g _24932_ (.A(_03755_), .B(_03756_), .Y(mem_la_addr[6]));
NAND_g _24933_ (.A(_02602_), .B(mem_la_addr[6]), .Y(_03757_));
NAND_g _24934_ (.A(mem_addr[6]), .B(_02603_), .Y(_03758_));
NAND_g _24935_ (.A(_03757_), .B(_03758_), .Y(_00808_));
NAND_g _24936_ (.A(reg_out[7]), .B(_12542_), .Y(_03759_));
NAND_g _24937_ (.A(_12581_), .B(_03759_), .Y(_03760_));
NAND_g _24938_ (.A(_02594_), .B(_03760_), .Y(_03761_));
NAND_g _24939_ (.A(pcpi_rs1[7]), .B(_02593_), .Y(_03762_));
NAND_g _24940_ (.A(_03761_), .B(_03762_), .Y(mem_la_addr[7]));
NAND_g _24941_ (.A(_02602_), .B(mem_la_addr[7]), .Y(_03763_));
NAND_g _24942_ (.A(mem_addr[7]), .B(_02603_), .Y(_03764_));
NAND_g _24943_ (.A(_03763_), .B(_03764_), .Y(_00809_));
NAND_g _24944_ (.A(reg_out[8]), .B(_12542_), .Y(_03765_));
NAND_g _24945_ (.A(_12587_), .B(_03765_), .Y(_03766_));
NAND_g _24946_ (.A(_02594_), .B(_03766_), .Y(_03767_));
NAND_g _24947_ (.A(pcpi_rs1[8]), .B(_02593_), .Y(_03768_));
NAND_g _24948_ (.A(_03767_), .B(_03768_), .Y(mem_la_addr[8]));
NAND_g _24949_ (.A(_02602_), .B(mem_la_addr[8]), .Y(_03769_));
NAND_g _24950_ (.A(mem_addr[8]), .B(_02603_), .Y(_03770_));
NAND_g _24951_ (.A(_03769_), .B(_03770_), .Y(_00810_));
NAND_g _24952_ (.A(reg_out[9]), .B(_12542_), .Y(_03771_));
NAND_g _24953_ (.A(_12593_), .B(_03771_), .Y(_03772_));
NAND_g _24954_ (.A(_02594_), .B(_03772_), .Y(_03773_));
NAND_g _24955_ (.A(pcpi_rs1[9]), .B(_02593_), .Y(_03774_));
NAND_g _24956_ (.A(_03773_), .B(_03774_), .Y(mem_la_addr[9]));
NAND_g _24957_ (.A(_02602_), .B(mem_la_addr[9]), .Y(_03775_));
NAND_g _24958_ (.A(mem_addr[9]), .B(_02603_), .Y(_03776_));
NAND_g _24959_ (.A(_03775_), .B(_03776_), .Y(_00811_));
NAND_g _24960_ (.A(reg_out[10]), .B(_12542_), .Y(_03777_));
NAND_g _24961_ (.A(_12599_), .B(_03777_), .Y(_03778_));
NAND_g _24962_ (.A(_02594_), .B(_03778_), .Y(_03779_));
NAND_g _24963_ (.A(pcpi_rs1[10]), .B(_02593_), .Y(_03780_));
NAND_g _24964_ (.A(_03779_), .B(_03780_), .Y(mem_la_addr[10]));
NAND_g _24965_ (.A(mem_addr[10]), .B(_02603_), .Y(_03781_));
NAND_g _24966_ (.A(_02602_), .B(mem_la_addr[10]), .Y(_03782_));
NAND_g _24967_ (.A(_03781_), .B(_03782_), .Y(_00812_));
NAND_g _24968_ (.A(reg_out[11]), .B(_12542_), .Y(_03783_));
NAND_g _24969_ (.A(_12605_), .B(_03783_), .Y(_03784_));
NAND_g _24970_ (.A(_02594_), .B(_03784_), .Y(_03785_));
NAND_g _24971_ (.A(pcpi_rs1[11]), .B(_02593_), .Y(_03786_));
NAND_g _24972_ (.A(_03785_), .B(_03786_), .Y(mem_la_addr[11]));
NAND_g _24973_ (.A(_02602_), .B(mem_la_addr[11]), .Y(_03787_));
NAND_g _24974_ (.A(mem_addr[11]), .B(_02603_), .Y(_03788_));
NAND_g _24975_ (.A(_03787_), .B(_03788_), .Y(_00813_));
NAND_g _24976_ (.A(reg_out[12]), .B(_12542_), .Y(_03789_));
NAND_g _24977_ (.A(_12611_), .B(_03789_), .Y(_03790_));
NAND_g _24978_ (.A(_02594_), .B(_03790_), .Y(_03791_));
NAND_g _24979_ (.A(pcpi_rs1[12]), .B(_02593_), .Y(_03792_));
NAND_g _24980_ (.A(_03791_), .B(_03792_), .Y(mem_la_addr[12]));
NAND_g _24981_ (.A(_02602_), .B(mem_la_addr[12]), .Y(_03793_));
NAND_g _24982_ (.A(mem_addr[12]), .B(_02603_), .Y(_03794_));
NAND_g _24983_ (.A(_03793_), .B(_03794_), .Y(_00814_));
NAND_g _24984_ (.A(reg_out[13]), .B(_12542_), .Y(_03795_));
NAND_g _24985_ (.A(_12617_), .B(_03795_), .Y(_03796_));
NAND_g _24986_ (.A(_02594_), .B(_03796_), .Y(_03797_));
NAND_g _24987_ (.A(pcpi_rs1[13]), .B(_02593_), .Y(_03798_));
NAND_g _24988_ (.A(_03797_), .B(_03798_), .Y(mem_la_addr[13]));
NAND_g _24989_ (.A(_02602_), .B(mem_la_addr[13]), .Y(_03799_));
NAND_g _24990_ (.A(mem_addr[13]), .B(_02603_), .Y(_03800_));
NAND_g _24991_ (.A(_03799_), .B(_03800_), .Y(_00815_));
NAND_g _24992_ (.A(reg_out[14]), .B(_12542_), .Y(_03801_));
NAND_g _24993_ (.A(_12623_), .B(_03801_), .Y(_03802_));
NAND_g _24994_ (.A(_02594_), .B(_03802_), .Y(_03803_));
NAND_g _24995_ (.A(pcpi_rs1[14]), .B(_02593_), .Y(_03804_));
NAND_g _24996_ (.A(_03803_), .B(_03804_), .Y(mem_la_addr[14]));
NAND_g _24997_ (.A(mem_addr[14]), .B(_02603_), .Y(_03805_));
NAND_g _24998_ (.A(_02602_), .B(mem_la_addr[14]), .Y(_03806_));
NAND_g _24999_ (.A(_03805_), .B(_03806_), .Y(_00816_));
NAND_g _25000_ (.A(reg_out[15]), .B(_12542_), .Y(_03807_));
NAND_g _25001_ (.A(_12629_), .B(_03807_), .Y(_03808_));
NAND_g _25002_ (.A(_02594_), .B(_03808_), .Y(_03809_));
NAND_g _25003_ (.A(pcpi_rs1[15]), .B(_02593_), .Y(_03810_));
NAND_g _25004_ (.A(_03809_), .B(_03810_), .Y(mem_la_addr[15]));
NAND_g _25005_ (.A(_02602_), .B(mem_la_addr[15]), .Y(_03811_));
NAND_g _25006_ (.A(mem_addr[15]), .B(_02603_), .Y(_03812_));
NAND_g _25007_ (.A(_03811_), .B(_03812_), .Y(_00817_));
NAND_g _25008_ (.A(reg_out[16]), .B(_12542_), .Y(_03813_));
NAND_g _25009_ (.A(_12635_), .B(_03813_), .Y(_03814_));
NAND_g _25010_ (.A(_02594_), .B(_03814_), .Y(_03815_));
NAND_g _25011_ (.A(pcpi_rs1[16]), .B(_02593_), .Y(_03816_));
NAND_g _25012_ (.A(_03815_), .B(_03816_), .Y(mem_la_addr[16]));
NAND_g _25013_ (.A(_02602_), .B(mem_la_addr[16]), .Y(_03817_));
NAND_g _25014_ (.A(mem_addr[16]), .B(_02603_), .Y(_03818_));
NAND_g _25015_ (.A(_03817_), .B(_03818_), .Y(_00818_));
NAND_g _25016_ (.A(reg_out[17]), .B(_12542_), .Y(_03819_));
NAND_g _25017_ (.A(_12641_), .B(_03819_), .Y(_03820_));
NAND_g _25018_ (.A(_02594_), .B(_03820_), .Y(_03821_));
NAND_g _25019_ (.A(pcpi_rs1[17]), .B(_02593_), .Y(_03822_));
NAND_g _25020_ (.A(_03821_), .B(_03822_), .Y(mem_la_addr[17]));
NAND_g _25021_ (.A(_02602_), .B(mem_la_addr[17]), .Y(_03823_));
NAND_g _25022_ (.A(mem_addr[17]), .B(_02603_), .Y(_03824_));
NAND_g _25023_ (.A(_03823_), .B(_03824_), .Y(_00819_));
NAND_g _25024_ (.A(reg_out[18]), .B(_12542_), .Y(_03825_));
NAND_g _25025_ (.A(_12647_), .B(_03825_), .Y(_03826_));
NAND_g _25026_ (.A(_02594_), .B(_03826_), .Y(_03827_));
NAND_g _25027_ (.A(pcpi_rs1[18]), .B(_02593_), .Y(_03828_));
NAND_g _25028_ (.A(_03827_), .B(_03828_), .Y(mem_la_addr[18]));
NAND_g _25029_ (.A(_02602_), .B(mem_la_addr[18]), .Y(_03829_));
NAND_g _25030_ (.A(mem_addr[18]), .B(_02603_), .Y(_03830_));
NAND_g _25031_ (.A(_03829_), .B(_03830_), .Y(_00820_));
NAND_g _25032_ (.A(reg_out[19]), .B(_12542_), .Y(_03831_));
NAND_g _25033_ (.A(_12653_), .B(_03831_), .Y(_03832_));
NAND_g _25034_ (.A(_02594_), .B(_03832_), .Y(_03833_));
NAND_g _25035_ (.A(pcpi_rs1[19]), .B(_02593_), .Y(_03834_));
NAND_g _25036_ (.A(_03833_), .B(_03834_), .Y(mem_la_addr[19]));
NAND_g _25037_ (.A(_02602_), .B(mem_la_addr[19]), .Y(_03835_));
NAND_g _25038_ (.A(mem_addr[19]), .B(_02603_), .Y(_03836_));
NAND_g _25039_ (.A(_03835_), .B(_03836_), .Y(_00821_));
NAND_g _25040_ (.A(reg_out[20]), .B(_12542_), .Y(_03837_));
NAND_g _25041_ (.A(_12659_), .B(_03837_), .Y(_03838_));
NAND_g _25042_ (.A(_02594_), .B(_03838_), .Y(_03839_));
NAND_g _25043_ (.A(pcpi_rs1[20]), .B(_02593_), .Y(_03840_));
NAND_g _25044_ (.A(_03839_), .B(_03840_), .Y(mem_la_addr[20]));
NAND_g _25045_ (.A(_02602_), .B(mem_la_addr[20]), .Y(_03841_));
NAND_g _25046_ (.A(mem_addr[20]), .B(_02603_), .Y(_03842_));
NAND_g _25047_ (.A(_03841_), .B(_03842_), .Y(_00822_));
NAND_g _25048_ (.A(reg_out[21]), .B(_12542_), .Y(_03843_));
NAND_g _25049_ (.A(_12665_), .B(_03843_), .Y(_03844_));
NAND_g _25050_ (.A(_02594_), .B(_03844_), .Y(_03845_));
NAND_g _25051_ (.A(pcpi_rs1[21]), .B(_02593_), .Y(_03846_));
NAND_g _25052_ (.A(_03845_), .B(_03846_), .Y(mem_la_addr[21]));
NAND_g _25053_ (.A(_02602_), .B(mem_la_addr[21]), .Y(_03847_));
NAND_g _25054_ (.A(mem_addr[21]), .B(_02603_), .Y(_03848_));
NAND_g _25055_ (.A(_03847_), .B(_03848_), .Y(_00823_));
NAND_g _25056_ (.A(reg_out[22]), .B(_12542_), .Y(_03849_));
NAND_g _25057_ (.A(_12671_), .B(_03849_), .Y(_03850_));
NAND_g _25058_ (.A(_02594_), .B(_03850_), .Y(_03851_));
NAND_g _25059_ (.A(pcpi_rs1[22]), .B(_02593_), .Y(_03852_));
NAND_g _25060_ (.A(_03851_), .B(_03852_), .Y(mem_la_addr[22]));
NAND_g _25061_ (.A(_02602_), .B(mem_la_addr[22]), .Y(_03853_));
NAND_g _25062_ (.A(mem_addr[22]), .B(_02603_), .Y(_03854_));
NAND_g _25063_ (.A(_03853_), .B(_03854_), .Y(_00824_));
NAND_g _25064_ (.A(reg_out[23]), .B(_12542_), .Y(_03855_));
NAND_g _25065_ (.A(_12677_), .B(_03855_), .Y(_03856_));
NAND_g _25066_ (.A(_02594_), .B(_03856_), .Y(_03857_));
NAND_g _25067_ (.A(pcpi_rs1[23]), .B(_02593_), .Y(_03858_));
NAND_g _25068_ (.A(_03857_), .B(_03858_), .Y(mem_la_addr[23]));
NAND_g _25069_ (.A(mem_addr[23]), .B(_02603_), .Y(_03859_));
NAND_g _25070_ (.A(_02602_), .B(mem_la_addr[23]), .Y(_03860_));
NAND_g _25071_ (.A(_03859_), .B(_03860_), .Y(_00825_));
NAND_g _25072_ (.A(reg_out[24]), .B(_12542_), .Y(_03861_));
NAND_g _25073_ (.A(_12682_), .B(_03861_), .Y(_03862_));
NAND_g _25074_ (.A(_02594_), .B(_03862_), .Y(_03863_));
NAND_g _25075_ (.A(pcpi_rs1[24]), .B(_02593_), .Y(_03864_));
NAND_g _25076_ (.A(_03863_), .B(_03864_), .Y(mem_la_addr[24]));
NAND_g _25077_ (.A(_02602_), .B(mem_la_addr[24]), .Y(_03865_));
NAND_g _25078_ (.A(mem_addr[24]), .B(_02603_), .Y(_03866_));
NAND_g _25079_ (.A(_03865_), .B(_03866_), .Y(_00826_));
NAND_g _25080_ (.A(reg_out[25]), .B(_12542_), .Y(_03867_));
NAND_g _25081_ (.A(_12688_), .B(_03867_), .Y(_03868_));
NAND_g _25082_ (.A(_02594_), .B(_03868_), .Y(_03869_));
NAND_g _25083_ (.A(pcpi_rs1[25]), .B(_02593_), .Y(_03870_));
NAND_g _25084_ (.A(_03869_), .B(_03870_), .Y(mem_la_addr[25]));
NAND_g _25085_ (.A(_02602_), .B(mem_la_addr[25]), .Y(_03871_));
NAND_g _25086_ (.A(mem_addr[25]), .B(_02603_), .Y(_03872_));
NAND_g _25087_ (.A(_03871_), .B(_03872_), .Y(_00827_));
NAND_g _25088_ (.A(reg_out[26]), .B(_12542_), .Y(_03873_));
NAND_g _25089_ (.A(_12693_), .B(_03873_), .Y(_03874_));
NAND_g _25090_ (.A(_02594_), .B(_03874_), .Y(_03875_));
NAND_g _25091_ (.A(pcpi_rs1[26]), .B(_02593_), .Y(_03876_));
NAND_g _25092_ (.A(_03875_), .B(_03876_), .Y(mem_la_addr[26]));
NAND_g _25093_ (.A(mem_addr[26]), .B(_02603_), .Y(_03877_));
NAND_g _25094_ (.A(_02602_), .B(mem_la_addr[26]), .Y(_03878_));
NAND_g _25095_ (.A(_03877_), .B(_03878_), .Y(_00828_));
NAND_g _25096_ (.A(reg_out[27]), .B(_12542_), .Y(_03879_));
NAND_g _25097_ (.A(_12699_), .B(_03879_), .Y(_03880_));
NAND_g _25098_ (.A(_02594_), .B(_03880_), .Y(_03881_));
NAND_g _25099_ (.A(pcpi_rs1[27]), .B(_02593_), .Y(_03882_));
NAND_g _25100_ (.A(_03881_), .B(_03882_), .Y(mem_la_addr[27]));
NAND_g _25101_ (.A(mem_addr[27]), .B(_02603_), .Y(_03883_));
NAND_g _25102_ (.A(_02602_), .B(mem_la_addr[27]), .Y(_03884_));
NAND_g _25103_ (.A(_03883_), .B(_03884_), .Y(_00829_));
NAND_g _25104_ (.A(reg_out[28]), .B(_12542_), .Y(_03885_));
NAND_g _25105_ (.A(_12704_), .B(_03885_), .Y(_03886_));
NAND_g _25106_ (.A(_02594_), .B(_03886_), .Y(_03887_));
NAND_g _25107_ (.A(pcpi_rs1[28]), .B(_02593_), .Y(_03888_));
NAND_g _25108_ (.A(_03887_), .B(_03888_), .Y(mem_la_addr[28]));
NAND_g _25109_ (.A(_02602_), .B(mem_la_addr[28]), .Y(_03889_));
NAND_g _25110_ (.A(mem_addr[28]), .B(_02603_), .Y(_03890_));
NAND_g _25111_ (.A(_03889_), .B(_03890_), .Y(_00830_));
NAND_g _25112_ (.A(reg_out[29]), .B(_12542_), .Y(_03891_));
NAND_g _25113_ (.A(_12710_), .B(_03891_), .Y(_03892_));
NAND_g _25114_ (.A(_02594_), .B(_03892_), .Y(_03893_));
NAND_g _25115_ (.A(pcpi_rs1[29]), .B(_02593_), .Y(_03894_));
NAND_g _25116_ (.A(_03893_), .B(_03894_), .Y(mem_la_addr[29]));
NAND_g _25117_ (.A(_02602_), .B(mem_la_addr[29]), .Y(_03895_));
NAND_g _25118_ (.A(mem_addr[29]), .B(_02603_), .Y(_03896_));
NAND_g _25119_ (.A(_03895_), .B(_03896_), .Y(_00831_));
NAND_g _25120_ (.A(reg_out[30]), .B(_12542_), .Y(_03897_));
NAND_g _25121_ (.A(_12716_), .B(_03897_), .Y(_03898_));
NAND_g _25122_ (.A(_02594_), .B(_03898_), .Y(_03899_));
NAND_g _25123_ (.A(pcpi_rs1[30]), .B(_02593_), .Y(_03900_));
NAND_g _25124_ (.A(_03899_), .B(_03900_), .Y(mem_la_addr[30]));
NAND_g _25125_ (.A(_02602_), .B(mem_la_addr[30]), .Y(_03901_));
NAND_g _25126_ (.A(mem_addr[30]), .B(_02603_), .Y(_03902_));
NAND_g _25127_ (.A(_03901_), .B(_03902_), .Y(_00832_));
NAND_g _25128_ (.A(reg_out[31]), .B(_12542_), .Y(_03903_));
NAND_g _25129_ (.A(_12721_), .B(_03903_), .Y(_03904_));
NAND_g _25130_ (.A(_02594_), .B(_03904_), .Y(_03905_));
NAND_g _25131_ (.A(pcpi_rs1[31]), .B(_02593_), .Y(_03906_));
NAND_g _25132_ (.A(_03905_), .B(_03906_), .Y(mem_la_addr[31]));
NAND_g _25133_ (.A(_02602_), .B(mem_la_addr[31]), .Y(_03907_));
NAND_g _25134_ (.A(mem_addr[31]), .B(_02603_), .Y(_03908_));
NAND_g _25135_ (.A(_03907_), .B(_03908_), .Y(_00833_));
NAND_g _25136_ (.A(mem_wordsize[0]), .B(mem_wordsize[1]), .Y(_03909_));
AND_g _25137_ (.A(pcpi_rs2[0]), .B(_03909_), .Y(mem_la_wdata[0]));
AND_g _25138_ (.A(_02598_), .B(_02600_), .Y(_03910_));
NAND_g _25139_ (.A(_02598_), .B(_02600_), .Y(_03911_));
NAND_g _25140_ (.A(mem_la_wdata[0]), .B(_03910_), .Y(_03912_));
NAND_g _25141_ (.A(mem_wdata[0]), .B(_03911_), .Y(_03913_));
NAND_g _25142_ (.A(_03912_), .B(_03913_), .Y(_00834_));
AND_g _25143_ (.A(pcpi_rs2[1]), .B(_03909_), .Y(mem_la_wdata[1]));
NAND_g _25144_ (.A(_03910_), .B(mem_la_wdata[1]), .Y(_03914_));
NAND_g _25145_ (.A(mem_wdata[1]), .B(_03911_), .Y(_03915_));
NAND_g _25146_ (.A(_03914_), .B(_03915_), .Y(_00835_));
AND_g _25147_ (.A(pcpi_rs2[2]), .B(_03909_), .Y(mem_la_wdata[2]));
NAND_g _25148_ (.A(_03910_), .B(mem_la_wdata[2]), .Y(_03916_));
NAND_g _25149_ (.A(mem_wdata[2]), .B(_03911_), .Y(_03917_));
NAND_g _25150_ (.A(_03916_), .B(_03917_), .Y(_00836_));
AND_g _25151_ (.A(pcpi_rs2[3]), .B(_03909_), .Y(mem_la_wdata[3]));
NAND_g _25152_ (.A(_03910_), .B(mem_la_wdata[3]), .Y(_03918_));
NAND_g _25153_ (.A(mem_wdata[3]), .B(_03911_), .Y(_03919_));
NAND_g _25154_ (.A(_03918_), .B(_03919_), .Y(_00837_));
AND_g _25155_ (.A(pcpi_rs2[4]), .B(_03909_), .Y(mem_la_wdata[4]));
NAND_g _25156_ (.A(_03910_), .B(mem_la_wdata[4]), .Y(_03920_));
NAND_g _25157_ (.A(mem_wdata[4]), .B(_03911_), .Y(_03921_));
NAND_g _25158_ (.A(_03920_), .B(_03921_), .Y(_00838_));
AND_g _25159_ (.A(pcpi_rs2[5]), .B(_03909_), .Y(mem_la_wdata[5]));
NAND_g _25160_ (.A(_03910_), .B(mem_la_wdata[5]), .Y(_03922_));
NAND_g _25161_ (.A(mem_wdata[5]), .B(_03911_), .Y(_03923_));
NAND_g _25162_ (.A(_03922_), .B(_03923_), .Y(_00839_));
AND_g _25163_ (.A(pcpi_rs2[6]), .B(_03909_), .Y(mem_la_wdata[6]));
NAND_g _25164_ (.A(_03910_), .B(mem_la_wdata[6]), .Y(_03924_));
NAND_g _25165_ (.A(mem_wdata[6]), .B(_03911_), .Y(_03925_));
NAND_g _25166_ (.A(_03924_), .B(_03925_), .Y(_00840_));
AND_g _25167_ (.A(pcpi_rs2[7]), .B(_03909_), .Y(mem_la_wdata[7]));
NAND_g _25168_ (.A(_03910_), .B(mem_la_wdata[7]), .Y(_03926_));
NAND_g _25169_ (.A(mem_wdata[7]), .B(_03911_), .Y(_03927_));
NAND_g _25170_ (.A(_03926_), .B(_03927_), .Y(_00841_));
AND_g _25171_ (.A(_11012_), .B(mem_wordsize[1]), .Y(_03928_));
NAND_g _25172_ (.A(pcpi_rs2[0]), .B(_03928_), .Y(_03929_));
NAND_g _25173_ (.A(pcpi_rs2[8]), .B(_11013_), .Y(_03930_));
NAND_g _25174_ (.A(_03929_), .B(_03930_), .Y(mem_la_wdata[8]));
NAND_g _25175_ (.A(mem_wdata[8]), .B(_03911_), .Y(_03931_));
NAND_g _25176_ (.A(_03910_), .B(mem_la_wdata[8]), .Y(_03932_));
NAND_g _25177_ (.A(_03931_), .B(_03932_), .Y(_00842_));
NAND_g _25178_ (.A(pcpi_rs2[1]), .B(_03928_), .Y(_03933_));
NAND_g _25179_ (.A(pcpi_rs2[9]), .B(_11013_), .Y(_03934_));
NAND_g _25180_ (.A(_03933_), .B(_03934_), .Y(mem_la_wdata[9]));
NAND_g _25181_ (.A(mem_wdata[9]), .B(_03911_), .Y(_03935_));
NAND_g _25182_ (.A(_03910_), .B(mem_la_wdata[9]), .Y(_03936_));
NAND_g _25183_ (.A(_03935_), .B(_03936_), .Y(_00843_));
NAND_g _25184_ (.A(pcpi_rs2[2]), .B(_03928_), .Y(_03937_));
NAND_g _25185_ (.A(pcpi_rs2[10]), .B(_11013_), .Y(_03938_));
NAND_g _25186_ (.A(_03937_), .B(_03938_), .Y(mem_la_wdata[10]));
NAND_g _25187_ (.A(mem_wdata[10]), .B(_03911_), .Y(_03939_));
NAND_g _25188_ (.A(_03910_), .B(mem_la_wdata[10]), .Y(_03940_));
NAND_g _25189_ (.A(_03939_), .B(_03940_), .Y(_00844_));
NAND_g _25190_ (.A(pcpi_rs2[3]), .B(_03928_), .Y(_03941_));
NAND_g _25191_ (.A(pcpi_rs2[11]), .B(_11013_), .Y(_03942_));
NAND_g _25192_ (.A(_03941_), .B(_03942_), .Y(mem_la_wdata[11]));
NAND_g _25193_ (.A(mem_wdata[11]), .B(_03911_), .Y(_03943_));
NAND_g _25194_ (.A(_03910_), .B(mem_la_wdata[11]), .Y(_03944_));
NAND_g _25195_ (.A(_03943_), .B(_03944_), .Y(_00845_));
NAND_g _25196_ (.A(pcpi_rs2[4]), .B(_03928_), .Y(_03945_));
NAND_g _25197_ (.A(pcpi_rs2[12]), .B(_11013_), .Y(_03946_));
NAND_g _25198_ (.A(_03945_), .B(_03946_), .Y(mem_la_wdata[12]));
NAND_g _25199_ (.A(mem_wdata[12]), .B(_03911_), .Y(_03947_));
NAND_g _25200_ (.A(_03910_), .B(mem_la_wdata[12]), .Y(_03948_));
NAND_g _25201_ (.A(_03947_), .B(_03948_), .Y(_00846_));
NAND_g _25202_ (.A(pcpi_rs2[5]), .B(_03928_), .Y(_03949_));
NAND_g _25203_ (.A(pcpi_rs2[13]), .B(_11013_), .Y(_03950_));
NAND_g _25204_ (.A(_03949_), .B(_03950_), .Y(mem_la_wdata[13]));
NAND_g _25205_ (.A(mem_wdata[13]), .B(_03911_), .Y(_03951_));
NAND_g _25206_ (.A(_03910_), .B(mem_la_wdata[13]), .Y(_03952_));
NAND_g _25207_ (.A(_03951_), .B(_03952_), .Y(_00847_));
NAND_g _25208_ (.A(pcpi_rs2[6]), .B(_03928_), .Y(_03953_));
NAND_g _25209_ (.A(pcpi_rs2[14]), .B(_11013_), .Y(_03954_));
NAND_g _25210_ (.A(_03953_), .B(_03954_), .Y(mem_la_wdata[14]));
NAND_g _25211_ (.A(mem_wdata[14]), .B(_03911_), .Y(_03955_));
NAND_g _25212_ (.A(_03910_), .B(mem_la_wdata[14]), .Y(_03956_));
NAND_g _25213_ (.A(_03955_), .B(_03956_), .Y(_00848_));
NAND_g _25214_ (.A(pcpi_rs2[7]), .B(_03928_), .Y(_03957_));
NAND_g _25215_ (.A(pcpi_rs2[15]), .B(_11013_), .Y(_03958_));
NAND_g _25216_ (.A(_03957_), .B(_03958_), .Y(mem_la_wdata[15]));
NAND_g _25217_ (.A(mem_wdata[15]), .B(_03911_), .Y(_03959_));
NAND_g _25218_ (.A(_03910_), .B(mem_la_wdata[15]), .Y(_03960_));
NAND_g _25219_ (.A(_03959_), .B(_03960_), .Y(_00849_));
NOR_g _25220_ (.A(mem_wordsize[0]), .B(mem_wordsize[1]), .Y(_03961_));
NAND_g _25221_ (.A(_11012_), .B(_11013_), .Y(_03962_));
NAND_g _25222_ (.A(pcpi_rs2[16]), .B(_03961_), .Y(_03963_));
NAND_g _25223_ (.A(mem_la_wdata[0]), .B(_03962_), .Y(_03964_));
NAND_g _25224_ (.A(_03963_), .B(_03964_), .Y(mem_la_wdata[16]));
NAND_g _25225_ (.A(_03910_), .B(mem_la_wdata[16]), .Y(_03965_));
NAND_g _25226_ (.A(mem_wdata[16]), .B(_03911_), .Y(_03966_));
NAND_g _25227_ (.A(_03965_), .B(_03966_), .Y(_00850_));
NAND_g _25228_ (.A(pcpi_rs2[17]), .B(_03961_), .Y(_03967_));
NAND_g _25229_ (.A(mem_la_wdata[1]), .B(_03962_), .Y(_03968_));
NAND_g _25230_ (.A(_03967_), .B(_03968_), .Y(mem_la_wdata[17]));
NAND_g _25231_ (.A(_03910_), .B(mem_la_wdata[17]), .Y(_03969_));
NAND_g _25232_ (.A(mem_wdata[17]), .B(_03911_), .Y(_03970_));
NAND_g _25233_ (.A(_03969_), .B(_03970_), .Y(_00851_));
NAND_g _25234_ (.A(pcpi_rs2[18]), .B(_03961_), .Y(_03971_));
NAND_g _25235_ (.A(mem_la_wdata[2]), .B(_03962_), .Y(_03972_));
NAND_g _25236_ (.A(_03971_), .B(_03972_), .Y(mem_la_wdata[18]));
NAND_g _25237_ (.A(_03910_), .B(mem_la_wdata[18]), .Y(_03973_));
NAND_g _25238_ (.A(mem_wdata[18]), .B(_03911_), .Y(_03974_));
NAND_g _25239_ (.A(_03973_), .B(_03974_), .Y(_00852_));
NAND_g _25240_ (.A(pcpi_rs2[19]), .B(_03961_), .Y(_03975_));
NAND_g _25241_ (.A(mem_la_wdata[3]), .B(_03962_), .Y(_03976_));
NAND_g _25242_ (.A(_03975_), .B(_03976_), .Y(mem_la_wdata[19]));
NAND_g _25243_ (.A(_03910_), .B(mem_la_wdata[19]), .Y(_03977_));
NAND_g _25244_ (.A(mem_wdata[19]), .B(_03911_), .Y(_03978_));
NAND_g _25245_ (.A(_03977_), .B(_03978_), .Y(_00853_));
NAND_g _25246_ (.A(pcpi_rs2[20]), .B(_03961_), .Y(_03979_));
NAND_g _25247_ (.A(mem_la_wdata[4]), .B(_03962_), .Y(_03980_));
NAND_g _25248_ (.A(_03979_), .B(_03980_), .Y(mem_la_wdata[20]));
NAND_g _25249_ (.A(_03910_), .B(mem_la_wdata[20]), .Y(_03981_));
NAND_g _25250_ (.A(mem_wdata[20]), .B(_03911_), .Y(_03982_));
NAND_g _25251_ (.A(_03981_), .B(_03982_), .Y(_00854_));
NAND_g _25252_ (.A(pcpi_rs2[21]), .B(_03961_), .Y(_03983_));
NAND_g _25253_ (.A(mem_la_wdata[5]), .B(_03962_), .Y(_03984_));
NAND_g _25254_ (.A(_03983_), .B(_03984_), .Y(mem_la_wdata[21]));
NAND_g _25255_ (.A(_03910_), .B(mem_la_wdata[21]), .Y(_03985_));
NAND_g _25256_ (.A(mem_wdata[21]), .B(_03911_), .Y(_03986_));
NAND_g _25257_ (.A(_03985_), .B(_03986_), .Y(_00855_));
NAND_g _25258_ (.A(pcpi_rs2[22]), .B(_03961_), .Y(_03987_));
NAND_g _25259_ (.A(mem_la_wdata[6]), .B(_03962_), .Y(_03988_));
NAND_g _25260_ (.A(_03987_), .B(_03988_), .Y(mem_la_wdata[22]));
NAND_g _25261_ (.A(_03910_), .B(mem_la_wdata[22]), .Y(_03989_));
NAND_g _25262_ (.A(mem_wdata[22]), .B(_03911_), .Y(_03990_));
NAND_g _25263_ (.A(_03989_), .B(_03990_), .Y(_00856_));
NAND_g _25264_ (.A(pcpi_rs2[23]), .B(_03961_), .Y(_03991_));
NAND_g _25265_ (.A(mem_la_wdata[7]), .B(_03962_), .Y(_03992_));
NAND_g _25266_ (.A(_03991_), .B(_03992_), .Y(mem_la_wdata[23]));
NAND_g _25267_ (.A(_03910_), .B(mem_la_wdata[23]), .Y(_03993_));
NAND_g _25268_ (.A(mem_wdata[23]), .B(_03911_), .Y(_03994_));
NAND_g _25269_ (.A(_03993_), .B(_03994_), .Y(_00857_));
NAND_g _25270_ (.A(pcpi_rs2[24]), .B(_03961_), .Y(_03995_));
AND_g _25271_ (.A(mem_wordsize[0]), .B(_11013_), .Y(_03996_));
NAND_g _25272_ (.A(pcpi_rs2[8]), .B(_03996_), .Y(_03997_));
AND_g _25273_ (.A(_03929_), .B(_03997_), .Y(_03998_));
NAND_g _25274_ (.A(_03995_), .B(_03998_), .Y(mem_la_wdata[24]));
NAND_g _25275_ (.A(mem_wdata[24]), .B(_03911_), .Y(_03999_));
NAND_g _25276_ (.A(_03910_), .B(mem_la_wdata[24]), .Y(_04000_));
NAND_g _25277_ (.A(_03999_), .B(_04000_), .Y(_00858_));
NAND_g _25278_ (.A(pcpi_rs2[25]), .B(_03961_), .Y(_04001_));
NAND_g _25279_ (.A(pcpi_rs2[9]), .B(_03996_), .Y(_04002_));
AND_g _25280_ (.A(_03933_), .B(_04002_), .Y(_04003_));
NAND_g _25281_ (.A(_04001_), .B(_04003_), .Y(mem_la_wdata[25]));
NAND_g _25282_ (.A(mem_wdata[25]), .B(_03911_), .Y(_04004_));
NAND_g _25283_ (.A(_03910_), .B(mem_la_wdata[25]), .Y(_04005_));
NAND_g _25284_ (.A(_04004_), .B(_04005_), .Y(_00859_));
NAND_g _25285_ (.A(pcpi_rs2[10]), .B(_03996_), .Y(_04006_));
NAND_g _25286_ (.A(pcpi_rs2[26]), .B(_03961_), .Y(_04007_));
AND_g _25287_ (.A(_03937_), .B(_04006_), .Y(_04008_));
NAND_g _25288_ (.A(_04007_), .B(_04008_), .Y(mem_la_wdata[26]));
NAND_g _25289_ (.A(mem_wdata[26]), .B(_03911_), .Y(_04009_));
NAND_g _25290_ (.A(_03910_), .B(mem_la_wdata[26]), .Y(_04010_));
NAND_g _25291_ (.A(_04009_), .B(_04010_), .Y(_00860_));
NAND_g _25292_ (.A(pcpi_rs2[27]), .B(_03961_), .Y(_04011_));
NAND_g _25293_ (.A(pcpi_rs2[11]), .B(_03996_), .Y(_04012_));
AND_g _25294_ (.A(_03941_), .B(_04012_), .Y(_04013_));
NAND_g _25295_ (.A(_04011_), .B(_04013_), .Y(mem_la_wdata[27]));
NAND_g _25296_ (.A(mem_wdata[27]), .B(_03911_), .Y(_04014_));
NAND_g _25297_ (.A(_03910_), .B(mem_la_wdata[27]), .Y(_04015_));
NAND_g _25298_ (.A(_04014_), .B(_04015_), .Y(_00861_));
NAND_g _25299_ (.A(pcpi_rs2[12]), .B(_03996_), .Y(_04016_));
NAND_g _25300_ (.A(pcpi_rs2[28]), .B(_03961_), .Y(_04017_));
AND_g _25301_ (.A(_03945_), .B(_04016_), .Y(_04018_));
NAND_g _25302_ (.A(_04017_), .B(_04018_), .Y(mem_la_wdata[28]));
NAND_g _25303_ (.A(mem_wdata[28]), .B(_03911_), .Y(_04019_));
NAND_g _25304_ (.A(_03910_), .B(mem_la_wdata[28]), .Y(_04020_));
NAND_g _25305_ (.A(_04019_), .B(_04020_), .Y(_00862_));
NAND_g _25306_ (.A(pcpi_rs2[13]), .B(_03996_), .Y(_04021_));
NAND_g _25307_ (.A(pcpi_rs2[29]), .B(_03961_), .Y(_04022_));
AND_g _25308_ (.A(_03949_), .B(_04021_), .Y(_04023_));
NAND_g _25309_ (.A(_04022_), .B(_04023_), .Y(mem_la_wdata[29]));
NAND_g _25310_ (.A(mem_wdata[29]), .B(_03911_), .Y(_04024_));
NAND_g _25311_ (.A(_03910_), .B(mem_la_wdata[29]), .Y(_04025_));
NAND_g _25312_ (.A(_04024_), .B(_04025_), .Y(_00863_));
NAND_g _25313_ (.A(pcpi_rs2[14]), .B(_03996_), .Y(_04026_));
NAND_g _25314_ (.A(pcpi_rs2[30]), .B(_03961_), .Y(_04027_));
AND_g _25315_ (.A(_03953_), .B(_04026_), .Y(_04028_));
NAND_g _25316_ (.A(_04027_), .B(_04028_), .Y(mem_la_wdata[30]));
NAND_g _25317_ (.A(mem_wdata[30]), .B(_03911_), .Y(_04029_));
NAND_g _25318_ (.A(_03910_), .B(mem_la_wdata[30]), .Y(_04030_));
NAND_g _25319_ (.A(_04029_), .B(_04030_), .Y(_00864_));
NAND_g _25320_ (.A(pcpi_rs2[15]), .B(_03996_), .Y(_04031_));
NAND_g _25321_ (.A(pcpi_rs2[31]), .B(_03961_), .Y(_04032_));
AND_g _25322_ (.A(_03957_), .B(_04031_), .Y(_04033_));
NAND_g _25323_ (.A(_04032_), .B(_04033_), .Y(mem_la_wdata[31]));
NAND_g _25324_ (.A(mem_wdata[31]), .B(_03911_), .Y(_04034_));
NAND_g _25325_ (.A(_03910_), .B(mem_la_wdata[31]), .Y(_04035_));
NAND_g _25326_ (.A(_04034_), .B(_04035_), .Y(_00865_));
NAND_g _25327_ (.A(mem_wstrb[0]), .B(_02603_), .Y(_04036_));
AND_g _25328_ (.A(mem_wordsize[0]), .B(pcpi_rs1[1]), .Y(_04037_));
NAND_g _25329_ (.A(mem_wordsize[0]), .B(pcpi_rs1[1]), .Y(_04038_));
AND_g _25330_ (.A(_11013_), .B(_04038_), .Y(_04039_));
NAND_g _25331_ (.A(_11013_), .B(_04038_), .Y(_04040_));
NOR_g _25332_ (.A(pcpi_rs1[0]), .B(pcpi_rs1[1]), .Y(_04041_));
NAND_g _25333_ (.A(_11012_), .B(_04041_), .Y(_04042_));
NAND_g _25334_ (.A(_04040_), .B(_04042_), .Y(mem_la_wstrb[0]));
NOR_g _25335_ (.A(_02601_), .B(_03911_), .Y(_04043_));
NAND_g _25336_ (.A(mem_la_wstrb[0]), .B(_04043_), .Y(_04044_));
NAND_g _25337_ (.A(_04036_), .B(_04044_), .Y(_00866_));
AND_g _25338_ (.A(pcpi_rs1[0]), .B(_11136_), .Y(_04045_));
NAND_g _25339_ (.A(_11012_), .B(_04045_), .Y(_04046_));
NAND_g _25340_ (.A(_04040_), .B(_04046_), .Y(mem_la_wstrb[1]));
NAND_g _25341_ (.A(_04043_), .B(mem_la_wstrb[1]), .Y(_04047_));
NAND_g _25342_ (.A(mem_wstrb[1]), .B(_02603_), .Y(_04048_));
NAND_g _25343_ (.A(_04047_), .B(_04048_), .Y(_00867_));
NAND_g _25344_ (.A(_11012_), .B(pcpi_rs1[1]), .Y(_04049_));
AND_g _25345_ (.A(pcpi_rs1[1]), .B(_03928_), .Y(_04050_));
NAND_g _25346_ (.A(_11135_), .B(_04050_), .Y(_04051_));
AND_g _25347_ (.A(_11013_), .B(_04037_), .Y(_04052_));
NAND_g _25348_ (.A(_11013_), .B(_04037_), .Y(_04053_));
NAND_g _25349_ (.A(_04051_), .B(_04053_), .Y(_04054_));
NOT_g _25350_ (.A(_04054_), .Y(_04055_));
NAND_g _25351_ (.A(_03962_), .B(_04055_), .Y(mem_la_wstrb[2]));
NAND_g _25352_ (.A(_04043_), .B(mem_la_wstrb[2]), .Y(_04056_));
NAND_g _25353_ (.A(mem_wstrb[2]), .B(_02603_), .Y(_04057_));
NAND_g _25354_ (.A(_04056_), .B(_04057_), .Y(_00868_));
NAND_g _25355_ (.A(mem_wstrb[3]), .B(_02603_), .Y(_04058_));
AND_g _25356_ (.A(pcpi_rs1[0]), .B(_04050_), .Y(_04059_));
NOR_g _25357_ (.A(_03961_), .B(_04059_), .Y(_04060_));
NAND_g _25358_ (.A(_04053_), .B(_04060_), .Y(mem_la_wstrb[3]));
NAND_g _25359_ (.A(_04043_), .B(mem_la_wstrb[3]), .Y(_04061_));
NAND_g _25360_ (.A(_04058_), .B(_04061_), .Y(_00869_));
NAND_g _25361_ (.A(_10898_), .B(_02611_), .Y(_04062_));
AND_g _25362_ (.A(_02609_), .B(_04062_), .Y(_04063_));
NAND_g _25363_ (.A(_02608_), .B(_04063_), .Y(_04064_));
NAND_g _25364_ (.A(mem_state[0]), .B(_04064_), .Y(_04065_));
AND_g _25365_ (.A(mem_state[0]), .B(_11084_), .Y(_04066_));
AND_g _25366_ (.A(_11908_), .B(_04066_), .Y(_04067_));
AND_g _25367_ (.A(_11910_), .B(_02598_), .Y(_04068_));
NAND_g _25368_ (.A(_04067_), .B(_04068_), .Y(_04069_));
NAND_g _25369_ (.A(_02595_), .B(_03707_), .Y(_04070_));
AND_g _25370_ (.A(_04069_), .B(_04070_), .Y(_04071_));
NAND_g _25371_ (.A(_04065_), .B(_04071_), .Y(_00870_));
NAND_g _25372_ (.A(mem_state[1]), .B(_04064_), .Y(_04072_));
AND_g _25373_ (.A(_03911_), .B(_04069_), .Y(_04073_));
NAND_g _25374_ (.A(_04072_), .B(_04073_), .Y(_00871_));
NAND_g _25375_ (.A(_11262_), .B(_12542_), .Y(_04074_));
AND_g _25376_ (.A(reg_next_pc[0]), .B(resetn), .Y(_04075_));
AND_g _25377_ (.A(_04074_), .B(_04075_), .Y(_00879_));
NOR_g _25378_ (.A(decoded_imm[31]), .B(_12314_), .Y(_04076_));
NAND_g _25379_ (.A(mem_rdata_q[31]), .B(_12520_), .Y(_04077_));
NAND_g _25380_ (.A(mem_rdata_q[31]), .B(_12484_), .Y(_04078_));
AND_g _25381_ (.A(_12314_), .B(_04078_), .Y(_04079_));
NAND_g _25382_ (.A(instr_jal), .B(decoded_imm_j[31]), .Y(_04080_));
NOR_g _25383_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(is_sb_sh_sw), .Y(_04081_));
NAND_g _25384_ (.A(_10902_), .B(_10980_), .Y(_04082_));
NAND_g _25385_ (.A(mem_rdata_q[31]), .B(_04082_), .Y(_04083_));
AND_g _25386_ (.A(_04080_), .B(_04083_), .Y(_04084_));
AND_g _25387_ (.A(_04079_), .B(_04084_), .Y(_04085_));
AND_g _25388_ (.A(_04077_), .B(_04085_), .Y(_04086_));
NOR_g _25389_ (.A(_04076_), .B(_04086_), .Y(_00880_));
NOR_g _25390_ (.A(decoded_imm[30]), .B(_12314_), .Y(_04087_));
NAND_g _25391_ (.A(mem_rdata_q[30]), .B(_12520_), .Y(_04088_));
AND_g _25392_ (.A(_04085_), .B(_04088_), .Y(_04089_));
NOR_g _25393_ (.A(_04087_), .B(_04089_), .Y(_00881_));
NOR_g _25394_ (.A(decoded_imm[29]), .B(_12314_), .Y(_04090_));
NAND_g _25395_ (.A(mem_rdata_q[29]), .B(_12520_), .Y(_04091_));
AND_g _25396_ (.A(_04085_), .B(_04091_), .Y(_04092_));
NOR_g _25397_ (.A(_04090_), .B(_04092_), .Y(_00882_));
NOR_g _25398_ (.A(decoded_imm[28]), .B(_12314_), .Y(_04093_));
NAND_g _25399_ (.A(mem_rdata_q[28]), .B(_12520_), .Y(_04094_));
AND_g _25400_ (.A(_04085_), .B(_04094_), .Y(_04095_));
NOR_g _25401_ (.A(_04093_), .B(_04095_), .Y(_00883_));
NOR_g _25402_ (.A(decoded_imm[27]), .B(_12314_), .Y(_04096_));
NAND_g _25403_ (.A(mem_rdata_q[27]), .B(_12520_), .Y(_04097_));
AND_g _25404_ (.A(_04085_), .B(_04097_), .Y(_04098_));
NOR_g _25405_ (.A(_04096_), .B(_04098_), .Y(_00884_));
NOR_g _25406_ (.A(decoded_imm[26]), .B(_12314_), .Y(_04099_));
NAND_g _25407_ (.A(mem_rdata_q[26]), .B(_12520_), .Y(_04100_));
AND_g _25408_ (.A(_04085_), .B(_04100_), .Y(_04101_));
NOR_g _25409_ (.A(_04099_), .B(_04101_), .Y(_00885_));
NOR_g _25410_ (.A(decoded_imm[25]), .B(_12314_), .Y(_04102_));
NAND_g _25411_ (.A(mem_rdata_q[25]), .B(_12520_), .Y(_04103_));
AND_g _25412_ (.A(_04085_), .B(_04103_), .Y(_04104_));
NOR_g _25413_ (.A(_04102_), .B(_04104_), .Y(_00886_));
NOR_g _25414_ (.A(decoded_imm[24]), .B(_12314_), .Y(_04105_));
NAND_g _25415_ (.A(mem_rdata_q[24]), .B(_12520_), .Y(_04106_));
AND_g _25416_ (.A(_04085_), .B(_04106_), .Y(_04107_));
NOR_g _25417_ (.A(_04105_), .B(_04107_), .Y(_00887_));
NOR_g _25418_ (.A(decoded_imm[23]), .B(_12314_), .Y(_04108_));
NAND_g _25419_ (.A(mem_rdata_q[23]), .B(_12520_), .Y(_04109_));
AND_g _25420_ (.A(_04085_), .B(_04109_), .Y(_04110_));
NOR_g _25421_ (.A(_04108_), .B(_04110_), .Y(_00888_));
NOR_g _25422_ (.A(decoded_imm[22]), .B(_12314_), .Y(_04111_));
NAND_g _25423_ (.A(mem_rdata_q[22]), .B(_12520_), .Y(_04112_));
AND_g _25424_ (.A(_04085_), .B(_04112_), .Y(_04113_));
NOR_g _25425_ (.A(_04111_), .B(_04113_), .Y(_00889_));
NOR_g _25426_ (.A(decoded_imm[21]), .B(_12314_), .Y(_04114_));
NAND_g _25427_ (.A(mem_rdata_q[21]), .B(_12520_), .Y(_04115_));
AND_g _25428_ (.A(_04085_), .B(_04115_), .Y(_04116_));
NOR_g _25429_ (.A(_04114_), .B(_04116_), .Y(_00890_));
NOR_g _25430_ (.A(decoded_imm[20]), .B(_12314_), .Y(_04117_));
NAND_g _25431_ (.A(mem_rdata_q[20]), .B(_12520_), .Y(_04118_));
AND_g _25432_ (.A(_04085_), .B(_04118_), .Y(_04119_));
NOR_g _25433_ (.A(_04117_), .B(_04119_), .Y(_00891_));
NOR_g _25434_ (.A(decoded_imm[19]), .B(_12314_), .Y(_04120_));
AND_g _25435_ (.A(_04079_), .B(_04083_), .Y(_04121_));
NAND_g _25436_ (.A(mem_rdata_q[19]), .B(_12520_), .Y(_04122_));
NAND_g _25437_ (.A(instr_jal), .B(decoded_imm_j[19]), .Y(_04123_));
AND_g _25438_ (.A(_04122_), .B(_04123_), .Y(_04124_));
AND_g _25439_ (.A(_04121_), .B(_04124_), .Y(_04125_));
NOR_g _25440_ (.A(_04120_), .B(_04125_), .Y(_00892_));
NOR_g _25441_ (.A(decoded_imm[18]), .B(_12314_), .Y(_04126_));
NAND_g _25442_ (.A(instr_jal), .B(decoded_imm_j[18]), .Y(_04127_));
NAND_g _25443_ (.A(mem_rdata_q[18]), .B(_12520_), .Y(_04128_));
AND_g _25444_ (.A(_04127_), .B(_04128_), .Y(_04129_));
AND_g _25445_ (.A(_04121_), .B(_04129_), .Y(_04130_));
NOR_g _25446_ (.A(_04126_), .B(_04130_), .Y(_00893_));
NOR_g _25447_ (.A(decoded_imm[17]), .B(_12314_), .Y(_04131_));
NAND_g _25448_ (.A(mem_rdata_q[17]), .B(_12520_), .Y(_04132_));
NAND_g _25449_ (.A(instr_jal), .B(decoded_imm_j[17]), .Y(_04133_));
AND_g _25450_ (.A(_04132_), .B(_04133_), .Y(_04134_));
AND_g _25451_ (.A(_04121_), .B(_04134_), .Y(_04135_));
NOR_g _25452_ (.A(_04131_), .B(_04135_), .Y(_00894_));
NOR_g _25453_ (.A(decoded_imm[16]), .B(_12314_), .Y(_04136_));
NAND_g _25454_ (.A(mem_rdata_q[16]), .B(_12520_), .Y(_04137_));
NAND_g _25455_ (.A(instr_jal), .B(decoded_imm_j[16]), .Y(_04138_));
AND_g _25456_ (.A(_04137_), .B(_04138_), .Y(_04139_));
AND_g _25457_ (.A(_04121_), .B(_04139_), .Y(_04140_));
NOR_g _25458_ (.A(_04136_), .B(_04140_), .Y(_00895_));
NOR_g _25459_ (.A(decoded_imm[15]), .B(_12314_), .Y(_04141_));
NAND_g _25460_ (.A(mem_rdata_q[15]), .B(_12520_), .Y(_04142_));
NAND_g _25461_ (.A(instr_jal), .B(decoded_imm_j[15]), .Y(_04143_));
AND_g _25462_ (.A(_04142_), .B(_04143_), .Y(_04144_));
AND_g _25463_ (.A(_04121_), .B(_04144_), .Y(_04145_));
NOR_g _25464_ (.A(_04141_), .B(_04145_), .Y(_00896_));
NOR_g _25465_ (.A(decoded_imm[14]), .B(_12314_), .Y(_04146_));
NOR_g _25466_ (.A(_11079_), .B(_12519_), .Y(_04147_));
AND_g _25467_ (.A(instr_jal), .B(decoded_imm_j[14]), .Y(_04148_));
NOR_g _25468_ (.A(_04147_), .B(_04148_), .Y(_04149_));
AND_g _25469_ (.A(_04121_), .B(_04149_), .Y(_04150_));
NOR_g _25470_ (.A(_04146_), .B(_04150_), .Y(_00897_));
NOR_g _25471_ (.A(decoded_imm[13]), .B(_12314_), .Y(_04151_));
AND_g _25472_ (.A(instr_jal), .B(decoded_imm_j[13]), .Y(_04152_));
NOR_g _25473_ (.A(_11078_), .B(_12519_), .Y(_04153_));
NOR_g _25474_ (.A(_04152_), .B(_04153_), .Y(_04154_));
AND_g _25475_ (.A(_04121_), .B(_04154_), .Y(_04155_));
NOR_g _25476_ (.A(_04151_), .B(_04155_), .Y(_00898_));
NOR_g _25477_ (.A(decoded_imm[12]), .B(_12314_), .Y(_04156_));
NOR_g _25478_ (.A(_11077_), .B(_12519_), .Y(_04157_));
AND_g _25479_ (.A(instr_jal), .B(decoded_imm_j[12]), .Y(_04158_));
NOR_g _25480_ (.A(_04157_), .B(_04158_), .Y(_04159_));
AND_g _25481_ (.A(_04121_), .B(_04159_), .Y(_04160_));
NOR_g _25482_ (.A(_04156_), .B(_04160_), .Y(_00899_));
NOR_g _25483_ (.A(decoded_imm[11]), .B(_12314_), .Y(_04161_));
NAND_g _25484_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(mem_rdata_q[7]), .Y(_04162_));
NAND_g _25485_ (.A(is_sb_sh_sw), .B(mem_rdata_q[31]), .Y(_04163_));
NAND_g _25486_ (.A(instr_jal), .B(decoded_imm_j[11]), .Y(_04164_));
AND_g _25487_ (.A(_04163_), .B(_04164_), .Y(_04165_));
AND_g _25488_ (.A(_04162_), .B(_04165_), .Y(_04166_));
AND_g _25489_ (.A(_04079_), .B(_04166_), .Y(_04167_));
NOR_g _25490_ (.A(_04161_), .B(_04167_), .Y(_00900_));
NAND_g _25491_ (.A(_12485_), .B(_04081_), .Y(_04168_));
NAND_g _25492_ (.A(mem_rdata_q[30]), .B(_04168_), .Y(_04169_));
NAND_g _25493_ (.A(instr_jal), .B(decoded_imm_j[10]), .Y(_04170_));
NOR_g _25494_ (.A(decoded_imm[10]), .B(_12314_), .Y(_04171_));
AND_g _25495_ (.A(_12314_), .B(_04170_), .Y(_04172_));
AND_g _25496_ (.A(_04169_), .B(_04172_), .Y(_04173_));
NOR_g _25497_ (.A(_04171_), .B(_04173_), .Y(_00901_));
NAND_g _25498_ (.A(mem_rdata_q[29]), .B(_04168_), .Y(_04174_));
NAND_g _25499_ (.A(decoded_imm_j[9]), .B(instr_jal), .Y(_04175_));
NOR_g _25500_ (.A(decoded_imm[9]), .B(_12314_), .Y(_04176_));
AND_g _25501_ (.A(_12314_), .B(_04175_), .Y(_04177_));
AND_g _25502_ (.A(_04174_), .B(_04177_), .Y(_04178_));
NOR_g _25503_ (.A(_04176_), .B(_04178_), .Y(_00902_));
NAND_g _25504_ (.A(mem_rdata_q[28]), .B(_04168_), .Y(_04179_));
NAND_g _25505_ (.A(decoded_imm_j[8]), .B(instr_jal), .Y(_04180_));
NOR_g _25506_ (.A(decoded_imm[8]), .B(_12314_), .Y(_04181_));
AND_g _25507_ (.A(_12314_), .B(_04180_), .Y(_04182_));
AND_g _25508_ (.A(_04179_), .B(_04182_), .Y(_04183_));
NOR_g _25509_ (.A(_04181_), .B(_04183_), .Y(_00903_));
NAND_g _25510_ (.A(mem_rdata_q[27]), .B(_04168_), .Y(_04184_));
NAND_g _25511_ (.A(instr_jal), .B(decoded_imm_j[7]), .Y(_04185_));
NOR_g _25512_ (.A(decoded_imm[7]), .B(_12314_), .Y(_04186_));
AND_g _25513_ (.A(_12314_), .B(_04185_), .Y(_04187_));
AND_g _25514_ (.A(_04184_), .B(_04187_), .Y(_04188_));
NOR_g _25515_ (.A(_04186_), .B(_04188_), .Y(_00904_));
NAND_g _25516_ (.A(mem_rdata_q[26]), .B(_04168_), .Y(_04189_));
NAND_g _25517_ (.A(instr_jal), .B(decoded_imm_j[6]), .Y(_04190_));
NOR_g _25518_ (.A(decoded_imm[6]), .B(_12314_), .Y(_04191_));
AND_g _25519_ (.A(_12314_), .B(_04190_), .Y(_04192_));
AND_g _25520_ (.A(_04189_), .B(_04192_), .Y(_04193_));
NOR_g _25521_ (.A(_04191_), .B(_04193_), .Y(_00905_));
NAND_g _25522_ (.A(mem_rdata_q[25]), .B(_04168_), .Y(_04194_));
NAND_g _25523_ (.A(decoded_imm_j[5]), .B(instr_jal), .Y(_04195_));
NOR_g _25524_ (.A(decoded_imm[5]), .B(_12314_), .Y(_04196_));
AND_g _25525_ (.A(_12314_), .B(_04195_), .Y(_04197_));
AND_g _25526_ (.A(_04194_), .B(_04197_), .Y(_04198_));
NOR_g _25527_ (.A(_04196_), .B(_04198_), .Y(_00906_));
NAND_g _25528_ (.A(mem_rdata_q[24]), .B(_12484_), .Y(_04199_));
NAND_g _25529_ (.A(mem_rdata_q[11]), .B(_04082_), .Y(_04200_));
NAND_g _25530_ (.A(instr_jal), .B(decoded_imm_j[4]), .Y(_04201_));
AND_g _25531_ (.A(_04200_), .B(_04201_), .Y(_04202_));
NAND_g _25532_ (.A(_04199_), .B(_04202_), .Y(_04203_));
NAND_g _25533_ (.A(_12314_), .B(_04203_), .Y(_04204_));
NAND_g _25534_ (.A(decoded_imm[4]), .B(_12315_), .Y(_04205_));
NAND_g _25535_ (.A(_04204_), .B(_04205_), .Y(_00907_));
NAND_g _25536_ (.A(mem_rdata_q[23]), .B(_12484_), .Y(_04206_));
NAND_g _25537_ (.A(mem_rdata_q[10]), .B(_04082_), .Y(_04207_));
NAND_g _25538_ (.A(instr_jal), .B(decoded_imm_j[3]), .Y(_04208_));
AND_g _25539_ (.A(_04207_), .B(_04208_), .Y(_04209_));
NAND_g _25540_ (.A(_04206_), .B(_04209_), .Y(_04210_));
NAND_g _25541_ (.A(_12314_), .B(_04210_), .Y(_04211_));
NAND_g _25542_ (.A(decoded_imm[3]), .B(_12315_), .Y(_04212_));
NAND_g _25543_ (.A(_04211_), .B(_04212_), .Y(_00908_));
NAND_g _25544_ (.A(mem_rdata_q[22]), .B(_12484_), .Y(_04213_));
NAND_g _25545_ (.A(instr_jal), .B(decoded_imm_j[2]), .Y(_04214_));
NAND_g _25546_ (.A(mem_rdata_q[9]), .B(_04082_), .Y(_04215_));
NOR_g _25547_ (.A(decoded_imm[2]), .B(_12314_), .Y(_04216_));
AND_g _25548_ (.A(_12314_), .B(_04214_), .Y(_04217_));
AND_g _25549_ (.A(_04213_), .B(_04217_), .Y(_04218_));
AND_g _25550_ (.A(_04215_), .B(_04218_), .Y(_04219_));
NOR_g _25551_ (.A(_04216_), .B(_04219_), .Y(_00909_));
NAND_g _25552_ (.A(mem_rdata_q[21]), .B(_12484_), .Y(_04220_));
NAND_g _25553_ (.A(mem_rdata_q[8]), .B(_04082_), .Y(_04221_));
NOR_g _25554_ (.A(_12315_), .B(_12727_), .Y(_04222_));
AND_g _25555_ (.A(_04221_), .B(_04222_), .Y(_04223_));
AND_g _25556_ (.A(_04220_), .B(_04223_), .Y(_04224_));
NOR_g _25557_ (.A(decoded_imm[1]), .B(_12314_), .Y(_04225_));
NOR_g _25558_ (.A(_04224_), .B(_04225_), .Y(_00910_));
AND_g _25559_ (.A(_11287_), .B(_11932_), .Y(_04226_));
NAND_g _25560_ (.A(_11287_), .B(_11932_), .Y(_04227_));
NAND_g _25561_ (.A(cpuregs_31[0]), .B(_04227_), .Y(_04228_));
NAND_g _25562_ (.A(_11301_), .B(_04226_), .Y(_04229_));
NAND_g _25563_ (.A(_04228_), .B(_04229_), .Y(_00911_));
NAND_g _25564_ (.A(cpuregs_31[1]), .B(_04227_), .Y(_04230_));
NAND_g _25565_ (.A(_11310_), .B(_04226_), .Y(_04231_));
NAND_g _25566_ (.A(_04230_), .B(_04231_), .Y(_00912_));
NAND_g _25567_ (.A(cpuregs_31[2]), .B(_04227_), .Y(_04232_));
NAND_g _25568_ (.A(_11319_), .B(_04226_), .Y(_04233_));
NAND_g _25569_ (.A(_04232_), .B(_04233_), .Y(_00913_));
NAND_g _25570_ (.A(cpuregs_31[3]), .B(_04227_), .Y(_04234_));
NAND_g _25571_ (.A(_11332_), .B(_04226_), .Y(_04235_));
NAND_g _25572_ (.A(_04234_), .B(_04235_), .Y(_00914_));
NAND_g _25573_ (.A(cpuregs_31[4]), .B(_04227_), .Y(_04236_));
NAND_g _25574_ (.A(_11345_), .B(_04226_), .Y(_04237_));
NAND_g _25575_ (.A(_04236_), .B(_04237_), .Y(_00915_));
NAND_g _25576_ (.A(cpuregs_31[5]), .B(_04227_), .Y(_04238_));
NAND_g _25577_ (.A(_11358_), .B(_04226_), .Y(_04239_));
NAND_g _25578_ (.A(_04238_), .B(_04239_), .Y(_00916_));
NAND_g _25579_ (.A(cpuregs_31[6]), .B(_04227_), .Y(_04240_));
NAND_g _25580_ (.A(_11371_), .B(_04226_), .Y(_04241_));
NAND_g _25581_ (.A(_04240_), .B(_04241_), .Y(_00917_));
NAND_g _25582_ (.A(cpuregs_31[7]), .B(_04227_), .Y(_04242_));
NAND_g _25583_ (.A(_11384_), .B(_04226_), .Y(_04243_));
NAND_g _25584_ (.A(_04242_), .B(_04243_), .Y(_00918_));
NAND_g _25585_ (.A(cpuregs_31[8]), .B(_04227_), .Y(_04244_));
NAND_g _25586_ (.A(_11397_), .B(_04226_), .Y(_04245_));
NAND_g _25587_ (.A(_04244_), .B(_04245_), .Y(_00919_));
NAND_g _25588_ (.A(cpuregs_31[9]), .B(_04227_), .Y(_04246_));
NAND_g _25589_ (.A(_11410_), .B(_04226_), .Y(_04247_));
NAND_g _25590_ (.A(_04246_), .B(_04247_), .Y(_00920_));
NAND_g _25591_ (.A(cpuregs_31[10]), .B(_04227_), .Y(_04248_));
NAND_g _25592_ (.A(_11423_), .B(_04226_), .Y(_04249_));
NAND_g _25593_ (.A(_04248_), .B(_04249_), .Y(_00921_));
NAND_g _25594_ (.A(cpuregs_31[11]), .B(_04227_), .Y(_04250_));
NAND_g _25595_ (.A(_11436_), .B(_04226_), .Y(_04251_));
NAND_g _25596_ (.A(_04250_), .B(_04251_), .Y(_00922_));
NAND_g _25597_ (.A(cpuregs_31[12]), .B(_04227_), .Y(_04252_));
NAND_g _25598_ (.A(_11449_), .B(_04226_), .Y(_04253_));
NAND_g _25599_ (.A(_04252_), .B(_04253_), .Y(_00923_));
NAND_g _25600_ (.A(cpuregs_31[13]), .B(_04227_), .Y(_04254_));
NAND_g _25601_ (.A(_11462_), .B(_04226_), .Y(_04255_));
NAND_g _25602_ (.A(_04254_), .B(_04255_), .Y(_00924_));
NAND_g _25603_ (.A(cpuregs_31[14]), .B(_04227_), .Y(_04256_));
NAND_g _25604_ (.A(_11475_), .B(_04226_), .Y(_04257_));
NAND_g _25605_ (.A(_04256_), .B(_04257_), .Y(_00925_));
NAND_g _25606_ (.A(cpuregs_31[15]), .B(_04227_), .Y(_04258_));
NAND_g _25607_ (.A(_11488_), .B(_04226_), .Y(_04259_));
NAND_g _25608_ (.A(_04258_), .B(_04259_), .Y(_00926_));
NAND_g _25609_ (.A(cpuregs_31[16]), .B(_04227_), .Y(_04260_));
NAND_g _25610_ (.A(_11501_), .B(_04226_), .Y(_04261_));
NAND_g _25611_ (.A(_04260_), .B(_04261_), .Y(_00927_));
NAND_g _25612_ (.A(_11514_), .B(_04226_), .Y(_04262_));
NAND_g _25613_ (.A(cpuregs_31[17]), .B(_04227_), .Y(_04263_));
NAND_g _25614_ (.A(_04262_), .B(_04263_), .Y(_00928_));
NAND_g _25615_ (.A(_11527_), .B(_04226_), .Y(_04264_));
NAND_g _25616_ (.A(cpuregs_31[18]), .B(_04227_), .Y(_04265_));
NAND_g _25617_ (.A(_04264_), .B(_04265_), .Y(_00929_));
NAND_g _25618_ (.A(_11540_), .B(_04226_), .Y(_04266_));
NAND_g _25619_ (.A(cpuregs_31[19]), .B(_04227_), .Y(_04267_));
NAND_g _25620_ (.A(_04266_), .B(_04267_), .Y(_00930_));
NAND_g _25621_ (.A(_11553_), .B(_04226_), .Y(_04268_));
NAND_g _25622_ (.A(cpuregs_31[20]), .B(_04227_), .Y(_04269_));
NAND_g _25623_ (.A(_04268_), .B(_04269_), .Y(_00931_));
NAND_g _25624_ (.A(_11566_), .B(_04226_), .Y(_04270_));
NAND_g _25625_ (.A(cpuregs_31[21]), .B(_04227_), .Y(_04271_));
NAND_g _25626_ (.A(_04270_), .B(_04271_), .Y(_00932_));
NAND_g _25627_ (.A(_11579_), .B(_04226_), .Y(_04272_));
NAND_g _25628_ (.A(cpuregs_31[22]), .B(_04227_), .Y(_04273_));
NAND_g _25629_ (.A(_04272_), .B(_04273_), .Y(_00933_));
NAND_g _25630_ (.A(_11592_), .B(_04226_), .Y(_04274_));
NAND_g _25631_ (.A(cpuregs_31[23]), .B(_04227_), .Y(_04275_));
NAND_g _25632_ (.A(_04274_), .B(_04275_), .Y(_00934_));
NAND_g _25633_ (.A(_11605_), .B(_04226_), .Y(_04276_));
NAND_g _25634_ (.A(cpuregs_31[24]), .B(_04227_), .Y(_04277_));
NAND_g _25635_ (.A(_04276_), .B(_04277_), .Y(_00935_));
NAND_g _25636_ (.A(_11618_), .B(_04226_), .Y(_04278_));
NAND_g _25637_ (.A(cpuregs_31[25]), .B(_04227_), .Y(_04279_));
NAND_g _25638_ (.A(_04278_), .B(_04279_), .Y(_00936_));
NAND_g _25639_ (.A(_11631_), .B(_04226_), .Y(_04280_));
NAND_g _25640_ (.A(cpuregs_31[26]), .B(_04227_), .Y(_04281_));
NAND_g _25641_ (.A(_04280_), .B(_04281_), .Y(_00937_));
NAND_g _25642_ (.A(_11644_), .B(_04226_), .Y(_04282_));
NAND_g _25643_ (.A(cpuregs_31[27]), .B(_04227_), .Y(_04283_));
NAND_g _25644_ (.A(_04282_), .B(_04283_), .Y(_00938_));
NAND_g _25645_ (.A(_11657_), .B(_04226_), .Y(_04284_));
NAND_g _25646_ (.A(cpuregs_31[28]), .B(_04227_), .Y(_04285_));
NAND_g _25647_ (.A(_04284_), .B(_04285_), .Y(_00939_));
NAND_g _25648_ (.A(_11670_), .B(_04226_), .Y(_04286_));
NAND_g _25649_ (.A(cpuregs_31[29]), .B(_04227_), .Y(_04287_));
NAND_g _25650_ (.A(_04286_), .B(_04287_), .Y(_00940_));
NAND_g _25651_ (.A(_11683_), .B(_04226_), .Y(_04288_));
NAND_g _25652_ (.A(cpuregs_31[30]), .B(_04227_), .Y(_04289_));
NAND_g _25653_ (.A(_04288_), .B(_04289_), .Y(_00941_));
NAND_g _25654_ (.A(_11695_), .B(_04226_), .Y(_04290_));
NAND_g _25655_ (.A(cpuregs_31[31]), .B(_04227_), .Y(_04291_));
NAND_g _25656_ (.A(_04290_), .B(_04291_), .Y(_00942_));
AND_g _25657_ (.A(_11285_), .B(_11767_), .Y(_04292_));
AND_g _25658_ (.A(_11932_), .B(_04292_), .Y(_04293_));
NAND_g _25659_ (.A(_11932_), .B(_04292_), .Y(_04294_));
NAND_g _25660_ (.A(cpuregs_3[0]), .B(_04294_), .Y(_04295_));
NAND_g _25661_ (.A(_11301_), .B(_04293_), .Y(_04296_));
NAND_g _25662_ (.A(_04295_), .B(_04296_), .Y(_00943_));
NAND_g _25663_ (.A(cpuregs_3[1]), .B(_04294_), .Y(_04297_));
NAND_g _25664_ (.A(_11310_), .B(_04293_), .Y(_04298_));
NAND_g _25665_ (.A(_04297_), .B(_04298_), .Y(_00944_));
NAND_g _25666_ (.A(cpuregs_3[2]), .B(_04294_), .Y(_04299_));
NAND_g _25667_ (.A(_11319_), .B(_04293_), .Y(_04300_));
NAND_g _25668_ (.A(_04299_), .B(_04300_), .Y(_00945_));
NAND_g _25669_ (.A(cpuregs_3[3]), .B(_04294_), .Y(_04301_));
NAND_g _25670_ (.A(_11332_), .B(_04293_), .Y(_04302_));
NAND_g _25671_ (.A(_04301_), .B(_04302_), .Y(_00946_));
NAND_g _25672_ (.A(cpuregs_3[4]), .B(_04294_), .Y(_04303_));
NAND_g _25673_ (.A(_11345_), .B(_04293_), .Y(_04304_));
NAND_g _25674_ (.A(_04303_), .B(_04304_), .Y(_00947_));
NAND_g _25675_ (.A(cpuregs_3[5]), .B(_04294_), .Y(_04305_));
NAND_g _25676_ (.A(_11358_), .B(_04293_), .Y(_04306_));
NAND_g _25677_ (.A(_04305_), .B(_04306_), .Y(_00948_));
NAND_g _25678_ (.A(cpuregs_3[6]), .B(_04294_), .Y(_04307_));
NAND_g _25679_ (.A(_11371_), .B(_04293_), .Y(_04308_));
NAND_g _25680_ (.A(_04307_), .B(_04308_), .Y(_00949_));
NAND_g _25681_ (.A(cpuregs_3[7]), .B(_04294_), .Y(_04309_));
NAND_g _25682_ (.A(_11384_), .B(_04293_), .Y(_04310_));
NAND_g _25683_ (.A(_04309_), .B(_04310_), .Y(_00950_));
NAND_g _25684_ (.A(cpuregs_3[8]), .B(_04294_), .Y(_04311_));
NAND_g _25685_ (.A(_11397_), .B(_04293_), .Y(_04312_));
NAND_g _25686_ (.A(_04311_), .B(_04312_), .Y(_00951_));
NAND_g _25687_ (.A(cpuregs_3[9]), .B(_04294_), .Y(_04313_));
NAND_g _25688_ (.A(_11410_), .B(_04293_), .Y(_04314_));
NAND_g _25689_ (.A(_04313_), .B(_04314_), .Y(_00952_));
NAND_g _25690_ (.A(cpuregs_3[10]), .B(_04294_), .Y(_04315_));
NAND_g _25691_ (.A(_11423_), .B(_04293_), .Y(_04316_));
NAND_g _25692_ (.A(_04315_), .B(_04316_), .Y(_00953_));
NAND_g _25693_ (.A(cpuregs_3[11]), .B(_04294_), .Y(_04317_));
NAND_g _25694_ (.A(_11436_), .B(_04293_), .Y(_04318_));
NAND_g _25695_ (.A(_04317_), .B(_04318_), .Y(_00954_));
NAND_g _25696_ (.A(cpuregs_3[12]), .B(_04294_), .Y(_04319_));
NAND_g _25697_ (.A(_11449_), .B(_04293_), .Y(_04320_));
NAND_g _25698_ (.A(_04319_), .B(_04320_), .Y(_00955_));
NAND_g _25699_ (.A(cpuregs_3[13]), .B(_04294_), .Y(_04321_));
NAND_g _25700_ (.A(_11462_), .B(_04293_), .Y(_04322_));
NAND_g _25701_ (.A(_04321_), .B(_04322_), .Y(_00956_));
NAND_g _25702_ (.A(cpuregs_3[14]), .B(_04294_), .Y(_04323_));
NAND_g _25703_ (.A(_11475_), .B(_04293_), .Y(_04324_));
NAND_g _25704_ (.A(_04323_), .B(_04324_), .Y(_00957_));
NAND_g _25705_ (.A(cpuregs_3[15]), .B(_04294_), .Y(_04325_));
NAND_g _25706_ (.A(_11488_), .B(_04293_), .Y(_04326_));
NAND_g _25707_ (.A(_04325_), .B(_04326_), .Y(_00958_));
NAND_g _25708_ (.A(cpuregs_3[16]), .B(_04294_), .Y(_04327_));
NAND_g _25709_ (.A(_11501_), .B(_04293_), .Y(_04328_));
NAND_g _25710_ (.A(_04327_), .B(_04328_), .Y(_00959_));
NOR_g _25711_ (.A(cpuregs_3[17]), .B(_04293_), .Y(_04329_));
NOR_g _25712_ (.A(_11514_), .B(_04294_), .Y(_04330_));
NOR_g _25713_ (.A(_04329_), .B(_04330_), .Y(_00960_));
NAND_g _25714_ (.A(_11527_), .B(_04293_), .Y(_04331_));
NAND_g _25715_ (.A(cpuregs_3[18]), .B(_04294_), .Y(_04332_));
NAND_g _25716_ (.A(_04331_), .B(_04332_), .Y(_00961_));
NAND_g _25717_ (.A(_11540_), .B(_04293_), .Y(_04333_));
NAND_g _25718_ (.A(cpuregs_3[19]), .B(_04294_), .Y(_04334_));
NAND_g _25719_ (.A(_04333_), .B(_04334_), .Y(_00962_));
NAND_g _25720_ (.A(_11553_), .B(_04293_), .Y(_04335_));
NAND_g _25721_ (.A(cpuregs_3[20]), .B(_04294_), .Y(_04336_));
NAND_g _25722_ (.A(_04335_), .B(_04336_), .Y(_00963_));
NAND_g _25723_ (.A(_11566_), .B(_04293_), .Y(_04337_));
NAND_g _25724_ (.A(cpuregs_3[21]), .B(_04294_), .Y(_04338_));
NAND_g _25725_ (.A(_04337_), .B(_04338_), .Y(_00964_));
NAND_g _25726_ (.A(_11579_), .B(_04293_), .Y(_04339_));
NAND_g _25727_ (.A(cpuregs_3[22]), .B(_04294_), .Y(_04340_));
NAND_g _25728_ (.A(_04339_), .B(_04340_), .Y(_00965_));
NAND_g _25729_ (.A(_11592_), .B(_04293_), .Y(_04341_));
NAND_g _25730_ (.A(cpuregs_3[23]), .B(_04294_), .Y(_04342_));
NAND_g _25731_ (.A(_04341_), .B(_04342_), .Y(_00966_));
NAND_g _25732_ (.A(_11605_), .B(_04293_), .Y(_04343_));
NAND_g _25733_ (.A(cpuregs_3[24]), .B(_04294_), .Y(_04344_));
NAND_g _25734_ (.A(_04343_), .B(_04344_), .Y(_00967_));
NAND_g _25735_ (.A(_11618_), .B(_04293_), .Y(_04345_));
NAND_g _25736_ (.A(cpuregs_3[25]), .B(_04294_), .Y(_04346_));
NAND_g _25737_ (.A(_04345_), .B(_04346_), .Y(_00968_));
NAND_g _25738_ (.A(_11631_), .B(_04293_), .Y(_04347_));
NAND_g _25739_ (.A(cpuregs_3[26]), .B(_04294_), .Y(_04348_));
NAND_g _25740_ (.A(_04347_), .B(_04348_), .Y(_00969_));
NAND_g _25741_ (.A(_11644_), .B(_04293_), .Y(_04349_));
NAND_g _25742_ (.A(cpuregs_3[27]), .B(_04294_), .Y(_04350_));
NAND_g _25743_ (.A(_04349_), .B(_04350_), .Y(_00970_));
NAND_g _25744_ (.A(_11657_), .B(_04293_), .Y(_04351_));
NAND_g _25745_ (.A(cpuregs_3[28]), .B(_04294_), .Y(_04352_));
NAND_g _25746_ (.A(_04351_), .B(_04352_), .Y(_00971_));
NAND_g _25747_ (.A(_11670_), .B(_04293_), .Y(_04353_));
NAND_g _25748_ (.A(cpuregs_3[29]), .B(_04294_), .Y(_04354_));
NAND_g _25749_ (.A(_04353_), .B(_04354_), .Y(_00972_));
NAND_g _25750_ (.A(_11683_), .B(_04293_), .Y(_04355_));
NAND_g _25751_ (.A(cpuregs_3[30]), .B(_04294_), .Y(_04356_));
NAND_g _25752_ (.A(_04355_), .B(_04356_), .Y(_00973_));
NAND_g _25753_ (.A(_11695_), .B(_04293_), .Y(_04357_));
NAND_g _25754_ (.A(cpuregs_3[31]), .B(_04294_), .Y(_04358_));
NAND_g _25755_ (.A(_04357_), .B(_04358_), .Y(_00974_));
NAND_g _25756_ (.A(_11279_), .B(_11282_), .Y(_04359_));
AND_g _25757_ (.A(_11287_), .B(_04359_), .Y(_04360_));
NAND_g _25758_ (.A(_11287_), .B(_04359_), .Y(_04361_));
NAND_g _25759_ (.A(cpuregs_28[0]), .B(_04361_), .Y(_04362_));
NAND_g _25760_ (.A(_11301_), .B(_04360_), .Y(_04363_));
NAND_g _25761_ (.A(_04362_), .B(_04363_), .Y(_00975_));
NAND_g _25762_ (.A(cpuregs_28[1]), .B(_04361_), .Y(_04364_));
NAND_g _25763_ (.A(_11310_), .B(_04360_), .Y(_04365_));
NAND_g _25764_ (.A(_04364_), .B(_04365_), .Y(_00976_));
NAND_g _25765_ (.A(cpuregs_28[2]), .B(_04361_), .Y(_04366_));
NAND_g _25766_ (.A(_11319_), .B(_04360_), .Y(_04367_));
NAND_g _25767_ (.A(_04366_), .B(_04367_), .Y(_00977_));
NAND_g _25768_ (.A(cpuregs_28[3]), .B(_04361_), .Y(_04368_));
NAND_g _25769_ (.A(_11332_), .B(_04360_), .Y(_04369_));
NAND_g _25770_ (.A(_04368_), .B(_04369_), .Y(_00978_));
NAND_g _25771_ (.A(cpuregs_28[4]), .B(_04361_), .Y(_04370_));
NAND_g _25772_ (.A(_11345_), .B(_04360_), .Y(_04371_));
NAND_g _25773_ (.A(_04370_), .B(_04371_), .Y(_00979_));
NAND_g _25774_ (.A(cpuregs_28[5]), .B(_04361_), .Y(_04372_));
NAND_g _25775_ (.A(_11358_), .B(_04360_), .Y(_04373_));
NAND_g _25776_ (.A(_04372_), .B(_04373_), .Y(_00980_));
NAND_g _25777_ (.A(cpuregs_28[6]), .B(_04361_), .Y(_04374_));
NAND_g _25778_ (.A(_11371_), .B(_04360_), .Y(_04375_));
NAND_g _25779_ (.A(_04374_), .B(_04375_), .Y(_00981_));
NAND_g _25780_ (.A(cpuregs_28[7]), .B(_04361_), .Y(_04376_));
NAND_g _25781_ (.A(_11384_), .B(_04360_), .Y(_04377_));
NAND_g _25782_ (.A(_04376_), .B(_04377_), .Y(_00982_));
NAND_g _25783_ (.A(cpuregs_28[8]), .B(_04361_), .Y(_04378_));
NAND_g _25784_ (.A(_11397_), .B(_04360_), .Y(_04379_));
NAND_g _25785_ (.A(_04378_), .B(_04379_), .Y(_00983_));
NAND_g _25786_ (.A(cpuregs_28[9]), .B(_04361_), .Y(_04380_));
NAND_g _25787_ (.A(_11410_), .B(_04360_), .Y(_04381_));
NAND_g _25788_ (.A(_04380_), .B(_04381_), .Y(_00984_));
NAND_g _25789_ (.A(cpuregs_28[10]), .B(_04361_), .Y(_04382_));
NAND_g _25790_ (.A(_11423_), .B(_04360_), .Y(_04383_));
NAND_g _25791_ (.A(_04382_), .B(_04383_), .Y(_00985_));
NAND_g _25792_ (.A(cpuregs_28[11]), .B(_04361_), .Y(_04384_));
NAND_g _25793_ (.A(_11436_), .B(_04360_), .Y(_04385_));
NAND_g _25794_ (.A(_04384_), .B(_04385_), .Y(_00986_));
NAND_g _25795_ (.A(cpuregs_28[12]), .B(_04361_), .Y(_04386_));
NAND_g _25796_ (.A(_11449_), .B(_04360_), .Y(_04387_));
NAND_g _25797_ (.A(_04386_), .B(_04387_), .Y(_00987_));
NAND_g _25798_ (.A(cpuregs_28[13]), .B(_04361_), .Y(_04388_));
NAND_g _25799_ (.A(_11462_), .B(_04360_), .Y(_04389_));
NAND_g _25800_ (.A(_04388_), .B(_04389_), .Y(_00988_));
NAND_g _25801_ (.A(cpuregs_28[14]), .B(_04361_), .Y(_04390_));
NAND_g _25802_ (.A(_11475_), .B(_04360_), .Y(_04391_));
NAND_g _25803_ (.A(_04390_), .B(_04391_), .Y(_00989_));
NAND_g _25804_ (.A(cpuregs_28[15]), .B(_04361_), .Y(_04392_));
NAND_g _25805_ (.A(_11488_), .B(_04360_), .Y(_04393_));
NAND_g _25806_ (.A(_04392_), .B(_04393_), .Y(_00990_));
NAND_g _25807_ (.A(cpuregs_28[16]), .B(_04361_), .Y(_04394_));
NAND_g _25808_ (.A(_11501_), .B(_04360_), .Y(_04395_));
NAND_g _25809_ (.A(_04394_), .B(_04395_), .Y(_00991_));
AND_g _25810_ (.A(_11098_), .B(_04361_), .Y(_04396_));
NOR_g _25811_ (.A(_11514_), .B(_04361_), .Y(_04397_));
NOR_g _25812_ (.A(_04396_), .B(_04397_), .Y(_00992_));
AND_g _25813_ (.A(_11099_), .B(_04361_), .Y(_04398_));
NOR_g _25814_ (.A(_11527_), .B(_04361_), .Y(_04399_));
NOR_g _25815_ (.A(_04398_), .B(_04399_), .Y(_00993_));
NOR_g _25816_ (.A(cpuregs_28[19]), .B(_04360_), .Y(_04400_));
NOR_g _25817_ (.A(_11540_), .B(_04361_), .Y(_04401_));
NOR_g _25818_ (.A(_04400_), .B(_04401_), .Y(_00994_));
AND_g _25819_ (.A(_11100_), .B(_04361_), .Y(_04402_));
NOR_g _25820_ (.A(_11553_), .B(_04361_), .Y(_04403_));
NOR_g _25821_ (.A(_04402_), .B(_04403_), .Y(_00995_));
NOR_g _25822_ (.A(cpuregs_28[21]), .B(_04360_), .Y(_04404_));
NOR_g _25823_ (.A(_11566_), .B(_04361_), .Y(_04405_));
NOR_g _25824_ (.A(_04404_), .B(_04405_), .Y(_00996_));
NOR_g _25825_ (.A(cpuregs_28[22]), .B(_04360_), .Y(_04406_));
NOR_g _25826_ (.A(_11579_), .B(_04361_), .Y(_04407_));
NOR_g _25827_ (.A(_04406_), .B(_04407_), .Y(_00997_));
NOR_g _25828_ (.A(cpuregs_28[23]), .B(_04360_), .Y(_04408_));
NOR_g _25829_ (.A(_11592_), .B(_04361_), .Y(_04409_));
NOR_g _25830_ (.A(_04408_), .B(_04409_), .Y(_00998_));
NOR_g _25831_ (.A(cpuregs_28[24]), .B(_04360_), .Y(_04410_));
NOR_g _25832_ (.A(_11605_), .B(_04361_), .Y(_04411_));
NOR_g _25833_ (.A(_04410_), .B(_04411_), .Y(_00999_));
NOR_g _25834_ (.A(cpuregs_28[25]), .B(_04360_), .Y(_04412_));
NOR_g _25835_ (.A(_11618_), .B(_04361_), .Y(_04413_));
NOR_g _25836_ (.A(_04412_), .B(_04413_), .Y(_01000_));
NOR_g _25837_ (.A(cpuregs_28[26]), .B(_04360_), .Y(_04414_));
NOR_g _25838_ (.A(_11631_), .B(_04361_), .Y(_04415_));
NOR_g _25839_ (.A(_04414_), .B(_04415_), .Y(_01001_));
NOR_g _25840_ (.A(cpuregs_28[27]), .B(_04360_), .Y(_04416_));
NOR_g _25841_ (.A(_11644_), .B(_04361_), .Y(_04417_));
NOR_g _25842_ (.A(_04416_), .B(_04417_), .Y(_01002_));
NOR_g _25843_ (.A(cpuregs_28[28]), .B(_04360_), .Y(_04418_));
NOR_g _25844_ (.A(_11657_), .B(_04361_), .Y(_04419_));
NOR_g _25845_ (.A(_04418_), .B(_04419_), .Y(_01003_));
AND_g _25846_ (.A(_11101_), .B(_04361_), .Y(_04420_));
NOR_g _25847_ (.A(_11670_), .B(_04361_), .Y(_04421_));
NOR_g _25848_ (.A(_04420_), .B(_04421_), .Y(_01004_));
NOR_g _25849_ (.A(cpuregs_28[30]), .B(_04360_), .Y(_04422_));
NOR_g _25850_ (.A(_11683_), .B(_04361_), .Y(_04423_));
NOR_g _25851_ (.A(_04422_), .B(_04423_), .Y(_01005_));
NOR_g _25852_ (.A(cpuregs_28[31]), .B(_04360_), .Y(_04424_));
NOR_g _25853_ (.A(_11695_), .B(_04361_), .Y(_04425_));
NOR_g _25854_ (.A(_04424_), .B(_04425_), .Y(_01006_));
AND_g _25855_ (.A(_11044_), .B(_11286_), .Y(_04426_));
AND_g _25856_ (.A(_11765_), .B(_04426_), .Y(_04427_));
NAND_g _25857_ (.A(_11765_), .B(_04426_), .Y(_04428_));
NAND_g _25858_ (.A(_11301_), .B(_04427_), .Y(_04429_));
NAND_g _25859_ (.A(cpuregs_14[0]), .B(_04428_), .Y(_04430_));
NAND_g _25860_ (.A(_04429_), .B(_04430_), .Y(_01007_));
NAND_g _25861_ (.A(_11310_), .B(_04427_), .Y(_04431_));
NAND_g _25862_ (.A(cpuregs_14[1]), .B(_04428_), .Y(_04432_));
NAND_g _25863_ (.A(_04431_), .B(_04432_), .Y(_01008_));
NAND_g _25864_ (.A(_11319_), .B(_04427_), .Y(_04433_));
NAND_g _25865_ (.A(cpuregs_14[2]), .B(_04428_), .Y(_04434_));
NAND_g _25866_ (.A(_04433_), .B(_04434_), .Y(_01009_));
NAND_g _25867_ (.A(_11332_), .B(_04427_), .Y(_04435_));
NAND_g _25868_ (.A(cpuregs_14[3]), .B(_04428_), .Y(_04436_));
NAND_g _25869_ (.A(_04435_), .B(_04436_), .Y(_01010_));
NAND_g _25870_ (.A(_11345_), .B(_04427_), .Y(_04437_));
NAND_g _25871_ (.A(cpuregs_14[4]), .B(_04428_), .Y(_04438_));
NAND_g _25872_ (.A(_04437_), .B(_04438_), .Y(_01011_));
NAND_g _25873_ (.A(_11358_), .B(_04427_), .Y(_04439_));
NAND_g _25874_ (.A(cpuregs_14[5]), .B(_04428_), .Y(_04440_));
NAND_g _25875_ (.A(_04439_), .B(_04440_), .Y(_01012_));
NAND_g _25876_ (.A(_11371_), .B(_04427_), .Y(_04441_));
NAND_g _25877_ (.A(cpuregs_14[6]), .B(_04428_), .Y(_04442_));
NAND_g _25878_ (.A(_04441_), .B(_04442_), .Y(_01013_));
NAND_g _25879_ (.A(_11384_), .B(_04427_), .Y(_04443_));
NAND_g _25880_ (.A(cpuregs_14[7]), .B(_04428_), .Y(_04444_));
NAND_g _25881_ (.A(_04443_), .B(_04444_), .Y(_01014_));
NAND_g _25882_ (.A(_11397_), .B(_04427_), .Y(_04445_));
NAND_g _25883_ (.A(cpuregs_14[8]), .B(_04428_), .Y(_04446_));
NAND_g _25884_ (.A(_04445_), .B(_04446_), .Y(_01015_));
NAND_g _25885_ (.A(_11410_), .B(_04427_), .Y(_04447_));
NAND_g _25886_ (.A(cpuregs_14[9]), .B(_04428_), .Y(_04448_));
NAND_g _25887_ (.A(_04447_), .B(_04448_), .Y(_01016_));
NAND_g _25888_ (.A(_11423_), .B(_04427_), .Y(_04449_));
NAND_g _25889_ (.A(cpuregs_14[10]), .B(_04428_), .Y(_04450_));
NAND_g _25890_ (.A(_04449_), .B(_04450_), .Y(_01017_));
NAND_g _25891_ (.A(_11436_), .B(_04427_), .Y(_04451_));
NAND_g _25892_ (.A(cpuregs_14[11]), .B(_04428_), .Y(_04452_));
NAND_g _25893_ (.A(_04451_), .B(_04452_), .Y(_01018_));
NAND_g _25894_ (.A(_11449_), .B(_04427_), .Y(_04453_));
NAND_g _25895_ (.A(cpuregs_14[12]), .B(_04428_), .Y(_04454_));
NAND_g _25896_ (.A(_04453_), .B(_04454_), .Y(_01019_));
NAND_g _25897_ (.A(_11462_), .B(_04427_), .Y(_04455_));
NAND_g _25898_ (.A(cpuregs_14[13]), .B(_04428_), .Y(_04456_));
NAND_g _25899_ (.A(_04455_), .B(_04456_), .Y(_01020_));
NAND_g _25900_ (.A(_11475_), .B(_04427_), .Y(_04457_));
NAND_g _25901_ (.A(cpuregs_14[14]), .B(_04428_), .Y(_04458_));
NAND_g _25902_ (.A(_04457_), .B(_04458_), .Y(_01021_));
NAND_g _25903_ (.A(_11488_), .B(_04427_), .Y(_04459_));
NAND_g _25904_ (.A(cpuregs_14[15]), .B(_04428_), .Y(_04460_));
NAND_g _25905_ (.A(_04459_), .B(_04460_), .Y(_01022_));
NAND_g _25906_ (.A(_11501_), .B(_04427_), .Y(_04461_));
NAND_g _25907_ (.A(cpuregs_14[16]), .B(_04428_), .Y(_04462_));
NAND_g _25908_ (.A(_04461_), .B(_04462_), .Y(_01023_));
NAND_g _25909_ (.A(_11514_), .B(_04427_), .Y(_04463_));
NAND_g _25910_ (.A(cpuregs_14[17]), .B(_04428_), .Y(_04464_));
NAND_g _25911_ (.A(_04463_), .B(_04464_), .Y(_01024_));
NAND_g _25912_ (.A(_11527_), .B(_04427_), .Y(_04465_));
NAND_g _25913_ (.A(cpuregs_14[18]), .B(_04428_), .Y(_04466_));
NAND_g _25914_ (.A(_04465_), .B(_04466_), .Y(_01025_));
NAND_g _25915_ (.A(_11540_), .B(_04427_), .Y(_04467_));
NAND_g _25916_ (.A(cpuregs_14[19]), .B(_04428_), .Y(_04468_));
NAND_g _25917_ (.A(_04467_), .B(_04468_), .Y(_01026_));
NAND_g _25918_ (.A(_11553_), .B(_04427_), .Y(_04469_));
NAND_g _25919_ (.A(cpuregs_14[20]), .B(_04428_), .Y(_04470_));
NAND_g _25920_ (.A(_04469_), .B(_04470_), .Y(_01027_));
NAND_g _25921_ (.A(_11566_), .B(_04427_), .Y(_04471_));
NAND_g _25922_ (.A(cpuregs_14[21]), .B(_04428_), .Y(_04472_));
NAND_g _25923_ (.A(_04471_), .B(_04472_), .Y(_01028_));
NAND_g _25924_ (.A(_11579_), .B(_04427_), .Y(_04473_));
NAND_g _25925_ (.A(cpuregs_14[22]), .B(_04428_), .Y(_04474_));
NAND_g _25926_ (.A(_04473_), .B(_04474_), .Y(_01029_));
NAND_g _25927_ (.A(_11592_), .B(_04427_), .Y(_04475_));
NAND_g _25928_ (.A(cpuregs_14[23]), .B(_04428_), .Y(_04476_));
NAND_g _25929_ (.A(_04475_), .B(_04476_), .Y(_01030_));
NAND_g _25930_ (.A(_11605_), .B(_04427_), .Y(_04477_));
NAND_g _25931_ (.A(cpuregs_14[24]), .B(_04428_), .Y(_04478_));
NAND_g _25932_ (.A(_04477_), .B(_04478_), .Y(_01031_));
NAND_g _25933_ (.A(_11618_), .B(_04427_), .Y(_04479_));
NAND_g _25934_ (.A(cpuregs_14[25]), .B(_04428_), .Y(_04480_));
NAND_g _25935_ (.A(_04479_), .B(_04480_), .Y(_01032_));
NAND_g _25936_ (.A(_11631_), .B(_04427_), .Y(_04481_));
NAND_g _25937_ (.A(cpuregs_14[26]), .B(_04428_), .Y(_04482_));
NAND_g _25938_ (.A(_04481_), .B(_04482_), .Y(_01033_));
NAND_g _25939_ (.A(_11644_), .B(_04427_), .Y(_04483_));
NAND_g _25940_ (.A(cpuregs_14[27]), .B(_04428_), .Y(_04484_));
NAND_g _25941_ (.A(_04483_), .B(_04484_), .Y(_01034_));
NAND_g _25942_ (.A(_11657_), .B(_04427_), .Y(_04485_));
NAND_g _25943_ (.A(cpuregs_14[28]), .B(_04428_), .Y(_04486_));
NAND_g _25944_ (.A(_04485_), .B(_04486_), .Y(_01035_));
NAND_g _25945_ (.A(_11670_), .B(_04427_), .Y(_04487_));
NAND_g _25946_ (.A(cpuregs_14[29]), .B(_04428_), .Y(_04488_));
NAND_g _25947_ (.A(_04487_), .B(_04488_), .Y(_01036_));
NAND_g _25948_ (.A(_11683_), .B(_04427_), .Y(_04489_));
NAND_g _25949_ (.A(cpuregs_14[30]), .B(_04428_), .Y(_04490_));
NAND_g _25950_ (.A(_04489_), .B(_04490_), .Y(_01037_));
NAND_g _25951_ (.A(_11695_), .B(_04427_), .Y(_04491_));
NAND_g _25952_ (.A(cpuregs_14[31]), .B(_04428_), .Y(_04492_));
NAND_g _25953_ (.A(_04491_), .B(_04492_), .Y(_01038_));
AND_g _25954_ (.A(_11765_), .B(_12000_), .Y(_04493_));
NAND_g _25955_ (.A(_11765_), .B(_12000_), .Y(_04494_));
NAND_g _25956_ (.A(cpuregs_26[0]), .B(_04494_), .Y(_04495_));
NAND_g _25957_ (.A(_11301_), .B(_04493_), .Y(_04496_));
NAND_g _25958_ (.A(_04495_), .B(_04496_), .Y(_01039_));
NAND_g _25959_ (.A(cpuregs_26[1]), .B(_04494_), .Y(_04497_));
NAND_g _25960_ (.A(_11310_), .B(_04493_), .Y(_04498_));
NAND_g _25961_ (.A(_04497_), .B(_04498_), .Y(_01040_));
NAND_g _25962_ (.A(cpuregs_26[2]), .B(_04494_), .Y(_04499_));
NAND_g _25963_ (.A(_11319_), .B(_04493_), .Y(_04500_));
NAND_g _25964_ (.A(_04499_), .B(_04500_), .Y(_01041_));
NAND_g _25965_ (.A(cpuregs_26[3]), .B(_04494_), .Y(_04501_));
NAND_g _25966_ (.A(_11332_), .B(_04493_), .Y(_04502_));
NAND_g _25967_ (.A(_04501_), .B(_04502_), .Y(_01042_));
NAND_g _25968_ (.A(cpuregs_26[4]), .B(_04494_), .Y(_04503_));
NAND_g _25969_ (.A(_11345_), .B(_04493_), .Y(_04504_));
NAND_g _25970_ (.A(_04503_), .B(_04504_), .Y(_01043_));
NAND_g _25971_ (.A(cpuregs_26[5]), .B(_04494_), .Y(_04505_));
NAND_g _25972_ (.A(_11358_), .B(_04493_), .Y(_04506_));
NAND_g _25973_ (.A(_04505_), .B(_04506_), .Y(_01044_));
NAND_g _25974_ (.A(cpuregs_26[6]), .B(_04494_), .Y(_04507_));
NAND_g _25975_ (.A(_11371_), .B(_04493_), .Y(_04508_));
NAND_g _25976_ (.A(_04507_), .B(_04508_), .Y(_01045_));
NAND_g _25977_ (.A(cpuregs_26[7]), .B(_04494_), .Y(_04509_));
NAND_g _25978_ (.A(_11384_), .B(_04493_), .Y(_04510_));
NAND_g _25979_ (.A(_04509_), .B(_04510_), .Y(_01046_));
NAND_g _25980_ (.A(cpuregs_26[8]), .B(_04494_), .Y(_04511_));
NAND_g _25981_ (.A(_11397_), .B(_04493_), .Y(_04512_));
NAND_g _25982_ (.A(_04511_), .B(_04512_), .Y(_01047_));
NAND_g _25983_ (.A(cpuregs_26[9]), .B(_04494_), .Y(_04513_));
NAND_g _25984_ (.A(_11410_), .B(_04493_), .Y(_04514_));
NAND_g _25985_ (.A(_04513_), .B(_04514_), .Y(_01048_));
NAND_g _25986_ (.A(cpuregs_26[10]), .B(_04494_), .Y(_04515_));
NAND_g _25987_ (.A(_11423_), .B(_04493_), .Y(_04516_));
NAND_g _25988_ (.A(_04515_), .B(_04516_), .Y(_01049_));
NAND_g _25989_ (.A(cpuregs_26[11]), .B(_04494_), .Y(_04517_));
NAND_g _25990_ (.A(_11436_), .B(_04493_), .Y(_04518_));
NAND_g _25991_ (.A(_04517_), .B(_04518_), .Y(_01050_));
NAND_g _25992_ (.A(cpuregs_26[12]), .B(_04494_), .Y(_04519_));
NAND_g _25993_ (.A(_11449_), .B(_04493_), .Y(_04520_));
NAND_g _25994_ (.A(_04519_), .B(_04520_), .Y(_01051_));
NAND_g _25995_ (.A(cpuregs_26[13]), .B(_04494_), .Y(_04521_));
NAND_g _25996_ (.A(_11462_), .B(_04493_), .Y(_04522_));
NAND_g _25997_ (.A(_04521_), .B(_04522_), .Y(_01052_));
NAND_g _25998_ (.A(cpuregs_26[14]), .B(_04494_), .Y(_04523_));
NAND_g _25999_ (.A(_11475_), .B(_04493_), .Y(_04524_));
NAND_g _26000_ (.A(_04523_), .B(_04524_), .Y(_01053_));
NAND_g _26001_ (.A(cpuregs_26[15]), .B(_04494_), .Y(_04525_));
NAND_g _26002_ (.A(_11488_), .B(_04493_), .Y(_04526_));
NAND_g _26003_ (.A(_04525_), .B(_04526_), .Y(_01054_));
NAND_g _26004_ (.A(cpuregs_26[16]), .B(_04494_), .Y(_04527_));
NAND_g _26005_ (.A(_11501_), .B(_04493_), .Y(_04528_));
NAND_g _26006_ (.A(_04527_), .B(_04528_), .Y(_01055_));
NAND_g _26007_ (.A(_11514_), .B(_04493_), .Y(_04529_));
NAND_g _26008_ (.A(cpuregs_26[17]), .B(_04494_), .Y(_04530_));
NAND_g _26009_ (.A(_04529_), .B(_04530_), .Y(_01056_));
NAND_g _26010_ (.A(_11527_), .B(_04493_), .Y(_04531_));
NAND_g _26011_ (.A(cpuregs_26[18]), .B(_04494_), .Y(_04532_));
NAND_g _26012_ (.A(_04531_), .B(_04532_), .Y(_01057_));
NAND_g _26013_ (.A(_11540_), .B(_04493_), .Y(_04533_));
NAND_g _26014_ (.A(cpuregs_26[19]), .B(_04494_), .Y(_04534_));
NAND_g _26015_ (.A(_04533_), .B(_04534_), .Y(_01058_));
NAND_g _26016_ (.A(_11553_), .B(_04493_), .Y(_04535_));
NAND_g _26017_ (.A(cpuregs_26[20]), .B(_04494_), .Y(_04536_));
NAND_g _26018_ (.A(_04535_), .B(_04536_), .Y(_01059_));
NAND_g _26019_ (.A(_11566_), .B(_04493_), .Y(_04537_));
NAND_g _26020_ (.A(cpuregs_26[21]), .B(_04494_), .Y(_04538_));
NAND_g _26021_ (.A(_04537_), .B(_04538_), .Y(_01060_));
NAND_g _26022_ (.A(_11579_), .B(_04493_), .Y(_04539_));
NAND_g _26023_ (.A(cpuregs_26[22]), .B(_04494_), .Y(_04540_));
NAND_g _26024_ (.A(_04539_), .B(_04540_), .Y(_01061_));
NAND_g _26025_ (.A(_11592_), .B(_04493_), .Y(_04541_));
NAND_g _26026_ (.A(cpuregs_26[23]), .B(_04494_), .Y(_04542_));
NAND_g _26027_ (.A(_04541_), .B(_04542_), .Y(_01062_));
NAND_g _26028_ (.A(_11605_), .B(_04493_), .Y(_04543_));
NAND_g _26029_ (.A(cpuregs_26[24]), .B(_04494_), .Y(_04544_));
NAND_g _26030_ (.A(_04543_), .B(_04544_), .Y(_01063_));
NAND_g _26031_ (.A(_11618_), .B(_04493_), .Y(_04545_));
NAND_g _26032_ (.A(cpuregs_26[25]), .B(_04494_), .Y(_04546_));
NAND_g _26033_ (.A(_04545_), .B(_04546_), .Y(_01064_));
NAND_g _26034_ (.A(_11631_), .B(_04493_), .Y(_04547_));
NAND_g _26035_ (.A(cpuregs_26[26]), .B(_04494_), .Y(_04548_));
NAND_g _26036_ (.A(_04547_), .B(_04548_), .Y(_01065_));
NAND_g _26037_ (.A(_11644_), .B(_04493_), .Y(_04549_));
NAND_g _26038_ (.A(cpuregs_26[27]), .B(_04494_), .Y(_04550_));
NAND_g _26039_ (.A(_04549_), .B(_04550_), .Y(_01066_));
NAND_g _26040_ (.A(_11657_), .B(_04493_), .Y(_04551_));
NAND_g _26041_ (.A(cpuregs_26[28]), .B(_04494_), .Y(_04552_));
NAND_g _26042_ (.A(_04551_), .B(_04552_), .Y(_01067_));
NAND_g _26043_ (.A(_11670_), .B(_04493_), .Y(_04553_));
NAND_g _26044_ (.A(cpuregs_26[29]), .B(_04494_), .Y(_04554_));
NAND_g _26045_ (.A(_04553_), .B(_04554_), .Y(_01068_));
NAND_g _26046_ (.A(_11683_), .B(_04493_), .Y(_04555_));
NAND_g _26047_ (.A(cpuregs_26[30]), .B(_04494_), .Y(_04556_));
NAND_g _26048_ (.A(_04555_), .B(_04556_), .Y(_01069_));
NAND_g _26049_ (.A(_11695_), .B(_04493_), .Y(_04557_));
NAND_g _26050_ (.A(cpuregs_26[31]), .B(_04494_), .Y(_04558_));
NAND_g _26051_ (.A(_04557_), .B(_04558_), .Y(_01070_));
AND_g _26052_ (.A(_11289_), .B(_11768_), .Y(_04559_));
NAND_g _26053_ (.A(_11289_), .B(_11768_), .Y(_04560_));
NAND_g _26054_ (.A(cpuregs_5[0]), .B(_04560_), .Y(_04561_));
NAND_g _26055_ (.A(_11301_), .B(_04559_), .Y(_04562_));
NAND_g _26056_ (.A(_04561_), .B(_04562_), .Y(_01071_));
NAND_g _26057_ (.A(cpuregs_5[1]), .B(_04560_), .Y(_04563_));
NAND_g _26058_ (.A(_11310_), .B(_04559_), .Y(_04564_));
NAND_g _26059_ (.A(_04563_), .B(_04564_), .Y(_01072_));
NAND_g _26060_ (.A(cpuregs_5[2]), .B(_04560_), .Y(_04565_));
NAND_g _26061_ (.A(_11319_), .B(_04559_), .Y(_04566_));
NAND_g _26062_ (.A(_04565_), .B(_04566_), .Y(_01073_));
NAND_g _26063_ (.A(cpuregs_5[3]), .B(_04560_), .Y(_04567_));
NAND_g _26064_ (.A(_11332_), .B(_04559_), .Y(_04568_));
NAND_g _26065_ (.A(_04567_), .B(_04568_), .Y(_01074_));
NAND_g _26066_ (.A(cpuregs_5[4]), .B(_04560_), .Y(_04569_));
NAND_g _26067_ (.A(_11345_), .B(_04559_), .Y(_04570_));
NAND_g _26068_ (.A(_04569_), .B(_04570_), .Y(_01075_));
NAND_g _26069_ (.A(cpuregs_5[5]), .B(_04560_), .Y(_04571_));
NAND_g _26070_ (.A(_11358_), .B(_04559_), .Y(_04572_));
NAND_g _26071_ (.A(_04571_), .B(_04572_), .Y(_01076_));
NAND_g _26072_ (.A(cpuregs_5[6]), .B(_04560_), .Y(_04573_));
NAND_g _26073_ (.A(_11371_), .B(_04559_), .Y(_04574_));
NAND_g _26074_ (.A(_04573_), .B(_04574_), .Y(_01077_));
NAND_g _26075_ (.A(cpuregs_5[7]), .B(_04560_), .Y(_04575_));
NAND_g _26076_ (.A(_11384_), .B(_04559_), .Y(_04576_));
NAND_g _26077_ (.A(_04575_), .B(_04576_), .Y(_01078_));
NAND_g _26078_ (.A(cpuregs_5[8]), .B(_04560_), .Y(_04577_));
NAND_g _26079_ (.A(_11397_), .B(_04559_), .Y(_04578_));
NAND_g _26080_ (.A(_04577_), .B(_04578_), .Y(_01079_));
NAND_g _26081_ (.A(cpuregs_5[9]), .B(_04560_), .Y(_04579_));
NAND_g _26082_ (.A(_11410_), .B(_04559_), .Y(_04580_));
NAND_g _26083_ (.A(_04579_), .B(_04580_), .Y(_01080_));
NAND_g _26084_ (.A(cpuregs_5[10]), .B(_04560_), .Y(_04581_));
NAND_g _26085_ (.A(_11423_), .B(_04559_), .Y(_04582_));
NAND_g _26086_ (.A(_04581_), .B(_04582_), .Y(_01081_));
NAND_g _26087_ (.A(cpuregs_5[11]), .B(_04560_), .Y(_04583_));
NAND_g _26088_ (.A(_11436_), .B(_04559_), .Y(_04584_));
NAND_g _26089_ (.A(_04583_), .B(_04584_), .Y(_01082_));
NAND_g _26090_ (.A(cpuregs_5[12]), .B(_04560_), .Y(_04585_));
NAND_g _26091_ (.A(_11449_), .B(_04559_), .Y(_04586_));
NAND_g _26092_ (.A(_04585_), .B(_04586_), .Y(_01083_));
NAND_g _26093_ (.A(cpuregs_5[13]), .B(_04560_), .Y(_04587_));
NAND_g _26094_ (.A(_11462_), .B(_04559_), .Y(_04588_));
NAND_g _26095_ (.A(_04587_), .B(_04588_), .Y(_01084_));
NAND_g _26096_ (.A(cpuregs_5[14]), .B(_04560_), .Y(_04589_));
NAND_g _26097_ (.A(_11475_), .B(_04559_), .Y(_04590_));
NAND_g _26098_ (.A(_04589_), .B(_04590_), .Y(_01085_));
NAND_g _26099_ (.A(cpuregs_5[15]), .B(_04560_), .Y(_04591_));
NAND_g _26100_ (.A(_11488_), .B(_04559_), .Y(_04592_));
NAND_g _26101_ (.A(_04591_), .B(_04592_), .Y(_01086_));
NAND_g _26102_ (.A(cpuregs_5[16]), .B(_04560_), .Y(_04593_));
NAND_g _26103_ (.A(_11501_), .B(_04559_), .Y(_04594_));
NAND_g _26104_ (.A(_04593_), .B(_04594_), .Y(_01087_));
NOR_g _26105_ (.A(cpuregs_5[17]), .B(_04559_), .Y(_04595_));
NOR_g _26106_ (.A(_11514_), .B(_04560_), .Y(_04596_));
NOR_g _26107_ (.A(_04595_), .B(_04596_), .Y(_01088_));
NAND_g _26108_ (.A(cpuregs_5[18]), .B(_04560_), .Y(_04597_));
NAND_g _26109_ (.A(_11527_), .B(_04559_), .Y(_04598_));
NAND_g _26110_ (.A(_04597_), .B(_04598_), .Y(_01089_));
NAND_g _26111_ (.A(cpuregs_5[19]), .B(_04560_), .Y(_04599_));
NAND_g _26112_ (.A(_11540_), .B(_04559_), .Y(_04600_));
NAND_g _26113_ (.A(_04599_), .B(_04600_), .Y(_01090_));
NAND_g _26114_ (.A(cpuregs_5[20]), .B(_04560_), .Y(_04601_));
NAND_g _26115_ (.A(_11553_), .B(_04559_), .Y(_04602_));
NAND_g _26116_ (.A(_04601_), .B(_04602_), .Y(_01091_));
NAND_g _26117_ (.A(cpuregs_5[21]), .B(_04560_), .Y(_04603_));
NAND_g _26118_ (.A(_11566_), .B(_04559_), .Y(_04604_));
NAND_g _26119_ (.A(_04603_), .B(_04604_), .Y(_01092_));
NAND_g _26120_ (.A(cpuregs_5[22]), .B(_04560_), .Y(_04605_));
NAND_g _26121_ (.A(_11579_), .B(_04559_), .Y(_04606_));
NAND_g _26122_ (.A(_04605_), .B(_04606_), .Y(_01093_));
NAND_g _26123_ (.A(cpuregs_5[23]), .B(_04560_), .Y(_04607_));
NAND_g _26124_ (.A(_11592_), .B(_04559_), .Y(_04608_));
NAND_g _26125_ (.A(_04607_), .B(_04608_), .Y(_01094_));
NAND_g _26126_ (.A(cpuregs_5[24]), .B(_04560_), .Y(_04609_));
NAND_g _26127_ (.A(_11605_), .B(_04559_), .Y(_04610_));
NAND_g _26128_ (.A(_04609_), .B(_04610_), .Y(_01095_));
NAND_g _26129_ (.A(cpuregs_5[25]), .B(_04560_), .Y(_04611_));
NAND_g _26130_ (.A(_11618_), .B(_04559_), .Y(_04612_));
NAND_g _26131_ (.A(_04611_), .B(_04612_), .Y(_01096_));
NAND_g _26132_ (.A(cpuregs_5[26]), .B(_04560_), .Y(_04613_));
NAND_g _26133_ (.A(_11631_), .B(_04559_), .Y(_04614_));
NAND_g _26134_ (.A(_04613_), .B(_04614_), .Y(_01097_));
NAND_g _26135_ (.A(cpuregs_5[27]), .B(_04560_), .Y(_04615_));
NAND_g _26136_ (.A(_11644_), .B(_04559_), .Y(_04616_));
NAND_g _26137_ (.A(_04615_), .B(_04616_), .Y(_01098_));
NAND_g _26138_ (.A(cpuregs_5[28]), .B(_04560_), .Y(_04617_));
NAND_g _26139_ (.A(_11657_), .B(_04559_), .Y(_04618_));
NAND_g _26140_ (.A(_04617_), .B(_04618_), .Y(_01099_));
NAND_g _26141_ (.A(cpuregs_5[29]), .B(_04560_), .Y(_04619_));
NAND_g _26142_ (.A(_11670_), .B(_04559_), .Y(_04620_));
NAND_g _26143_ (.A(_04619_), .B(_04620_), .Y(_01100_));
NAND_g _26144_ (.A(cpuregs_5[30]), .B(_04560_), .Y(_04621_));
NAND_g _26145_ (.A(_11683_), .B(_04559_), .Y(_04622_));
NAND_g _26146_ (.A(_04621_), .B(_04622_), .Y(_01101_));
NAND_g _26147_ (.A(cpuregs_5[31]), .B(_04560_), .Y(_04623_));
NAND_g _26148_ (.A(_11695_), .B(_04559_), .Y(_04624_));
NAND_g _26149_ (.A(_04623_), .B(_04624_), .Y(_01102_));
AND_g _26150_ (.A(_11278_), .B(_04426_), .Y(_04625_));
NAND_g _26151_ (.A(_11278_), .B(_04426_), .Y(_04626_));
NAND_g _26152_ (.A(_11301_), .B(_04625_), .Y(_04627_));
NAND_g _26153_ (.A(cpuregs_12[0]), .B(_04626_), .Y(_04628_));
NAND_g _26154_ (.A(_04627_), .B(_04628_), .Y(_01103_));
NAND_g _26155_ (.A(_11310_), .B(_04625_), .Y(_04629_));
NAND_g _26156_ (.A(cpuregs_12[1]), .B(_04626_), .Y(_04630_));
NAND_g _26157_ (.A(_04629_), .B(_04630_), .Y(_01104_));
NAND_g _26158_ (.A(_11319_), .B(_04625_), .Y(_04631_));
NAND_g _26159_ (.A(cpuregs_12[2]), .B(_04626_), .Y(_04632_));
NAND_g _26160_ (.A(_04631_), .B(_04632_), .Y(_01105_));
NAND_g _26161_ (.A(_11332_), .B(_04625_), .Y(_04633_));
NAND_g _26162_ (.A(cpuregs_12[3]), .B(_04626_), .Y(_04634_));
NAND_g _26163_ (.A(_04633_), .B(_04634_), .Y(_01106_));
NAND_g _26164_ (.A(_11345_), .B(_04625_), .Y(_04635_));
NAND_g _26165_ (.A(cpuregs_12[4]), .B(_04626_), .Y(_04636_));
NAND_g _26166_ (.A(_04635_), .B(_04636_), .Y(_01107_));
NAND_g _26167_ (.A(_11358_), .B(_04625_), .Y(_04637_));
NAND_g _26168_ (.A(cpuregs_12[5]), .B(_04626_), .Y(_04638_));
NAND_g _26169_ (.A(_04637_), .B(_04638_), .Y(_01108_));
NAND_g _26170_ (.A(_11371_), .B(_04625_), .Y(_04639_));
NAND_g _26171_ (.A(cpuregs_12[6]), .B(_04626_), .Y(_04640_));
NAND_g _26172_ (.A(_04639_), .B(_04640_), .Y(_01109_));
NAND_g _26173_ (.A(_11384_), .B(_04625_), .Y(_04641_));
NAND_g _26174_ (.A(cpuregs_12[7]), .B(_04626_), .Y(_04642_));
NAND_g _26175_ (.A(_04641_), .B(_04642_), .Y(_01110_));
NAND_g _26176_ (.A(_11397_), .B(_04625_), .Y(_04643_));
NAND_g _26177_ (.A(cpuregs_12[8]), .B(_04626_), .Y(_04644_));
NAND_g _26178_ (.A(_04643_), .B(_04644_), .Y(_01111_));
NAND_g _26179_ (.A(_11410_), .B(_04625_), .Y(_04645_));
NAND_g _26180_ (.A(cpuregs_12[9]), .B(_04626_), .Y(_04646_));
NAND_g _26181_ (.A(_04645_), .B(_04646_), .Y(_01112_));
NAND_g _26182_ (.A(_11423_), .B(_04625_), .Y(_04647_));
NAND_g _26183_ (.A(cpuregs_12[10]), .B(_04626_), .Y(_04648_));
NAND_g _26184_ (.A(_04647_), .B(_04648_), .Y(_01113_));
NAND_g _26185_ (.A(_11436_), .B(_04625_), .Y(_04649_));
NAND_g _26186_ (.A(cpuregs_12[11]), .B(_04626_), .Y(_04650_));
NAND_g _26187_ (.A(_04649_), .B(_04650_), .Y(_01114_));
NAND_g _26188_ (.A(_11449_), .B(_04625_), .Y(_04651_));
NAND_g _26189_ (.A(cpuregs_12[12]), .B(_04626_), .Y(_04652_));
NAND_g _26190_ (.A(_04651_), .B(_04652_), .Y(_01115_));
NAND_g _26191_ (.A(_11462_), .B(_04625_), .Y(_04653_));
NAND_g _26192_ (.A(cpuregs_12[13]), .B(_04626_), .Y(_04654_));
NAND_g _26193_ (.A(_04653_), .B(_04654_), .Y(_01116_));
NAND_g _26194_ (.A(_11475_), .B(_04625_), .Y(_04655_));
NAND_g _26195_ (.A(cpuregs_12[14]), .B(_04626_), .Y(_04656_));
NAND_g _26196_ (.A(_04655_), .B(_04656_), .Y(_01117_));
NAND_g _26197_ (.A(_11488_), .B(_04625_), .Y(_04657_));
NAND_g _26198_ (.A(cpuregs_12[15]), .B(_04626_), .Y(_04658_));
NAND_g _26199_ (.A(_04657_), .B(_04658_), .Y(_01118_));
NAND_g _26200_ (.A(_11501_), .B(_04625_), .Y(_04659_));
NAND_g _26201_ (.A(cpuregs_12[16]), .B(_04626_), .Y(_04660_));
NAND_g _26202_ (.A(_04659_), .B(_04660_), .Y(_01119_));
NAND_g _26203_ (.A(_11514_), .B(_04625_), .Y(_04661_));
NAND_g _26204_ (.A(cpuregs_12[17]), .B(_04626_), .Y(_04662_));
NAND_g _26205_ (.A(_04661_), .B(_04662_), .Y(_01120_));
NAND_g _26206_ (.A(_11527_), .B(_04625_), .Y(_04663_));
NAND_g _26207_ (.A(cpuregs_12[18]), .B(_04626_), .Y(_04664_));
NAND_g _26208_ (.A(_04663_), .B(_04664_), .Y(_01121_));
NAND_g _26209_ (.A(_11540_), .B(_04625_), .Y(_04665_));
NAND_g _26210_ (.A(cpuregs_12[19]), .B(_04626_), .Y(_04666_));
NAND_g _26211_ (.A(_04665_), .B(_04666_), .Y(_01122_));
NAND_g _26212_ (.A(_11553_), .B(_04625_), .Y(_04667_));
NAND_g _26213_ (.A(cpuregs_12[20]), .B(_04626_), .Y(_04668_));
NAND_g _26214_ (.A(_04667_), .B(_04668_), .Y(_01123_));
NAND_g _26215_ (.A(_11566_), .B(_04625_), .Y(_04669_));
NAND_g _26216_ (.A(cpuregs_12[21]), .B(_04626_), .Y(_04670_));
NAND_g _26217_ (.A(_04669_), .B(_04670_), .Y(_01124_));
NAND_g _26218_ (.A(_11579_), .B(_04625_), .Y(_04671_));
NAND_g _26219_ (.A(cpuregs_12[22]), .B(_04626_), .Y(_04672_));
NAND_g _26220_ (.A(_04671_), .B(_04672_), .Y(_01125_));
NAND_g _26221_ (.A(_11592_), .B(_04625_), .Y(_04673_));
NAND_g _26222_ (.A(cpuregs_12[23]), .B(_04626_), .Y(_04674_));
NAND_g _26223_ (.A(_04673_), .B(_04674_), .Y(_01126_));
NAND_g _26224_ (.A(_11605_), .B(_04625_), .Y(_04675_));
NAND_g _26225_ (.A(cpuregs_12[24]), .B(_04626_), .Y(_04676_));
NAND_g _26226_ (.A(_04675_), .B(_04676_), .Y(_01127_));
NAND_g _26227_ (.A(_11618_), .B(_04625_), .Y(_04677_));
NAND_g _26228_ (.A(cpuregs_12[25]), .B(_04626_), .Y(_04678_));
NAND_g _26229_ (.A(_04677_), .B(_04678_), .Y(_01128_));
NAND_g _26230_ (.A(_11631_), .B(_04625_), .Y(_04679_));
NAND_g _26231_ (.A(cpuregs_12[26]), .B(_04626_), .Y(_04680_));
NAND_g _26232_ (.A(_04679_), .B(_04680_), .Y(_01129_));
NAND_g _26233_ (.A(_11644_), .B(_04625_), .Y(_04681_));
NAND_g _26234_ (.A(cpuregs_12[27]), .B(_04626_), .Y(_04682_));
NAND_g _26235_ (.A(_04681_), .B(_04682_), .Y(_01130_));
NAND_g _26236_ (.A(_11657_), .B(_04625_), .Y(_04683_));
NAND_g _26237_ (.A(cpuregs_12[28]), .B(_04626_), .Y(_04684_));
NAND_g _26238_ (.A(_04683_), .B(_04684_), .Y(_01131_));
NAND_g _26239_ (.A(_11670_), .B(_04625_), .Y(_04685_));
NAND_g _26240_ (.A(cpuregs_12[29]), .B(_04626_), .Y(_04686_));
NAND_g _26241_ (.A(_04685_), .B(_04686_), .Y(_01132_));
NAND_g _26242_ (.A(_11683_), .B(_04625_), .Y(_04687_));
NAND_g _26243_ (.A(cpuregs_12[30]), .B(_04626_), .Y(_04688_));
NAND_g _26244_ (.A(_04687_), .B(_04688_), .Y(_01133_));
NAND_g _26245_ (.A(_11695_), .B(_04625_), .Y(_04689_));
NAND_g _26246_ (.A(cpuregs_12[31]), .B(_04626_), .Y(_04690_));
NAND_g _26247_ (.A(_04689_), .B(_04690_), .Y(_01134_));
AND_g _26248_ (.A(_11768_), .B(_11932_), .Y(_04691_));
NAND_g _26249_ (.A(_11768_), .B(_11932_), .Y(_04692_));
NAND_g _26250_ (.A(cpuregs_7[0]), .B(_04692_), .Y(_04693_));
NAND_g _26251_ (.A(_11301_), .B(_04691_), .Y(_04694_));
NAND_g _26252_ (.A(_04693_), .B(_04694_), .Y(_01135_));
NAND_g _26253_ (.A(cpuregs_7[1]), .B(_04692_), .Y(_04695_));
NAND_g _26254_ (.A(_11310_), .B(_04691_), .Y(_04696_));
NAND_g _26255_ (.A(_04695_), .B(_04696_), .Y(_01136_));
NAND_g _26256_ (.A(cpuregs_7[2]), .B(_04692_), .Y(_04697_));
NAND_g _26257_ (.A(_11319_), .B(_04691_), .Y(_04698_));
NAND_g _26258_ (.A(_04697_), .B(_04698_), .Y(_01137_));
NAND_g _26259_ (.A(cpuregs_7[3]), .B(_04692_), .Y(_04699_));
NAND_g _26260_ (.A(_11332_), .B(_04691_), .Y(_04700_));
NAND_g _26261_ (.A(_04699_), .B(_04700_), .Y(_01138_));
NAND_g _26262_ (.A(cpuregs_7[4]), .B(_04692_), .Y(_04701_));
NAND_g _26263_ (.A(_11345_), .B(_04691_), .Y(_04702_));
NAND_g _26264_ (.A(_04701_), .B(_04702_), .Y(_01139_));
NAND_g _26265_ (.A(cpuregs_7[5]), .B(_04692_), .Y(_04703_));
NAND_g _26266_ (.A(_11358_), .B(_04691_), .Y(_04704_));
NAND_g _26267_ (.A(_04703_), .B(_04704_), .Y(_01140_));
NAND_g _26268_ (.A(cpuregs_7[6]), .B(_04692_), .Y(_04705_));
NAND_g _26269_ (.A(_11371_), .B(_04691_), .Y(_04706_));
NAND_g _26270_ (.A(_04705_), .B(_04706_), .Y(_01141_));
NAND_g _26271_ (.A(cpuregs_7[7]), .B(_04692_), .Y(_04707_));
NAND_g _26272_ (.A(_11384_), .B(_04691_), .Y(_04708_));
NAND_g _26273_ (.A(_04707_), .B(_04708_), .Y(_01142_));
NAND_g _26274_ (.A(cpuregs_7[8]), .B(_04692_), .Y(_04709_));
NAND_g _26275_ (.A(_11397_), .B(_04691_), .Y(_04710_));
NAND_g _26276_ (.A(_04709_), .B(_04710_), .Y(_01143_));
NAND_g _26277_ (.A(cpuregs_7[9]), .B(_04692_), .Y(_04711_));
NAND_g _26278_ (.A(_11410_), .B(_04691_), .Y(_04712_));
NAND_g _26279_ (.A(_04711_), .B(_04712_), .Y(_01144_));
NAND_g _26280_ (.A(cpuregs_7[10]), .B(_04692_), .Y(_04713_));
NAND_g _26281_ (.A(_11423_), .B(_04691_), .Y(_04714_));
NAND_g _26282_ (.A(_04713_), .B(_04714_), .Y(_01145_));
NAND_g _26283_ (.A(cpuregs_7[11]), .B(_04692_), .Y(_04715_));
NAND_g _26284_ (.A(_11436_), .B(_04691_), .Y(_04716_));
NAND_g _26285_ (.A(_04715_), .B(_04716_), .Y(_01146_));
NAND_g _26286_ (.A(cpuregs_7[12]), .B(_04692_), .Y(_04717_));
NAND_g _26287_ (.A(_11449_), .B(_04691_), .Y(_04718_));
NAND_g _26288_ (.A(_04717_), .B(_04718_), .Y(_01147_));
NAND_g _26289_ (.A(cpuregs_7[13]), .B(_04692_), .Y(_04719_));
NAND_g _26290_ (.A(_11462_), .B(_04691_), .Y(_04720_));
NAND_g _26291_ (.A(_04719_), .B(_04720_), .Y(_01148_));
NAND_g _26292_ (.A(cpuregs_7[14]), .B(_04692_), .Y(_04721_));
NAND_g _26293_ (.A(_11475_), .B(_04691_), .Y(_04722_));
NAND_g _26294_ (.A(_04721_), .B(_04722_), .Y(_01149_));
NAND_g _26295_ (.A(cpuregs_7[15]), .B(_04692_), .Y(_04723_));
NAND_g _26296_ (.A(_11488_), .B(_04691_), .Y(_04724_));
NAND_g _26297_ (.A(_04723_), .B(_04724_), .Y(_01150_));
NAND_g _26298_ (.A(cpuregs_7[16]), .B(_04692_), .Y(_04725_));
NAND_g _26299_ (.A(_11501_), .B(_04691_), .Y(_04726_));
NAND_g _26300_ (.A(_04725_), .B(_04726_), .Y(_01151_));
NOR_g _26301_ (.A(cpuregs_7[17]), .B(_04691_), .Y(_04727_));
NOR_g _26302_ (.A(_11514_), .B(_04692_), .Y(_04728_));
NOR_g _26303_ (.A(_04727_), .B(_04728_), .Y(_01152_));
NAND_g _26304_ (.A(_11527_), .B(_04691_), .Y(_04729_));
NAND_g _26305_ (.A(cpuregs_7[18]), .B(_04692_), .Y(_04730_));
NAND_g _26306_ (.A(_04729_), .B(_04730_), .Y(_01153_));
NAND_g _26307_ (.A(_11540_), .B(_04691_), .Y(_04731_));
NAND_g _26308_ (.A(cpuregs_7[19]), .B(_04692_), .Y(_04732_));
NAND_g _26309_ (.A(_04731_), .B(_04732_), .Y(_01154_));
NAND_g _26310_ (.A(_11553_), .B(_04691_), .Y(_04733_));
NAND_g _26311_ (.A(cpuregs_7[20]), .B(_04692_), .Y(_04734_));
NAND_g _26312_ (.A(_04733_), .B(_04734_), .Y(_01155_));
NAND_g _26313_ (.A(_11566_), .B(_04691_), .Y(_04735_));
NAND_g _26314_ (.A(cpuregs_7[21]), .B(_04692_), .Y(_04736_));
NAND_g _26315_ (.A(_04735_), .B(_04736_), .Y(_01156_));
NAND_g _26316_ (.A(_11579_), .B(_04691_), .Y(_04737_));
NAND_g _26317_ (.A(cpuregs_7[22]), .B(_04692_), .Y(_04738_));
NAND_g _26318_ (.A(_04737_), .B(_04738_), .Y(_01157_));
NAND_g _26319_ (.A(_11592_), .B(_04691_), .Y(_04739_));
NAND_g _26320_ (.A(cpuregs_7[23]), .B(_04692_), .Y(_04740_));
NAND_g _26321_ (.A(_04739_), .B(_04740_), .Y(_01158_));
NAND_g _26322_ (.A(_11605_), .B(_04691_), .Y(_04741_));
NAND_g _26323_ (.A(cpuregs_7[24]), .B(_04692_), .Y(_04742_));
NAND_g _26324_ (.A(_04741_), .B(_04742_), .Y(_01159_));
NAND_g _26325_ (.A(_11618_), .B(_04691_), .Y(_04743_));
NAND_g _26326_ (.A(cpuregs_7[25]), .B(_04692_), .Y(_04744_));
NAND_g _26327_ (.A(_04743_), .B(_04744_), .Y(_01160_));
NAND_g _26328_ (.A(_11631_), .B(_04691_), .Y(_04745_));
NAND_g _26329_ (.A(cpuregs_7[26]), .B(_04692_), .Y(_04746_));
NAND_g _26330_ (.A(_04745_), .B(_04746_), .Y(_01161_));
NAND_g _26331_ (.A(_11644_), .B(_04691_), .Y(_04747_));
NAND_g _26332_ (.A(cpuregs_7[27]), .B(_04692_), .Y(_04748_));
NAND_g _26333_ (.A(_04747_), .B(_04748_), .Y(_01162_));
NAND_g _26334_ (.A(_11657_), .B(_04691_), .Y(_04749_));
NAND_g _26335_ (.A(cpuregs_7[28]), .B(_04692_), .Y(_04750_));
NAND_g _26336_ (.A(_04749_), .B(_04750_), .Y(_01163_));
NAND_g _26337_ (.A(_11670_), .B(_04691_), .Y(_04751_));
NAND_g _26338_ (.A(cpuregs_7[29]), .B(_04692_), .Y(_04752_));
NAND_g _26339_ (.A(_04751_), .B(_04752_), .Y(_01164_));
NAND_g _26340_ (.A(_11683_), .B(_04691_), .Y(_04753_));
NAND_g _26341_ (.A(cpuregs_7[30]), .B(_04692_), .Y(_04754_));
NAND_g _26342_ (.A(_04753_), .B(_04754_), .Y(_01165_));
NAND_g _26343_ (.A(_11695_), .B(_04691_), .Y(_04755_));
NAND_g _26344_ (.A(cpuregs_7[31]), .B(_04692_), .Y(_04756_));
NAND_g _26345_ (.A(_04755_), .B(_04756_), .Y(_01166_));
NAND_g _26346_ (.A(_13409_), .B(_02239_), .Y(_04757_));
AND_g _26347_ (.A(_13726_), .B(_02618_), .Y(_04758_));
NOT_g _26348_ (.A(_04758_), .Y(dbg_ascii_state[24]));
NAND_g _26349_ (.A(_13412_), .B(_04758_), .Y(_04759_));
NOR_g _26350_ (.A(_13413_), .B(_02225_), .Y(_04760_));
NOT_g _26351_ (.A(_04760_), .Y(_04761_));
NAND_g _26352_ (.A(_04759_), .B(_04761_), .Y(_04762_));
NAND_g _26353_ (.A(cpu_state[0]), .B(_04762_), .Y(_04763_));
NAND_g _26354_ (.A(_04757_), .B(_04763_), .Y(_04764_));
NOR_g _26355_ (.A(reg_next_pc[0]), .B(reg_pc[1]), .Y(_04765_));
NOR_g _26356_ (.A(_11905_), .B(_04765_), .Y(_04766_));
NAND_g _26357_ (.A(_11135_), .B(_04049_), .Y(_04767_));
NAND_g _26358_ (.A(resetn), .B(_11013_), .Y(_04768_));
NOR_g _26359_ (.A(_11907_), .B(_04768_), .Y(_04769_));
AND_g _26360_ (.A(_04767_), .B(_04769_), .Y(_04770_));
NOR_g _26361_ (.A(_04766_), .B(_04770_), .Y(_04771_));
AND_g _26362_ (.A(resetn), .B(_04771_), .Y(_04772_));
AND_g _26363_ (.A(_04764_), .B(_04772_), .Y(_01167_));
NAND_g _26364_ (.A(cpu_state[1]), .B(_04762_), .Y(_04773_));
NAND_g _26365_ (.A(is_sb_sh_sw), .B(_14358_), .Y(_04774_));
NAND_g _26366_ (.A(_04773_), .B(_04774_), .Y(_04775_));
AND_g _26367_ (.A(_04772_), .B(_04775_), .Y(_01168_));
NAND_g _26368_ (.A(is_sll_srl_sra), .B(_14358_), .Y(_04776_));
AND_g _26369_ (.A(is_slli_srli_srai), .B(_13409_), .Y(_04777_));
NAND_g _26370_ (.A(_13390_), .B(_04759_), .Y(_04778_));
AND_g _26371_ (.A(cpu_state[2]), .B(_04778_), .Y(_04779_));
NOR_g _26372_ (.A(_04777_), .B(_04779_), .Y(_04780_));
NAND_g _26373_ (.A(_04776_), .B(_04780_), .Y(_04781_));
AND_g _26374_ (.A(_04772_), .B(_04781_), .Y(_01169_));
NOR_g _26375_ (.A(is_sll_srl_sra), .B(is_sb_sh_sw), .Y(_04782_));
NAND_g _26376_ (.A(_13832_), .B(_04782_), .Y(_04783_));
NAND_g _26377_ (.A(_13829_), .B(_04783_), .Y(_04784_));
NAND_g _26378_ (.A(_13409_), .B(_04784_), .Y(_04785_));
NAND_g _26379_ (.A(is_beq_bne_blt_bge_bltu_bgeu), .B(_11916_), .Y(_04786_));
NAND_g _26380_ (.A(_04759_), .B(_04786_), .Y(_04787_));
NAND_g _26381_ (.A(cpu_state[3]), .B(_04787_), .Y(_04788_));
NAND_g _26382_ (.A(_13724_), .B(_04782_), .Y(_04789_));
AND_g _26383_ (.A(_04788_), .B(_04789_), .Y(_04790_));
NAND_g _26384_ (.A(_04785_), .B(_04790_), .Y(_04791_));
AND_g _26385_ (.A(_04772_), .B(_04791_), .Y(_01170_));
NAND_g _26386_ (.A(cpu_state[4]), .B(_04772_), .Y(_04792_));
NOR_g _26387_ (.A(_04759_), .B(_04792_), .Y(_01171_));
AND_g _26388_ (.A(_11263_), .B(_04759_), .Y(_04793_));
NOR_g _26389_ (.A(cpu_state[5]), .B(_12537_), .Y(_04794_));
NOR_g _26390_ (.A(_04793_), .B(_04794_), .Y(_04795_));
AND_g _26391_ (.A(_04772_), .B(_04795_), .Y(_01172_));
NOR_g _26392_ (.A(dbg_ascii_state[27]), .B(dbg_ascii_state[18]), .Y(_04796_));
NOT_g _26393_ (.A(_04796_), .Y(dbg_ascii_state[38]));
NAND_g _26394_ (.A(cpu_state[6]), .B(_04796_), .Y(_04797_));
NAND_g _26395_ (.A(_11271_), .B(_04786_), .Y(_04798_));
NAND_g _26396_ (.A(resetn), .B(_02620_), .Y(_04799_));
NOR_g _26397_ (.A(_13416_), .B(_04799_), .Y(_04800_));
AND_g _26398_ (.A(_02244_), .B(_04800_), .Y(_04801_));
AND_g _26399_ (.A(_04798_), .B(_04801_), .Y(_04802_));
AND_g _26400_ (.A(_04797_), .B(_04802_), .Y(_04803_));
NAND_g _26401_ (.A(_02226_), .B(_04803_), .Y(_04804_));
AND_g _26402_ (.A(_04771_), .B(_04804_), .Y(_01173_));
AND_g _26403_ (.A(resetn), .B(_13409_), .Y(_04805_));
NAND_g _26404_ (.A(resetn), .B(_13409_), .Y(_04806_));
NAND_g _26405_ (.A(_13609_), .B(_04805_), .Y(_04807_));
NAND_g _26406_ (.A(resetn), .B(cpu_state[7]), .Y(_04808_));
AND_g _26407_ (.A(_04771_), .B(_04808_), .Y(_04809_));
NAND_g _26408_ (.A(_04807_), .B(_04809_), .Y(_01174_));
AND_g _26409_ (.A(_11278_), .B(_11697_), .Y(_04810_));
NAND_g _26410_ (.A(_11278_), .B(_11697_), .Y(_04811_));
NAND_g _26411_ (.A(cpuregs_8[0]), .B(_04811_), .Y(_04812_));
NAND_g _26412_ (.A(_11300_), .B(_04810_), .Y(_04813_));
NAND_g _26413_ (.A(_04812_), .B(_04813_), .Y(_01175_));
NAND_g _26414_ (.A(cpuregs_8[1]), .B(_04811_), .Y(_04814_));
NAND_g _26415_ (.A(_11309_), .B(_04810_), .Y(_04815_));
NAND_g _26416_ (.A(_04814_), .B(_04815_), .Y(_01176_));
NAND_g _26417_ (.A(cpuregs_8[2]), .B(_04811_), .Y(_04816_));
NAND_g _26418_ (.A(_11318_), .B(_04810_), .Y(_04817_));
NAND_g _26419_ (.A(_04816_), .B(_04817_), .Y(_01177_));
NAND_g _26420_ (.A(cpuregs_8[3]), .B(_04811_), .Y(_04818_));
NAND_g _26421_ (.A(_11331_), .B(_04810_), .Y(_04819_));
NAND_g _26422_ (.A(_04818_), .B(_04819_), .Y(_01178_));
NAND_g _26423_ (.A(cpuregs_8[4]), .B(_04811_), .Y(_04820_));
NAND_g _26424_ (.A(_11344_), .B(_04810_), .Y(_04821_));
NAND_g _26425_ (.A(_04820_), .B(_04821_), .Y(_01179_));
NAND_g _26426_ (.A(cpuregs_8[5]), .B(_04811_), .Y(_04822_));
NAND_g _26427_ (.A(_11357_), .B(_04810_), .Y(_04823_));
NAND_g _26428_ (.A(_04822_), .B(_04823_), .Y(_01180_));
NAND_g _26429_ (.A(cpuregs_8[6]), .B(_04811_), .Y(_04824_));
NAND_g _26430_ (.A(_11370_), .B(_04810_), .Y(_04825_));
NAND_g _26431_ (.A(_04824_), .B(_04825_), .Y(_01181_));
NAND_g _26432_ (.A(cpuregs_8[7]), .B(_04811_), .Y(_04826_));
NAND_g _26433_ (.A(_11383_), .B(_04810_), .Y(_04827_));
NAND_g _26434_ (.A(_04826_), .B(_04827_), .Y(_01182_));
NAND_g _26435_ (.A(cpuregs_8[8]), .B(_04811_), .Y(_04828_));
NAND_g _26436_ (.A(_11396_), .B(_04810_), .Y(_04829_));
NAND_g _26437_ (.A(_04828_), .B(_04829_), .Y(_01183_));
NAND_g _26438_ (.A(cpuregs_8[9]), .B(_04811_), .Y(_04830_));
NAND_g _26439_ (.A(_11409_), .B(_04810_), .Y(_04831_));
NAND_g _26440_ (.A(_04830_), .B(_04831_), .Y(_01184_));
NAND_g _26441_ (.A(cpuregs_8[10]), .B(_04811_), .Y(_04832_));
NAND_g _26442_ (.A(_11422_), .B(_04810_), .Y(_04833_));
NAND_g _26443_ (.A(_04832_), .B(_04833_), .Y(_01185_));
NAND_g _26444_ (.A(cpuregs_8[11]), .B(_04811_), .Y(_04834_));
NAND_g _26445_ (.A(_11435_), .B(_04810_), .Y(_04835_));
NAND_g _26446_ (.A(_04834_), .B(_04835_), .Y(_01186_));
NAND_g _26447_ (.A(cpuregs_8[12]), .B(_04811_), .Y(_04836_));
NAND_g _26448_ (.A(_11448_), .B(_04810_), .Y(_04837_));
NAND_g _26449_ (.A(_04836_), .B(_04837_), .Y(_01187_));
NAND_g _26450_ (.A(cpuregs_8[13]), .B(_04811_), .Y(_04838_));
NAND_g _26451_ (.A(_11461_), .B(_04810_), .Y(_04839_));
NAND_g _26452_ (.A(_04838_), .B(_04839_), .Y(_01188_));
NAND_g _26453_ (.A(cpuregs_8[14]), .B(_04811_), .Y(_04840_));
NAND_g _26454_ (.A(_11474_), .B(_04810_), .Y(_04841_));
NAND_g _26455_ (.A(_04840_), .B(_04841_), .Y(_01189_));
NAND_g _26456_ (.A(cpuregs_8[15]), .B(_04811_), .Y(_04842_));
NAND_g _26457_ (.A(_11487_), .B(_04810_), .Y(_04843_));
NAND_g _26458_ (.A(_04842_), .B(_04843_), .Y(_01190_));
NOR_g _26459_ (.A(_11500_), .B(_04811_), .Y(_04844_));
NOR_g _26460_ (.A(cpuregs_8[16]), .B(_04810_), .Y(_04845_));
NOR_g _26461_ (.A(_04844_), .B(_04845_), .Y(_01191_));
NAND_g _26462_ (.A(cpuregs_8[17]), .B(_04811_), .Y(_04846_));
NAND_g _26463_ (.A(_11513_), .B(_04810_), .Y(_04847_));
NAND_g _26464_ (.A(_04846_), .B(_04847_), .Y(_01192_));
NAND_g _26465_ (.A(cpuregs_8[18]), .B(_04811_), .Y(_04848_));
NAND_g _26466_ (.A(_11526_), .B(_04810_), .Y(_04849_));
NAND_g _26467_ (.A(_04848_), .B(_04849_), .Y(_01193_));
NAND_g _26468_ (.A(cpuregs_8[19]), .B(_04811_), .Y(_04850_));
NAND_g _26469_ (.A(_11539_), .B(_04810_), .Y(_04851_));
NAND_g _26470_ (.A(_04850_), .B(_04851_), .Y(_01194_));
NAND_g _26471_ (.A(cpuregs_8[20]), .B(_04811_), .Y(_04852_));
NAND_g _26472_ (.A(_11552_), .B(_04810_), .Y(_04853_));
NAND_g _26473_ (.A(_04852_), .B(_04853_), .Y(_01195_));
NAND_g _26474_ (.A(cpuregs_8[21]), .B(_04811_), .Y(_04854_));
NAND_g _26475_ (.A(_11565_), .B(_04810_), .Y(_04855_));
NAND_g _26476_ (.A(_04854_), .B(_04855_), .Y(_01196_));
NAND_g _26477_ (.A(cpuregs_8[22]), .B(_04811_), .Y(_04856_));
NAND_g _26478_ (.A(_11578_), .B(_04810_), .Y(_04857_));
NAND_g _26479_ (.A(_04856_), .B(_04857_), .Y(_01197_));
NAND_g _26480_ (.A(cpuregs_8[23]), .B(_04811_), .Y(_04858_));
NAND_g _26481_ (.A(_11591_), .B(_04810_), .Y(_04859_));
NAND_g _26482_ (.A(_04858_), .B(_04859_), .Y(_01198_));
NAND_g _26483_ (.A(cpuregs_8[24]), .B(_04811_), .Y(_04860_));
NAND_g _26484_ (.A(_11604_), .B(_04810_), .Y(_04861_));
NAND_g _26485_ (.A(_04860_), .B(_04861_), .Y(_01199_));
NAND_g _26486_ (.A(cpuregs_8[25]), .B(_04811_), .Y(_04862_));
NAND_g _26487_ (.A(_11617_), .B(_04810_), .Y(_04863_));
NAND_g _26488_ (.A(_04862_), .B(_04863_), .Y(_01200_));
NAND_g _26489_ (.A(cpuregs_8[26]), .B(_04811_), .Y(_04864_));
NAND_g _26490_ (.A(_11630_), .B(_04810_), .Y(_04865_));
NAND_g _26491_ (.A(_04864_), .B(_04865_), .Y(_01201_));
NAND_g _26492_ (.A(cpuregs_8[27]), .B(_04811_), .Y(_04866_));
NAND_g _26493_ (.A(_11643_), .B(_04810_), .Y(_04867_));
NAND_g _26494_ (.A(_04866_), .B(_04867_), .Y(_01202_));
NAND_g _26495_ (.A(cpuregs_8[28]), .B(_04811_), .Y(_04868_));
NAND_g _26496_ (.A(_11656_), .B(_04810_), .Y(_04869_));
NAND_g _26497_ (.A(_04868_), .B(_04869_), .Y(_01203_));
NAND_g _26498_ (.A(cpuregs_8[29]), .B(_04811_), .Y(_04870_));
NAND_g _26499_ (.A(_11669_), .B(_04810_), .Y(_04871_));
NAND_g _26500_ (.A(_04870_), .B(_04871_), .Y(_01204_));
NAND_g _26501_ (.A(cpuregs_8[30]), .B(_04811_), .Y(_04872_));
NAND_g _26502_ (.A(_11682_), .B(_04810_), .Y(_04873_));
NAND_g _26503_ (.A(_04872_), .B(_04873_), .Y(_01205_));
NAND_g _26504_ (.A(cpuregs_8[31]), .B(_04811_), .Y(_04874_));
NAND_g _26505_ (.A(_11694_), .B(_04810_), .Y(_04875_));
NAND_g _26506_ (.A(_04874_), .B(_04875_), .Y(_01206_));
NOR_g _26507_ (.A(pcpi_rs1[0]), .B(_13425_), .Y(_04876_));
NAND_g _26508_ (.A(cpuregs_7[0]), .B(_00012_[2]), .Y(_04877_));
NAND_g _26509_ (.A(cpuregs_3[0]), .B(_11214_), .Y(_04878_));
NAND_g _26510_ (.A(_04877_), .B(_04878_), .Y(_04879_));
AND_g _26511_ (.A(_00012_[0]), .B(_04879_), .Y(_04880_));
NAND_g _26512_ (.A(cpuregs_6[0]), .B(_00012_[2]), .Y(_04881_));
NAND_g _26513_ (.A(cpuregs_2[0]), .B(_11214_), .Y(_04882_));
AND_g _26514_ (.A(_04881_), .B(_04882_), .Y(_04883_));
NOR_g _26515_ (.A(_00012_[0]), .B(_04883_), .Y(_04884_));
NOR_g _26516_ (.A(_04880_), .B(_04884_), .Y(_04885_));
NAND_g _26517_ (.A(cpuregs_5[0]), .B(_00012_[2]), .Y(_04886_));
NAND_g _26518_ (.A(cpuregs_1[0]), .B(_11214_), .Y(_04887_));
NAND_g _26519_ (.A(_04886_), .B(_04887_), .Y(_04888_));
NAND_g _26520_ (.A(_00012_[0]), .B(_04888_), .Y(_04889_));
NAND_g _26521_ (.A(cpuregs_4[0]), .B(_00012_[2]), .Y(_04890_));
NAND_g _26522_ (.A(cpuregs_0[0]), .B(_11214_), .Y(_04891_));
AND_g _26523_ (.A(_04890_), .B(_04891_), .Y(_04892_));
NOR_g _26524_ (.A(_00012_[0]), .B(_04892_), .Y(_04893_));
NAND_g _26525_ (.A(_00012_[1]), .B(_04885_), .Y(_04894_));
NOR_g _26526_ (.A(_00012_[1]), .B(_04893_), .Y(_04895_));
NAND_g _26527_ (.A(_04889_), .B(_04895_), .Y(_04896_));
AND_g _26528_ (.A(_04894_), .B(_04896_), .Y(_04897_));
NAND_g _26529_ (.A(_11215_), .B(_04897_), .Y(_04898_));
NAND_g _26530_ (.A(cpuregs_13[0]), .B(_00012_[0]), .Y(_04899_));
NAND_g _26531_ (.A(cpuregs_12[0]), .B(_11212_), .Y(_04900_));
AND_g _26532_ (.A(_00012_[2]), .B(_04900_), .Y(_04901_));
NAND_g _26533_ (.A(_04899_), .B(_04901_), .Y(_04902_));
NAND_g _26534_ (.A(cpuregs_9[0]), .B(_00012_[0]), .Y(_04903_));
NAND_g _26535_ (.A(cpuregs_8[0]), .B(_11212_), .Y(_04904_));
AND_g _26536_ (.A(_11214_), .B(_04904_), .Y(_04905_));
NAND_g _26537_ (.A(_04903_), .B(_04905_), .Y(_04906_));
AND_g _26538_ (.A(_11213_), .B(_04906_), .Y(_04907_));
NAND_g _26539_ (.A(_04902_), .B(_04907_), .Y(_04908_));
NAND_g _26540_ (.A(cpuregs_15[0]), .B(_00012_[0]), .Y(_04909_));
NAND_g _26541_ (.A(cpuregs_14[0]), .B(_11212_), .Y(_04910_));
AND_g _26542_ (.A(_00012_[2]), .B(_04910_), .Y(_04911_));
NAND_g _26543_ (.A(_04909_), .B(_04911_), .Y(_04912_));
NAND_g _26544_ (.A(cpuregs_11[0]), .B(_00012_[0]), .Y(_04913_));
NAND_g _26545_ (.A(cpuregs_10[0]), .B(_11212_), .Y(_04914_));
AND_g _26546_ (.A(_11214_), .B(_04914_), .Y(_04915_));
NAND_g _26547_ (.A(_04913_), .B(_04915_), .Y(_04916_));
AND_g _26548_ (.A(_00012_[1]), .B(_04916_), .Y(_04917_));
NAND_g _26549_ (.A(_04912_), .B(_04917_), .Y(_04918_));
NAND_g _26550_ (.A(_04908_), .B(_04918_), .Y(_04919_));
NAND_g _26551_ (.A(_00012_[3]), .B(_04919_), .Y(_04920_));
AND_g _26552_ (.A(_04898_), .B(_04920_), .Y(_04921_));
NAND_g _26553_ (.A(_11216_), .B(_04921_), .Y(_04922_));
NAND_g _26554_ (.A(cpuregs_20[0]), .B(_11213_), .Y(_04923_));
NAND_g _26555_ (.A(cpuregs_22[0]), .B(_00012_[1]), .Y(_04924_));
AND_g _26556_ (.A(_00012_[2]), .B(_04924_), .Y(_04925_));
NAND_g _26557_ (.A(_04923_), .B(_04925_), .Y(_04926_));
NAND_g _26558_ (.A(cpuregs_16[0]), .B(_11213_), .Y(_04927_));
NAND_g _26559_ (.A(cpuregs_18[0]), .B(_00012_[1]), .Y(_04928_));
AND_g _26560_ (.A(_11214_), .B(_04928_), .Y(_04929_));
NAND_g _26561_ (.A(_04927_), .B(_04929_), .Y(_04930_));
AND_g _26562_ (.A(_11212_), .B(_04930_), .Y(_04931_));
NAND_g _26563_ (.A(_04926_), .B(_04931_), .Y(_04932_));
NAND_g _26564_ (.A(cpuregs_21[0]), .B(_11213_), .Y(_04933_));
NAND_g _26565_ (.A(cpuregs_23[0]), .B(_00012_[1]), .Y(_04934_));
AND_g _26566_ (.A(_00012_[2]), .B(_04934_), .Y(_04935_));
NAND_g _26567_ (.A(_04933_), .B(_04935_), .Y(_04936_));
NAND_g _26568_ (.A(cpuregs_17[0]), .B(_11213_), .Y(_04937_));
NAND_g _26569_ (.A(cpuregs_19[0]), .B(_00012_[1]), .Y(_04938_));
AND_g _26570_ (.A(_11214_), .B(_04938_), .Y(_04939_));
NAND_g _26571_ (.A(_04937_), .B(_04939_), .Y(_04940_));
AND_g _26572_ (.A(_00012_[0]), .B(_04940_), .Y(_04941_));
NAND_g _26573_ (.A(_04936_), .B(_04941_), .Y(_04942_));
NAND_g _26574_ (.A(_04932_), .B(_04942_), .Y(_04943_));
NAND_g _26575_ (.A(_11215_), .B(_04943_), .Y(_04944_));
NAND_g _26576_ (.A(cpuregs_26[0]), .B(_11214_), .Y(_04945_));
NAND_g _26577_ (.A(cpuregs_30[0]), .B(_00012_[2]), .Y(_04946_));
AND_g _26578_ (.A(_00012_[1]), .B(_04946_), .Y(_04947_));
NAND_g _26579_ (.A(_04945_), .B(_04947_), .Y(_04948_));
NAND_g _26580_ (.A(cpuregs_24[0]), .B(_11214_), .Y(_04949_));
NAND_g _26581_ (.A(cpuregs_28[0]), .B(_00012_[2]), .Y(_04950_));
AND_g _26582_ (.A(_11213_), .B(_04950_), .Y(_04951_));
NAND_g _26583_ (.A(_04949_), .B(_04951_), .Y(_04952_));
AND_g _26584_ (.A(_11212_), .B(_04952_), .Y(_04953_));
NAND_g _26585_ (.A(_04948_), .B(_04953_), .Y(_04954_));
NAND_g _26586_ (.A(cpuregs_27[0]), .B(_11214_), .Y(_04955_));
NAND_g _26587_ (.A(cpuregs_31[0]), .B(_00012_[2]), .Y(_04956_));
AND_g _26588_ (.A(_00012_[1]), .B(_04956_), .Y(_04957_));
NAND_g _26589_ (.A(_04955_), .B(_04957_), .Y(_04958_));
NAND_g _26590_ (.A(cpuregs_29[0]), .B(_00012_[2]), .Y(_04959_));
NAND_g _26591_ (.A(cpuregs_25[0]), .B(_11214_), .Y(_04960_));
AND_g _26592_ (.A(_11213_), .B(_04960_), .Y(_04961_));
NAND_g _26593_ (.A(_04959_), .B(_04961_), .Y(_04962_));
AND_g _26594_ (.A(_00012_[0]), .B(_04962_), .Y(_04963_));
NAND_g _26595_ (.A(_04958_), .B(_04963_), .Y(_04964_));
NAND_g _26596_ (.A(_04954_), .B(_04964_), .Y(_04965_));
NAND_g _26597_ (.A(_00012_[3]), .B(_04965_), .Y(_04966_));
AND_g _26598_ (.A(_00012_[4]), .B(_04944_), .Y(_04967_));
NAND_g _26599_ (.A(_04966_), .B(_04967_), .Y(_04968_));
AND_g _26600_ (.A(_13409_), .B(_04968_), .Y(_04969_));
AND_g _26601_ (.A(_04922_), .B(_04969_), .Y(_04970_));
AND_g _26602_ (.A(_13613_), .B(_04970_), .Y(_04971_));
XOR_g _26603_ (.A(decoded_imm[0]), .B(pcpi_rs1[0]), .Y(_04972_));
NAND_g _26604_ (.A(_13432_), .B(_04972_), .Y(_04973_));
NAND_g _26605_ (.A(reg_next_pc[0]), .B(_13714_), .Y(_04974_));
AND_g _26606_ (.A(_11136_), .B(_13382_), .Y(_04975_));
NOR_g _26607_ (.A(pcpi_rs1[4]), .B(_13382_), .Y(_04976_));
NOR_g _26608_ (.A(_04975_), .B(_04976_), .Y(_04977_));
AND_g _26609_ (.A(_13419_), .B(_04977_), .Y(_04978_));
NAND_g _26610_ (.A(_13389_), .B(_04978_), .Y(_04979_));
AND_g _26611_ (.A(_04974_), .B(_04979_), .Y(_04980_));
AND_g _26612_ (.A(_04973_), .B(_04980_), .Y(_04981_));
NAND_g _26613_ (.A(_13425_), .B(_04981_), .Y(_04982_));
NOR_g _26614_ (.A(_04971_), .B(_04982_), .Y(_04983_));
NOR_g _26615_ (.A(_04876_), .B(_04983_), .Y(_01207_));
NOR_g _26616_ (.A(pcpi_rs1[1]), .B(_13425_), .Y(_04984_));
NAND_g _26617_ (.A(cpuregs_7[1]), .B(_00012_[2]), .Y(_04985_));
NAND_g _26618_ (.A(cpuregs_3[1]), .B(_11214_), .Y(_04986_));
NAND_g _26619_ (.A(_04985_), .B(_04986_), .Y(_04987_));
AND_g _26620_ (.A(_00012_[0]), .B(_04987_), .Y(_04988_));
NAND_g _26621_ (.A(cpuregs_6[1]), .B(_00012_[2]), .Y(_04989_));
NAND_g _26622_ (.A(cpuregs_2[1]), .B(_11214_), .Y(_04990_));
AND_g _26623_ (.A(_04989_), .B(_04990_), .Y(_04991_));
NOR_g _26624_ (.A(_00012_[0]), .B(_04991_), .Y(_04992_));
NOR_g _26625_ (.A(_04988_), .B(_04992_), .Y(_04993_));
NAND_g _26626_ (.A(cpuregs_5[1]), .B(_00012_[2]), .Y(_04994_));
NAND_g _26627_ (.A(cpuregs_1[1]), .B(_11214_), .Y(_04995_));
NAND_g _26628_ (.A(_04994_), .B(_04995_), .Y(_04996_));
NAND_g _26629_ (.A(_00012_[0]), .B(_04996_), .Y(_04997_));
NAND_g _26630_ (.A(cpuregs_4[1]), .B(_00012_[2]), .Y(_04998_));
NAND_g _26631_ (.A(cpuregs_0[1]), .B(_11214_), .Y(_04999_));
AND_g _26632_ (.A(_04998_), .B(_04999_), .Y(_05000_));
NOR_g _26633_ (.A(_00012_[0]), .B(_05000_), .Y(_05001_));
NAND_g _26634_ (.A(_00012_[1]), .B(_04993_), .Y(_05002_));
NOR_g _26635_ (.A(_00012_[1]), .B(_05001_), .Y(_05003_));
NAND_g _26636_ (.A(_04997_), .B(_05003_), .Y(_05004_));
AND_g _26637_ (.A(_05002_), .B(_05004_), .Y(_05005_));
NAND_g _26638_ (.A(_11215_), .B(_05005_), .Y(_05006_));
NAND_g _26639_ (.A(cpuregs_13[1]), .B(_00012_[0]), .Y(_05007_));
NAND_g _26640_ (.A(cpuregs_12[1]), .B(_11212_), .Y(_05008_));
AND_g _26641_ (.A(_00012_[2]), .B(_05008_), .Y(_05009_));
NAND_g _26642_ (.A(_05007_), .B(_05009_), .Y(_05010_));
NAND_g _26643_ (.A(cpuregs_9[1]), .B(_00012_[0]), .Y(_05011_));
NAND_g _26644_ (.A(cpuregs_8[1]), .B(_11212_), .Y(_05012_));
AND_g _26645_ (.A(_11214_), .B(_05012_), .Y(_05013_));
NAND_g _26646_ (.A(_05011_), .B(_05013_), .Y(_05014_));
AND_g _26647_ (.A(_11213_), .B(_05014_), .Y(_05015_));
NAND_g _26648_ (.A(_05010_), .B(_05015_), .Y(_05016_));
NAND_g _26649_ (.A(cpuregs_15[1]), .B(_00012_[0]), .Y(_05017_));
NAND_g _26650_ (.A(cpuregs_14[1]), .B(_11212_), .Y(_05018_));
AND_g _26651_ (.A(_00012_[2]), .B(_05018_), .Y(_05019_));
NAND_g _26652_ (.A(_05017_), .B(_05019_), .Y(_05020_));
NAND_g _26653_ (.A(cpuregs_11[1]), .B(_00012_[0]), .Y(_05021_));
NAND_g _26654_ (.A(cpuregs_10[1]), .B(_11212_), .Y(_05022_));
AND_g _26655_ (.A(_11214_), .B(_05022_), .Y(_05023_));
NAND_g _26656_ (.A(_05021_), .B(_05023_), .Y(_05024_));
AND_g _26657_ (.A(_00012_[1]), .B(_05024_), .Y(_05025_));
NAND_g _26658_ (.A(_05020_), .B(_05025_), .Y(_05026_));
NAND_g _26659_ (.A(_05016_), .B(_05026_), .Y(_05027_));
NAND_g _26660_ (.A(_00012_[3]), .B(_05027_), .Y(_05028_));
AND_g _26661_ (.A(_05006_), .B(_05028_), .Y(_05029_));
NAND_g _26662_ (.A(_11216_), .B(_05029_), .Y(_05030_));
NAND_g _26663_ (.A(_11014_), .B(_00012_[2]), .Y(_05031_));
NOR_g _26664_ (.A(cpuregs_18[1]), .B(_00012_[2]), .Y(_05032_));
NOR_g _26665_ (.A(_00012_[0]), .B(_05032_), .Y(_05033_));
NAND_g _26666_ (.A(_05031_), .B(_05033_), .Y(_05034_));
NAND_g _26667_ (.A(_11177_), .B(_00012_[2]), .Y(_05035_));
NOR_g _26668_ (.A(cpuregs_19[1]), .B(_00012_[2]), .Y(_05036_));
NOR_g _26669_ (.A(_11212_), .B(_05036_), .Y(_05037_));
NAND_g _26670_ (.A(_05035_), .B(_05037_), .Y(_05038_));
AND_g _26671_ (.A(_05034_), .B(_05038_), .Y(_05039_));
NAND_g _26672_ (.A(_11193_), .B(_00012_[2]), .Y(_05040_));
NOR_g _26673_ (.A(cpuregs_16[1]), .B(_00012_[2]), .Y(_05041_));
NOR_g _26674_ (.A(_00012_[0]), .B(_05041_), .Y(_05042_));
NAND_g _26675_ (.A(_05040_), .B(_05042_), .Y(_05043_));
NAND_g _26676_ (.A(_11022_), .B(_00012_[2]), .Y(_05044_));
NOR_g _26677_ (.A(cpuregs_17[1]), .B(_00012_[2]), .Y(_05045_));
NOR_g _26678_ (.A(_11212_), .B(_05045_), .Y(_05046_));
NAND_g _26679_ (.A(_05044_), .B(_05046_), .Y(_05047_));
AND_g _26680_ (.A(_05043_), .B(_05047_), .Y(_05048_));
NAND_g _26681_ (.A(_00012_[1]), .B(_05039_), .Y(_05049_));
NAND_g _26682_ (.A(_11213_), .B(_05048_), .Y(_05050_));
AND_g _26683_ (.A(_05049_), .B(_05050_), .Y(_05051_));
NAND_g _26684_ (.A(_11215_), .B(_05051_), .Y(_05052_));
NAND_g _26685_ (.A(cpuregs_29[1]), .B(_11213_), .Y(_05053_));
NAND_g _26686_ (.A(cpuregs_31[1]), .B(_00012_[1]), .Y(_05054_));
AND_g _26687_ (.A(_00012_[2]), .B(_05054_), .Y(_05055_));
NAND_g _26688_ (.A(_05053_), .B(_05055_), .Y(_05056_));
NAND_g _26689_ (.A(cpuregs_25[1]), .B(_11213_), .Y(_05057_));
NAND_g _26690_ (.A(cpuregs_27[1]), .B(_00012_[1]), .Y(_05058_));
AND_g _26691_ (.A(_11214_), .B(_05058_), .Y(_05059_));
NAND_g _26692_ (.A(_05057_), .B(_05059_), .Y(_05060_));
AND_g _26693_ (.A(_00012_[0]), .B(_05060_), .Y(_05061_));
NAND_g _26694_ (.A(_05056_), .B(_05061_), .Y(_05062_));
NAND_g _26695_ (.A(cpuregs_28[1]), .B(_11213_), .Y(_05063_));
NAND_g _26696_ (.A(cpuregs_30[1]), .B(_00012_[1]), .Y(_05064_));
AND_g _26697_ (.A(_00012_[2]), .B(_05064_), .Y(_05065_));
NAND_g _26698_ (.A(_05063_), .B(_05065_), .Y(_05066_));
NAND_g _26699_ (.A(cpuregs_24[1]), .B(_11213_), .Y(_05067_));
NAND_g _26700_ (.A(cpuregs_26[1]), .B(_00012_[1]), .Y(_05068_));
AND_g _26701_ (.A(_11214_), .B(_05068_), .Y(_05069_));
NAND_g _26702_ (.A(_05067_), .B(_05069_), .Y(_05070_));
AND_g _26703_ (.A(_11212_), .B(_05070_), .Y(_05071_));
NAND_g _26704_ (.A(_05066_), .B(_05071_), .Y(_05072_));
NAND_g _26705_ (.A(_05062_), .B(_05072_), .Y(_05073_));
NAND_g _26706_ (.A(_00012_[3]), .B(_05073_), .Y(_05074_));
AND_g _26707_ (.A(_05052_), .B(_05074_), .Y(_05075_));
NAND_g _26708_ (.A(_00012_[4]), .B(_05075_), .Y(_05076_));
AND_g _26709_ (.A(_13409_), .B(_05076_), .Y(_05077_));
AND_g _26710_ (.A(_05030_), .B(_05077_), .Y(_05078_));
AND_g _26711_ (.A(_13613_), .B(_05078_), .Y(_05079_));
XOR_g _26712_ (.A(_13489_), .B(_13490_), .Y(_05080_));
NAND_g _26713_ (.A(_13432_), .B(_05080_), .Y(_05081_));
NAND_g _26714_ (.A(reg_pc[1]), .B(_13714_), .Y(_05082_));
NAND_g _26715_ (.A(pcpi_rs1[0]), .B(_13420_), .Y(_05083_));
NAND_g _26716_ (.A(pcpi_rs1[2]), .B(_13419_), .Y(_05084_));
NAND_g _26717_ (.A(pcpi_rs1[5]), .B(_13419_), .Y(_05085_));
NAND_g _26718_ (.A(_13383_), .B(_05085_), .Y(_05086_));
AND_g _26719_ (.A(_13382_), .B(_05084_), .Y(_05087_));
NAND_g _26720_ (.A(_05083_), .B(_05087_), .Y(_05088_));
AND_g _26721_ (.A(_05086_), .B(_05088_), .Y(_05089_));
NAND_g _26722_ (.A(_13389_), .B(_05089_), .Y(_05090_));
AND_g _26723_ (.A(_05082_), .B(_05090_), .Y(_05091_));
AND_g _26724_ (.A(_05081_), .B(_05091_), .Y(_05092_));
NAND_g _26725_ (.A(_13425_), .B(_05092_), .Y(_05093_));
NOR_g _26726_ (.A(_05079_), .B(_05093_), .Y(_05094_));
NOR_g _26727_ (.A(_04984_), .B(_05094_), .Y(_01208_));
NOR_g _26728_ (.A(pcpi_rs1[2]), .B(_13425_), .Y(_05095_));
NAND_g _26729_ (.A(cpuregs_13[2]), .B(_00012_[2]), .Y(_05096_));
NAND_g _26730_ (.A(cpuregs_9[2]), .B(_11214_), .Y(_05097_));
NAND_g _26731_ (.A(_05096_), .B(_05097_), .Y(_05098_));
NAND_g _26732_ (.A(_00012_[0]), .B(_05098_), .Y(_05099_));
NAND_g _26733_ (.A(cpuregs_12[2]), .B(_00012_[2]), .Y(_05100_));
NAND_g _26734_ (.A(cpuregs_8[2]), .B(_11214_), .Y(_05101_));
AND_g _26735_ (.A(_05100_), .B(_05101_), .Y(_05102_));
NOR_g _26736_ (.A(_00012_[0]), .B(_05102_), .Y(_05103_));
NAND_g _26737_ (.A(_10949_), .B(_00012_[2]), .Y(_05104_));
NOR_g _26738_ (.A(cpuregs_0[2]), .B(_00012_[2]), .Y(_05105_));
NOR_g _26739_ (.A(_00012_[0]), .B(_05105_), .Y(_05106_));
NAND_g _26740_ (.A(_05104_), .B(_05106_), .Y(_05107_));
NAND_g _26741_ (.A(_11107_), .B(_00012_[2]), .Y(_05108_));
NOR_g _26742_ (.A(cpuregs_1[2]), .B(_00012_[2]), .Y(_05109_));
NOR_g _26743_ (.A(_11212_), .B(_05109_), .Y(_05110_));
NAND_g _26744_ (.A(_05108_), .B(_05110_), .Y(_05111_));
NAND_g _26745_ (.A(cpuregs_11[2]), .B(_11214_), .Y(_05112_));
NAND_g _26746_ (.A(cpuregs_15[2]), .B(_00012_[2]), .Y(_05113_));
NAND_g _26747_ (.A(_05112_), .B(_05113_), .Y(_05114_));
AND_g _26748_ (.A(_00012_[0]), .B(_05114_), .Y(_05115_));
NAND_g _26749_ (.A(cpuregs_14[2]), .B(_00012_[2]), .Y(_05116_));
NAND_g _26750_ (.A(cpuregs_10[2]), .B(_11214_), .Y(_05117_));
AND_g _26751_ (.A(_05116_), .B(_05117_), .Y(_05118_));
NOR_g _26752_ (.A(_00012_[0]), .B(_05118_), .Y(_05119_));
NOR_g _26753_ (.A(_05115_), .B(_05119_), .Y(_05120_));
NAND_g _26754_ (.A(_10937_), .B(_00012_[2]), .Y(_05121_));
NOR_g _26755_ (.A(cpuregs_2[2]), .B(_00012_[2]), .Y(_05122_));
NOR_g _26756_ (.A(_00012_[0]), .B(_05122_), .Y(_05123_));
NAND_g _26757_ (.A(_05121_), .B(_05123_), .Y(_05124_));
NAND_g _26758_ (.A(_11123_), .B(_00012_[2]), .Y(_05125_));
NOR_g _26759_ (.A(cpuregs_3[2]), .B(_00012_[2]), .Y(_05126_));
NOR_g _26760_ (.A(_11212_), .B(_05126_), .Y(_05127_));
NAND_g _26761_ (.A(_05125_), .B(_05127_), .Y(_05128_));
AND_g _26762_ (.A(_05124_), .B(_05128_), .Y(_05129_));
NAND_g _26763_ (.A(_00012_[1]), .B(_05129_), .Y(_05130_));
AND_g _26764_ (.A(_11213_), .B(_05107_), .Y(_05131_));
NAND_g _26765_ (.A(_05111_), .B(_05131_), .Y(_05132_));
AND_g _26766_ (.A(_05130_), .B(_05132_), .Y(_05133_));
NAND_g _26767_ (.A(_11215_), .B(_05133_), .Y(_05134_));
NAND_g _26768_ (.A(_00012_[1]), .B(_05120_), .Y(_05135_));
NOR_g _26769_ (.A(_00012_[1]), .B(_05103_), .Y(_05136_));
NAND_g _26770_ (.A(_05099_), .B(_05136_), .Y(_05137_));
AND_g _26771_ (.A(_00012_[3]), .B(_05137_), .Y(_05138_));
NAND_g _26772_ (.A(_05135_), .B(_05138_), .Y(_05139_));
AND_g _26773_ (.A(_05134_), .B(_05139_), .Y(_05140_));
NAND_g _26774_ (.A(_11216_), .B(_05140_), .Y(_05141_));
NAND_g _26775_ (.A(cpuregs_20[2]), .B(_11213_), .Y(_05142_));
NAND_g _26776_ (.A(cpuregs_22[2]), .B(_00012_[1]), .Y(_05143_));
AND_g _26777_ (.A(_00012_[2]), .B(_05143_), .Y(_05144_));
NAND_g _26778_ (.A(_05142_), .B(_05144_), .Y(_05145_));
NAND_g _26779_ (.A(cpuregs_16[2]), .B(_11213_), .Y(_05146_));
NAND_g _26780_ (.A(cpuregs_18[2]), .B(_00012_[1]), .Y(_05147_));
AND_g _26781_ (.A(_11214_), .B(_05147_), .Y(_05148_));
NAND_g _26782_ (.A(_05146_), .B(_05148_), .Y(_05149_));
AND_g _26783_ (.A(_11212_), .B(_05149_), .Y(_05150_));
NAND_g _26784_ (.A(_05145_), .B(_05150_), .Y(_05151_));
NAND_g _26785_ (.A(cpuregs_21[2]), .B(_11213_), .Y(_05152_));
NAND_g _26786_ (.A(cpuregs_23[2]), .B(_00012_[1]), .Y(_05153_));
AND_g _26787_ (.A(_00012_[2]), .B(_05153_), .Y(_05154_));
NAND_g _26788_ (.A(_05152_), .B(_05154_), .Y(_05155_));
NAND_g _26789_ (.A(cpuregs_17[2]), .B(_11213_), .Y(_05156_));
NAND_g _26790_ (.A(cpuregs_19[2]), .B(_00012_[1]), .Y(_05157_));
AND_g _26791_ (.A(_11214_), .B(_05157_), .Y(_05158_));
NAND_g _26792_ (.A(_05156_), .B(_05158_), .Y(_05159_));
AND_g _26793_ (.A(_00012_[0]), .B(_05159_), .Y(_05160_));
NAND_g _26794_ (.A(_05155_), .B(_05160_), .Y(_05161_));
NAND_g _26795_ (.A(_05151_), .B(_05161_), .Y(_05162_));
NAND_g _26796_ (.A(_11215_), .B(_05162_), .Y(_05163_));
NAND_g _26797_ (.A(cpuregs_26[2]), .B(_11214_), .Y(_05164_));
NAND_g _26798_ (.A(cpuregs_30[2]), .B(_00012_[2]), .Y(_05165_));
AND_g _26799_ (.A(_00012_[1]), .B(_05165_), .Y(_05166_));
NAND_g _26800_ (.A(_05164_), .B(_05166_), .Y(_05167_));
NAND_g _26801_ (.A(cpuregs_24[2]), .B(_11214_), .Y(_05168_));
NAND_g _26802_ (.A(cpuregs_28[2]), .B(_00012_[2]), .Y(_05169_));
AND_g _26803_ (.A(_11213_), .B(_05169_), .Y(_05170_));
NAND_g _26804_ (.A(_05168_), .B(_05170_), .Y(_05171_));
AND_g _26805_ (.A(_11212_), .B(_05171_), .Y(_05172_));
NAND_g _26806_ (.A(_05167_), .B(_05172_), .Y(_05173_));
NAND_g _26807_ (.A(cpuregs_27[2]), .B(_11214_), .Y(_05174_));
NAND_g _26808_ (.A(cpuregs_31[2]), .B(_00012_[2]), .Y(_05175_));
AND_g _26809_ (.A(_00012_[1]), .B(_05175_), .Y(_05176_));
NAND_g _26810_ (.A(_05174_), .B(_05176_), .Y(_05177_));
NAND_g _26811_ (.A(cpuregs_29[2]), .B(_00012_[2]), .Y(_05178_));
NAND_g _26812_ (.A(cpuregs_25[2]), .B(_11214_), .Y(_05179_));
AND_g _26813_ (.A(_11213_), .B(_05179_), .Y(_05180_));
NAND_g _26814_ (.A(_05178_), .B(_05180_), .Y(_05181_));
AND_g _26815_ (.A(_00012_[0]), .B(_05181_), .Y(_05182_));
NAND_g _26816_ (.A(_05177_), .B(_05182_), .Y(_05183_));
NAND_g _26817_ (.A(_05173_), .B(_05183_), .Y(_05184_));
NAND_g _26818_ (.A(_00012_[3]), .B(_05184_), .Y(_05185_));
AND_g _26819_ (.A(_00012_[4]), .B(_05163_), .Y(_05186_));
NAND_g _26820_ (.A(_05185_), .B(_05186_), .Y(_05187_));
AND_g _26821_ (.A(_13409_), .B(_05187_), .Y(_05188_));
AND_g _26822_ (.A(_05141_), .B(_05188_), .Y(_05189_));
AND_g _26823_ (.A(_13613_), .B(_05189_), .Y(_05190_));
XOR_g _26824_ (.A(_13492_), .B(_13493_), .Y(_05191_));
NAND_g _26825_ (.A(_13432_), .B(_05191_), .Y(_05192_));
NAND_g _26826_ (.A(reg_pc[2]), .B(_13714_), .Y(_05193_));
NAND_g _26827_ (.A(pcpi_rs1[1]), .B(_13420_), .Y(_05194_));
NAND_g _26828_ (.A(pcpi_rs1[3]), .B(_13419_), .Y(_05195_));
NAND_g _26829_ (.A(pcpi_rs1[6]), .B(_13419_), .Y(_05196_));
NAND_g _26830_ (.A(_13383_), .B(_05196_), .Y(_05197_));
AND_g _26831_ (.A(_13382_), .B(_05195_), .Y(_05198_));
NAND_g _26832_ (.A(_05194_), .B(_05198_), .Y(_05199_));
AND_g _26833_ (.A(_05197_), .B(_05199_), .Y(_05200_));
NAND_g _26834_ (.A(_13389_), .B(_05200_), .Y(_05201_));
AND_g _26835_ (.A(_05193_), .B(_05201_), .Y(_05202_));
AND_g _26836_ (.A(_05192_), .B(_05202_), .Y(_05203_));
NAND_g _26837_ (.A(_13425_), .B(_05203_), .Y(_05204_));
NOR_g _26838_ (.A(_05190_), .B(_05204_), .Y(_05205_));
NOR_g _26839_ (.A(_05095_), .B(_05205_), .Y(_01209_));
NOR_g _26840_ (.A(pcpi_rs1[3]), .B(_13425_), .Y(_05206_));
NAND_g _26841_ (.A(cpuregs_13[3]), .B(_00012_[2]), .Y(_05207_));
NAND_g _26842_ (.A(cpuregs_9[3]), .B(_11214_), .Y(_05208_));
NAND_g _26843_ (.A(_05207_), .B(_05208_), .Y(_05209_));
NAND_g _26844_ (.A(_00012_[0]), .B(_05209_), .Y(_05210_));
NAND_g _26845_ (.A(cpuregs_12[3]), .B(_00012_[2]), .Y(_05211_));
NAND_g _26846_ (.A(cpuregs_8[3]), .B(_11214_), .Y(_05212_));
AND_g _26847_ (.A(_05211_), .B(_05212_), .Y(_05213_));
NOR_g _26848_ (.A(_00012_[0]), .B(_05213_), .Y(_05214_));
NAND_g _26849_ (.A(_10950_), .B(_00012_[2]), .Y(_05215_));
NOR_g _26850_ (.A(cpuregs_0[3]), .B(_00012_[2]), .Y(_05216_));
NOR_g _26851_ (.A(_00012_[0]), .B(_05216_), .Y(_05217_));
NAND_g _26852_ (.A(_05215_), .B(_05217_), .Y(_05218_));
NAND_g _26853_ (.A(_11108_), .B(_00012_[2]), .Y(_05219_));
NOR_g _26854_ (.A(cpuregs_1[3]), .B(_00012_[2]), .Y(_05220_));
NOR_g _26855_ (.A(_11212_), .B(_05220_), .Y(_05221_));
NAND_g _26856_ (.A(_05219_), .B(_05221_), .Y(_05222_));
NAND_g _26857_ (.A(cpuregs_11[3]), .B(_11214_), .Y(_05223_));
NAND_g _26858_ (.A(cpuregs_15[3]), .B(_00012_[2]), .Y(_05224_));
NAND_g _26859_ (.A(_05223_), .B(_05224_), .Y(_05225_));
AND_g _26860_ (.A(_00012_[0]), .B(_05225_), .Y(_05226_));
NAND_g _26861_ (.A(cpuregs_14[3]), .B(_00012_[2]), .Y(_05227_));
NAND_g _26862_ (.A(cpuregs_10[3]), .B(_11214_), .Y(_05228_));
AND_g _26863_ (.A(_05227_), .B(_05228_), .Y(_05229_));
NOR_g _26864_ (.A(_00012_[0]), .B(_05229_), .Y(_05230_));
NOR_g _26865_ (.A(_05226_), .B(_05230_), .Y(_05231_));
NAND_g _26866_ (.A(_10938_), .B(_00012_[2]), .Y(_05232_));
NOR_g _26867_ (.A(cpuregs_2[3]), .B(_00012_[2]), .Y(_05233_));
NOR_g _26868_ (.A(_00012_[0]), .B(_05233_), .Y(_05234_));
NAND_g _26869_ (.A(_05232_), .B(_05234_), .Y(_05235_));
NAND_g _26870_ (.A(_11124_), .B(_00012_[2]), .Y(_05236_));
NOR_g _26871_ (.A(cpuregs_3[3]), .B(_00012_[2]), .Y(_05237_));
NOR_g _26872_ (.A(_11212_), .B(_05237_), .Y(_05238_));
NAND_g _26873_ (.A(_05236_), .B(_05238_), .Y(_05239_));
AND_g _26874_ (.A(_05235_), .B(_05239_), .Y(_05240_));
NAND_g _26875_ (.A(_00012_[1]), .B(_05240_), .Y(_05241_));
AND_g _26876_ (.A(_11213_), .B(_05218_), .Y(_05242_));
NAND_g _26877_ (.A(_05222_), .B(_05242_), .Y(_05243_));
AND_g _26878_ (.A(_05241_), .B(_05243_), .Y(_05244_));
NAND_g _26879_ (.A(_11215_), .B(_05244_), .Y(_05245_));
NAND_g _26880_ (.A(_00012_[1]), .B(_05231_), .Y(_05246_));
NOR_g _26881_ (.A(_00012_[1]), .B(_05214_), .Y(_05247_));
NAND_g _26882_ (.A(_05210_), .B(_05247_), .Y(_05248_));
AND_g _26883_ (.A(_00012_[3]), .B(_05248_), .Y(_05249_));
NAND_g _26884_ (.A(_05246_), .B(_05249_), .Y(_05250_));
AND_g _26885_ (.A(_05245_), .B(_05250_), .Y(_05251_));
NAND_g _26886_ (.A(_11216_), .B(_05251_), .Y(_05252_));
NAND_g _26887_ (.A(cpuregs_20[3]), .B(_11213_), .Y(_05253_));
NAND_g _26888_ (.A(cpuregs_22[3]), .B(_00012_[1]), .Y(_05254_));
AND_g _26889_ (.A(_00012_[2]), .B(_05254_), .Y(_05255_));
NAND_g _26890_ (.A(_05253_), .B(_05255_), .Y(_05256_));
NAND_g _26891_ (.A(cpuregs_16[3]), .B(_11213_), .Y(_05257_));
NAND_g _26892_ (.A(cpuregs_18[3]), .B(_00012_[1]), .Y(_05258_));
AND_g _26893_ (.A(_11214_), .B(_05258_), .Y(_05259_));
NAND_g _26894_ (.A(_05257_), .B(_05259_), .Y(_05260_));
AND_g _26895_ (.A(_11212_), .B(_05260_), .Y(_05261_));
NAND_g _26896_ (.A(_05256_), .B(_05261_), .Y(_05262_));
NAND_g _26897_ (.A(cpuregs_21[3]), .B(_11213_), .Y(_05263_));
NAND_g _26898_ (.A(cpuregs_23[3]), .B(_00012_[1]), .Y(_05264_));
AND_g _26899_ (.A(_00012_[2]), .B(_05264_), .Y(_05265_));
NAND_g _26900_ (.A(_05263_), .B(_05265_), .Y(_05266_));
NAND_g _26901_ (.A(cpuregs_17[3]), .B(_11213_), .Y(_05267_));
NAND_g _26902_ (.A(cpuregs_19[3]), .B(_00012_[1]), .Y(_05268_));
AND_g _26903_ (.A(_11214_), .B(_05268_), .Y(_05269_));
NAND_g _26904_ (.A(_05267_), .B(_05269_), .Y(_05270_));
AND_g _26905_ (.A(_00012_[0]), .B(_05270_), .Y(_05271_));
NAND_g _26906_ (.A(_05266_), .B(_05271_), .Y(_05272_));
NAND_g _26907_ (.A(_05262_), .B(_05272_), .Y(_05273_));
NAND_g _26908_ (.A(_11215_), .B(_05273_), .Y(_05274_));
NAND_g _26909_ (.A(cpuregs_26[3]), .B(_11214_), .Y(_05275_));
NAND_g _26910_ (.A(cpuregs_30[3]), .B(_00012_[2]), .Y(_05276_));
AND_g _26911_ (.A(_00012_[1]), .B(_05276_), .Y(_05277_));
NAND_g _26912_ (.A(_05275_), .B(_05277_), .Y(_05278_));
NAND_g _26913_ (.A(cpuregs_24[3]), .B(_11214_), .Y(_05279_));
NAND_g _26914_ (.A(cpuregs_28[3]), .B(_00012_[2]), .Y(_05280_));
AND_g _26915_ (.A(_11213_), .B(_05280_), .Y(_05281_));
NAND_g _26916_ (.A(_05279_), .B(_05281_), .Y(_05282_));
AND_g _26917_ (.A(_11212_), .B(_05282_), .Y(_05283_));
NAND_g _26918_ (.A(_05278_), .B(_05283_), .Y(_05284_));
NAND_g _26919_ (.A(cpuregs_27[3]), .B(_11214_), .Y(_05285_));
NAND_g _26920_ (.A(cpuregs_31[3]), .B(_00012_[2]), .Y(_05286_));
AND_g _26921_ (.A(_00012_[1]), .B(_05286_), .Y(_05287_));
NAND_g _26922_ (.A(_05285_), .B(_05287_), .Y(_05288_));
NAND_g _26923_ (.A(cpuregs_29[3]), .B(_00012_[2]), .Y(_05289_));
NAND_g _26924_ (.A(cpuregs_25[3]), .B(_11214_), .Y(_05290_));
AND_g _26925_ (.A(_11213_), .B(_05290_), .Y(_05291_));
NAND_g _26926_ (.A(_05289_), .B(_05291_), .Y(_05292_));
AND_g _26927_ (.A(_00012_[0]), .B(_05292_), .Y(_05293_));
NAND_g _26928_ (.A(_05288_), .B(_05293_), .Y(_05294_));
NAND_g _26929_ (.A(_05284_), .B(_05294_), .Y(_05295_));
NAND_g _26930_ (.A(_00012_[3]), .B(_05295_), .Y(_05296_));
AND_g _26931_ (.A(_00012_[4]), .B(_05274_), .Y(_05297_));
NAND_g _26932_ (.A(_05296_), .B(_05297_), .Y(_05298_));
AND_g _26933_ (.A(_13409_), .B(_05298_), .Y(_05299_));
AND_g _26934_ (.A(_05252_), .B(_05299_), .Y(_05300_));
AND_g _26935_ (.A(_13613_), .B(_05300_), .Y(_05301_));
NAND_g _26936_ (.A(reg_pc[3]), .B(_13714_), .Y(_05302_));
NAND_g _26937_ (.A(pcpi_rs1[2]), .B(_13420_), .Y(_05303_));
NAND_g _26938_ (.A(pcpi_rs1[4]), .B(_13419_), .Y(_05304_));
NAND_g _26939_ (.A(pcpi_rs1[7]), .B(_13419_), .Y(_05305_));
AND_g _26940_ (.A(_13382_), .B(_05304_), .Y(_05306_));
NAND_g _26941_ (.A(_05303_), .B(_05306_), .Y(_05307_));
NAND_g _26942_ (.A(_13383_), .B(_05305_), .Y(_05308_));
AND_g _26943_ (.A(_05307_), .B(_05308_), .Y(_05309_));
NAND_g _26944_ (.A(_13389_), .B(_05309_), .Y(_05310_));
AND_g _26945_ (.A(_05302_), .B(_05310_), .Y(_05311_));
XOR_g _26946_ (.A(decoded_imm[3]), .B(pcpi_rs1[3]), .Y(_05312_));
XNOR_g _26947_ (.A(_13495_), .B(_05312_), .Y(_05313_));
NAND_g _26948_ (.A(_13432_), .B(_05313_), .Y(_05314_));
AND_g _26949_ (.A(_05311_), .B(_05314_), .Y(_05315_));
NAND_g _26950_ (.A(_13425_), .B(_05315_), .Y(_05316_));
NOR_g _26951_ (.A(_05301_), .B(_05316_), .Y(_05317_));
NOR_g _26952_ (.A(_05206_), .B(_05317_), .Y(_01210_));
NOR_g _26953_ (.A(pcpi_rs1[4]), .B(_13425_), .Y(_05318_));
NAND_g _26954_ (.A(cpuregs_7[4]), .B(_00012_[2]), .Y(_05319_));
NAND_g _26955_ (.A(cpuregs_3[4]), .B(_11214_), .Y(_05320_));
NAND_g _26956_ (.A(_05319_), .B(_05320_), .Y(_05321_));
AND_g _26957_ (.A(_00012_[0]), .B(_05321_), .Y(_05322_));
NAND_g _26958_ (.A(cpuregs_6[4]), .B(_00012_[2]), .Y(_05323_));
NAND_g _26959_ (.A(cpuregs_2[4]), .B(_11214_), .Y(_05324_));
AND_g _26960_ (.A(_05323_), .B(_05324_), .Y(_05325_));
NOR_g _26961_ (.A(_00012_[0]), .B(_05325_), .Y(_05326_));
NOR_g _26962_ (.A(_05322_), .B(_05326_), .Y(_05327_));
NAND_g _26963_ (.A(cpuregs_5[4]), .B(_00012_[2]), .Y(_05328_));
NAND_g _26964_ (.A(cpuregs_1[4]), .B(_11214_), .Y(_05329_));
NAND_g _26965_ (.A(_05328_), .B(_05329_), .Y(_05330_));
NAND_g _26966_ (.A(_00012_[0]), .B(_05330_), .Y(_05331_));
NAND_g _26967_ (.A(cpuregs_4[4]), .B(_00012_[2]), .Y(_05332_));
NAND_g _26968_ (.A(cpuregs_0[4]), .B(_11214_), .Y(_05333_));
AND_g _26969_ (.A(_05332_), .B(_05333_), .Y(_05334_));
NOR_g _26970_ (.A(_00012_[0]), .B(_05334_), .Y(_05335_));
NAND_g _26971_ (.A(_00012_[1]), .B(_05327_), .Y(_05336_));
NOR_g _26972_ (.A(_00012_[1]), .B(_05335_), .Y(_05337_));
NAND_g _26973_ (.A(_05331_), .B(_05337_), .Y(_05338_));
AND_g _26974_ (.A(_05336_), .B(_05338_), .Y(_05339_));
NAND_g _26975_ (.A(_11215_), .B(_05339_), .Y(_05340_));
NAND_g _26976_ (.A(cpuregs_13[4]), .B(_00012_[0]), .Y(_05341_));
NAND_g _26977_ (.A(cpuregs_12[4]), .B(_11212_), .Y(_05342_));
AND_g _26978_ (.A(_00012_[2]), .B(_05342_), .Y(_05343_));
NAND_g _26979_ (.A(_05341_), .B(_05343_), .Y(_05344_));
NAND_g _26980_ (.A(cpuregs_9[4]), .B(_00012_[0]), .Y(_05345_));
NAND_g _26981_ (.A(cpuregs_8[4]), .B(_11212_), .Y(_05346_));
AND_g _26982_ (.A(_11214_), .B(_05346_), .Y(_05347_));
NAND_g _26983_ (.A(_05345_), .B(_05347_), .Y(_05348_));
AND_g _26984_ (.A(_11213_), .B(_05348_), .Y(_05349_));
NAND_g _26985_ (.A(_05344_), .B(_05349_), .Y(_05350_));
NAND_g _26986_ (.A(cpuregs_15[4]), .B(_00012_[0]), .Y(_05351_));
NAND_g _26987_ (.A(cpuregs_14[4]), .B(_11212_), .Y(_05352_));
AND_g _26988_ (.A(_00012_[2]), .B(_05352_), .Y(_05353_));
NAND_g _26989_ (.A(_05351_), .B(_05353_), .Y(_05354_));
NAND_g _26990_ (.A(cpuregs_11[4]), .B(_00012_[0]), .Y(_05355_));
NAND_g _26991_ (.A(cpuregs_10[4]), .B(_11212_), .Y(_05356_));
AND_g _26992_ (.A(_11214_), .B(_05356_), .Y(_05357_));
NAND_g _26993_ (.A(_05355_), .B(_05357_), .Y(_05358_));
AND_g _26994_ (.A(_00012_[1]), .B(_05358_), .Y(_05359_));
NAND_g _26995_ (.A(_05354_), .B(_05359_), .Y(_05360_));
NAND_g _26996_ (.A(_05350_), .B(_05360_), .Y(_05361_));
NAND_g _26997_ (.A(_00012_[3]), .B(_05361_), .Y(_05362_));
AND_g _26998_ (.A(_05340_), .B(_05362_), .Y(_05363_));
NAND_g _26999_ (.A(_11216_), .B(_05363_), .Y(_05364_));
NAND_g _27000_ (.A(cpuregs_20[4]), .B(_11213_), .Y(_05365_));
NAND_g _27001_ (.A(cpuregs_22[4]), .B(_00012_[1]), .Y(_05366_));
AND_g _27002_ (.A(_00012_[2]), .B(_05366_), .Y(_05367_));
NAND_g _27003_ (.A(_05365_), .B(_05367_), .Y(_05368_));
NAND_g _27004_ (.A(cpuregs_16[4]), .B(_11213_), .Y(_05369_));
NAND_g _27005_ (.A(cpuregs_18[4]), .B(_00012_[1]), .Y(_05370_));
AND_g _27006_ (.A(_11214_), .B(_05370_), .Y(_05371_));
NAND_g _27007_ (.A(_05369_), .B(_05371_), .Y(_05372_));
AND_g _27008_ (.A(_11212_), .B(_05372_), .Y(_05373_));
NAND_g _27009_ (.A(_05368_), .B(_05373_), .Y(_05374_));
NAND_g _27010_ (.A(cpuregs_21[4]), .B(_11213_), .Y(_05375_));
NAND_g _27011_ (.A(cpuregs_23[4]), .B(_00012_[1]), .Y(_05376_));
AND_g _27012_ (.A(_00012_[2]), .B(_05376_), .Y(_05377_));
NAND_g _27013_ (.A(_05375_), .B(_05377_), .Y(_05378_));
NAND_g _27014_ (.A(cpuregs_17[4]), .B(_11213_), .Y(_05379_));
NAND_g _27015_ (.A(cpuregs_19[4]), .B(_00012_[1]), .Y(_05380_));
AND_g _27016_ (.A(_11214_), .B(_05380_), .Y(_05381_));
NAND_g _27017_ (.A(_05379_), .B(_05381_), .Y(_05382_));
AND_g _27018_ (.A(_00012_[0]), .B(_05382_), .Y(_05383_));
NAND_g _27019_ (.A(_05378_), .B(_05383_), .Y(_05384_));
NAND_g _27020_ (.A(_05374_), .B(_05384_), .Y(_05385_));
NAND_g _27021_ (.A(_11215_), .B(_05385_), .Y(_05386_));
NAND_g _27022_ (.A(cpuregs_26[4]), .B(_11214_), .Y(_05387_));
NAND_g _27023_ (.A(cpuregs_30[4]), .B(_00012_[2]), .Y(_05388_));
AND_g _27024_ (.A(_00012_[1]), .B(_05388_), .Y(_05389_));
NAND_g _27025_ (.A(_05387_), .B(_05389_), .Y(_05390_));
NAND_g _27026_ (.A(cpuregs_24[4]), .B(_11214_), .Y(_05391_));
NAND_g _27027_ (.A(cpuregs_28[4]), .B(_00012_[2]), .Y(_05392_));
AND_g _27028_ (.A(_11213_), .B(_05392_), .Y(_05393_));
NAND_g _27029_ (.A(_05391_), .B(_05393_), .Y(_05394_));
AND_g _27030_ (.A(_11212_), .B(_05394_), .Y(_05395_));
NAND_g _27031_ (.A(_05390_), .B(_05395_), .Y(_05396_));
NAND_g _27032_ (.A(cpuregs_27[4]), .B(_11214_), .Y(_05397_));
NAND_g _27033_ (.A(cpuregs_31[4]), .B(_00012_[2]), .Y(_05398_));
AND_g _27034_ (.A(_00012_[1]), .B(_05398_), .Y(_05399_));
NAND_g _27035_ (.A(_05397_), .B(_05399_), .Y(_05400_));
NAND_g _27036_ (.A(cpuregs_29[4]), .B(_00012_[2]), .Y(_05401_));
NAND_g _27037_ (.A(cpuregs_25[4]), .B(_11214_), .Y(_05402_));
AND_g _27038_ (.A(_11213_), .B(_05402_), .Y(_05403_));
NAND_g _27039_ (.A(_05401_), .B(_05403_), .Y(_05404_));
AND_g _27040_ (.A(_00012_[0]), .B(_05404_), .Y(_05405_));
NAND_g _27041_ (.A(_05400_), .B(_05405_), .Y(_05406_));
NAND_g _27042_ (.A(_05396_), .B(_05406_), .Y(_05407_));
NAND_g _27043_ (.A(_00012_[3]), .B(_05407_), .Y(_05408_));
AND_g _27044_ (.A(_00012_[4]), .B(_05386_), .Y(_05409_));
NAND_g _27045_ (.A(_05408_), .B(_05409_), .Y(_05410_));
AND_g _27046_ (.A(_13409_), .B(_05410_), .Y(_05411_));
AND_g _27047_ (.A(_05364_), .B(_05411_), .Y(_05412_));
AND_g _27048_ (.A(_13613_), .B(_05412_), .Y(_05413_));
XOR_g _27049_ (.A(_13484_), .B(_13497_), .Y(_05414_));
NAND_g _27050_ (.A(_13432_), .B(_05414_), .Y(_05415_));
NAND_g _27051_ (.A(reg_pc[4]), .B(_13714_), .Y(_05416_));
NAND_g _27052_ (.A(pcpi_rs1[3]), .B(_13420_), .Y(_05417_));
AND_g _27053_ (.A(_05085_), .B(_05417_), .Y(_05418_));
NAND_g _27054_ (.A(_13382_), .B(_05418_), .Y(_05419_));
NAND_g _27055_ (.A(pcpi_rs1[8]), .B(_13419_), .Y(_05420_));
AND_g _27056_ (.A(_05083_), .B(_05420_), .Y(_05421_));
NAND_g _27057_ (.A(_13383_), .B(_05421_), .Y(_05422_));
AND_g _27058_ (.A(_13389_), .B(_05419_), .Y(_05423_));
NAND_g _27059_ (.A(_05422_), .B(_05423_), .Y(_05424_));
AND_g _27060_ (.A(_05416_), .B(_05424_), .Y(_05425_));
AND_g _27061_ (.A(_05415_), .B(_05425_), .Y(_05426_));
NAND_g _27062_ (.A(_13425_), .B(_05426_), .Y(_05427_));
NOR_g _27063_ (.A(_05413_), .B(_05427_), .Y(_05428_));
NOR_g _27064_ (.A(_05318_), .B(_05428_), .Y(_01211_));
XOR_g _27065_ (.A(_13499_), .B(_13500_), .Y(_05429_));
NAND_g _27066_ (.A(_13432_), .B(_05429_), .Y(_05430_));
NAND_g _27067_ (.A(cpuregs_7[5]), .B(_00012_[2]), .Y(_05431_));
NAND_g _27068_ (.A(cpuregs_3[5]), .B(_11214_), .Y(_05432_));
NAND_g _27069_ (.A(_05431_), .B(_05432_), .Y(_05433_));
AND_g _27070_ (.A(_00012_[0]), .B(_05433_), .Y(_05434_));
NAND_g _27071_ (.A(cpuregs_6[5]), .B(_00012_[2]), .Y(_05435_));
NAND_g _27072_ (.A(cpuregs_2[5]), .B(_11214_), .Y(_05436_));
AND_g _27073_ (.A(_05435_), .B(_05436_), .Y(_05437_));
NOR_g _27074_ (.A(_00012_[0]), .B(_05437_), .Y(_05438_));
NOR_g _27075_ (.A(_05434_), .B(_05438_), .Y(_05439_));
NAND_g _27076_ (.A(cpuregs_5[5]), .B(_00012_[2]), .Y(_05440_));
NAND_g _27077_ (.A(cpuregs_1[5]), .B(_11214_), .Y(_05441_));
NAND_g _27078_ (.A(_05440_), .B(_05441_), .Y(_05442_));
NAND_g _27079_ (.A(_00012_[0]), .B(_05442_), .Y(_05443_));
NAND_g _27080_ (.A(cpuregs_4[5]), .B(_00012_[2]), .Y(_05444_));
NAND_g _27081_ (.A(cpuregs_0[5]), .B(_11214_), .Y(_05445_));
AND_g _27082_ (.A(_05444_), .B(_05445_), .Y(_05446_));
NOR_g _27083_ (.A(_00012_[0]), .B(_05446_), .Y(_05447_));
NAND_g _27084_ (.A(_00012_[1]), .B(_05439_), .Y(_05448_));
NOR_g _27085_ (.A(_00012_[1]), .B(_05447_), .Y(_05449_));
NAND_g _27086_ (.A(_05443_), .B(_05449_), .Y(_05450_));
AND_g _27087_ (.A(_05448_), .B(_05450_), .Y(_05451_));
NAND_g _27088_ (.A(_11215_), .B(_05451_), .Y(_05452_));
NAND_g _27089_ (.A(cpuregs_13[5]), .B(_00012_[0]), .Y(_05453_));
NAND_g _27090_ (.A(cpuregs_12[5]), .B(_11212_), .Y(_05454_));
AND_g _27091_ (.A(_00012_[2]), .B(_05454_), .Y(_05455_));
NAND_g _27092_ (.A(_05453_), .B(_05455_), .Y(_05456_));
NAND_g _27093_ (.A(cpuregs_9[5]), .B(_00012_[0]), .Y(_05457_));
NAND_g _27094_ (.A(cpuregs_8[5]), .B(_11212_), .Y(_05458_));
AND_g _27095_ (.A(_11214_), .B(_05458_), .Y(_05459_));
NAND_g _27096_ (.A(_05457_), .B(_05459_), .Y(_05460_));
AND_g _27097_ (.A(_11213_), .B(_05460_), .Y(_05461_));
NAND_g _27098_ (.A(_05456_), .B(_05461_), .Y(_05462_));
NAND_g _27099_ (.A(cpuregs_15[5]), .B(_00012_[0]), .Y(_05463_));
NAND_g _27100_ (.A(cpuregs_14[5]), .B(_11212_), .Y(_05464_));
AND_g _27101_ (.A(_00012_[2]), .B(_05464_), .Y(_05465_));
NAND_g _27102_ (.A(_05463_), .B(_05465_), .Y(_05466_));
NAND_g _27103_ (.A(cpuregs_11[5]), .B(_00012_[0]), .Y(_05467_));
NAND_g _27104_ (.A(cpuregs_10[5]), .B(_11212_), .Y(_05468_));
AND_g _27105_ (.A(_11214_), .B(_05468_), .Y(_05469_));
NAND_g _27106_ (.A(_05467_), .B(_05469_), .Y(_05470_));
AND_g _27107_ (.A(_00012_[1]), .B(_05470_), .Y(_05471_));
NAND_g _27108_ (.A(_05466_), .B(_05471_), .Y(_05472_));
NAND_g _27109_ (.A(_05462_), .B(_05472_), .Y(_05473_));
NAND_g _27110_ (.A(_00012_[3]), .B(_05473_), .Y(_05474_));
AND_g _27111_ (.A(_05452_), .B(_05474_), .Y(_05475_));
NAND_g _27112_ (.A(_11216_), .B(_05475_), .Y(_05476_));
NAND_g _27113_ (.A(cpuregs_20[5]), .B(_11213_), .Y(_05477_));
NAND_g _27114_ (.A(cpuregs_22[5]), .B(_00012_[1]), .Y(_05478_));
AND_g _27115_ (.A(_00012_[2]), .B(_05478_), .Y(_05479_));
NAND_g _27116_ (.A(_05477_), .B(_05479_), .Y(_05480_));
NAND_g _27117_ (.A(cpuregs_16[5]), .B(_11213_), .Y(_05481_));
NAND_g _27118_ (.A(cpuregs_18[5]), .B(_00012_[1]), .Y(_05482_));
AND_g _27119_ (.A(_11214_), .B(_05482_), .Y(_05483_));
NAND_g _27120_ (.A(_05481_), .B(_05483_), .Y(_05484_));
AND_g _27121_ (.A(_11212_), .B(_05484_), .Y(_05485_));
NAND_g _27122_ (.A(_05480_), .B(_05485_), .Y(_05486_));
NAND_g _27123_ (.A(cpuregs_21[5]), .B(_11213_), .Y(_05487_));
NAND_g _27124_ (.A(cpuregs_23[5]), .B(_00012_[1]), .Y(_05488_));
AND_g _27125_ (.A(_00012_[2]), .B(_05488_), .Y(_05489_));
NAND_g _27126_ (.A(_05487_), .B(_05489_), .Y(_05490_));
NAND_g _27127_ (.A(cpuregs_17[5]), .B(_11213_), .Y(_05491_));
NAND_g _27128_ (.A(cpuregs_19[5]), .B(_00012_[1]), .Y(_05492_));
AND_g _27129_ (.A(_11214_), .B(_05492_), .Y(_05493_));
NAND_g _27130_ (.A(_05491_), .B(_05493_), .Y(_05494_));
AND_g _27131_ (.A(_00012_[0]), .B(_05494_), .Y(_05495_));
NAND_g _27132_ (.A(_05490_), .B(_05495_), .Y(_05496_));
NAND_g _27133_ (.A(_05486_), .B(_05496_), .Y(_05497_));
NAND_g _27134_ (.A(_11215_), .B(_05497_), .Y(_05498_));
NAND_g _27135_ (.A(cpuregs_26[5]), .B(_11214_), .Y(_05499_));
NAND_g _27136_ (.A(cpuregs_30[5]), .B(_00012_[2]), .Y(_05500_));
AND_g _27137_ (.A(_00012_[1]), .B(_05500_), .Y(_05501_));
NAND_g _27138_ (.A(_05499_), .B(_05501_), .Y(_05502_));
NAND_g _27139_ (.A(cpuregs_24[5]), .B(_11214_), .Y(_05503_));
NAND_g _27140_ (.A(cpuregs_28[5]), .B(_00012_[2]), .Y(_05504_));
AND_g _27141_ (.A(_11213_), .B(_05504_), .Y(_05505_));
NAND_g _27142_ (.A(_05503_), .B(_05505_), .Y(_05506_));
AND_g _27143_ (.A(_11212_), .B(_05506_), .Y(_05507_));
NAND_g _27144_ (.A(_05502_), .B(_05507_), .Y(_05508_));
NAND_g _27145_ (.A(cpuregs_27[5]), .B(_11214_), .Y(_05509_));
NAND_g _27146_ (.A(cpuregs_31[5]), .B(_00012_[2]), .Y(_05510_));
AND_g _27147_ (.A(_00012_[1]), .B(_05510_), .Y(_05511_));
NAND_g _27148_ (.A(_05509_), .B(_05511_), .Y(_05512_));
NAND_g _27149_ (.A(cpuregs_29[5]), .B(_00012_[2]), .Y(_05513_));
NAND_g _27150_ (.A(cpuregs_25[5]), .B(_11214_), .Y(_05514_));
AND_g _27151_ (.A(_11213_), .B(_05514_), .Y(_05515_));
NAND_g _27152_ (.A(_05513_), .B(_05515_), .Y(_05516_));
AND_g _27153_ (.A(_00012_[0]), .B(_05516_), .Y(_05517_));
NAND_g _27154_ (.A(_05512_), .B(_05517_), .Y(_05518_));
NAND_g _27155_ (.A(_05508_), .B(_05518_), .Y(_05519_));
NAND_g _27156_ (.A(_00012_[3]), .B(_05519_), .Y(_05520_));
AND_g _27157_ (.A(_00012_[4]), .B(_05498_), .Y(_05521_));
NAND_g _27158_ (.A(_05520_), .B(_05521_), .Y(_05522_));
AND_g _27159_ (.A(_13409_), .B(_05522_), .Y(_05523_));
AND_g _27160_ (.A(_05476_), .B(_05523_), .Y(_05524_));
AND_g _27161_ (.A(_13613_), .B(_05524_), .Y(_05525_));
NAND_g _27162_ (.A(_13613_), .B(_05524_), .Y(_05526_));
NAND_g _27163_ (.A(reg_pc[5]), .B(_13714_), .Y(_05527_));
NAND_g _27164_ (.A(pcpi_rs1[4]), .B(_13420_), .Y(_05528_));
NAND_g _27165_ (.A(pcpi_rs1[9]), .B(_13419_), .Y(_05529_));
AND_g _27166_ (.A(_05194_), .B(_05529_), .Y(_05530_));
AND_g _27167_ (.A(_13382_), .B(_05528_), .Y(_05531_));
NAND_g _27168_ (.A(_05196_), .B(_05531_), .Y(_05532_));
NAND_g _27169_ (.A(_13383_), .B(_05530_), .Y(_05533_));
AND_g _27170_ (.A(_13389_), .B(_05532_), .Y(_05534_));
NAND_g _27171_ (.A(_05533_), .B(_05534_), .Y(_05535_));
AND_g _27172_ (.A(_05527_), .B(_05535_), .Y(_05536_));
AND_g _27173_ (.A(_05430_), .B(_05536_), .Y(_05537_));
AND_g _27174_ (.A(_13425_), .B(_05526_), .Y(_05538_));
AND_g _27175_ (.A(_05537_), .B(_05538_), .Y(_05539_));
NOR_g _27176_ (.A(pcpi_rs1[5]), .B(_13425_), .Y(_05540_));
NOR_g _27177_ (.A(_05539_), .B(_05540_), .Y(_01212_));
NOR_g _27178_ (.A(cpuregs_9[6]), .B(_00012_[2]), .Y(_05541_));
NOT_g _27179_ (.A(_05541_), .Y(_05542_));
NAND_g _27180_ (.A(_11143_), .B(_00012_[2]), .Y(_05543_));
AND_g _27181_ (.A(_00012_[0]), .B(_05543_), .Y(_05544_));
NAND_g _27182_ (.A(_05542_), .B(_05544_), .Y(_05545_));
NOR_g _27183_ (.A(cpuregs_8[6]), .B(_00012_[2]), .Y(_05546_));
NOR_g _27184_ (.A(cpuregs_12[6]), .B(_11214_), .Y(_05547_));
NOR_g _27185_ (.A(_05546_), .B(_05547_), .Y(_05548_));
NAND_g _27186_ (.A(_11212_), .B(_05548_), .Y(_05549_));
NAND_g _27187_ (.A(_05545_), .B(_05549_), .Y(_05550_));
NAND_g _27188_ (.A(_00012_[3]), .B(_05550_), .Y(_05551_));
NAND_g _27189_ (.A(cpuregs_4[6]), .B(_00012_[2]), .Y(_05552_));
NAND_g _27190_ (.A(cpuregs_0[6]), .B(_11214_), .Y(_05553_));
AND_g _27191_ (.A(_05552_), .B(_05553_), .Y(_05554_));
NAND_g _27192_ (.A(_11212_), .B(_05554_), .Y(_05555_));
NAND_g _27193_ (.A(cpuregs_5[6]), .B(_00012_[2]), .Y(_05556_));
NAND_g _27194_ (.A(cpuregs_1[6]), .B(_11214_), .Y(_05557_));
AND_g _27195_ (.A(_00012_[0]), .B(_05557_), .Y(_05558_));
NAND_g _27196_ (.A(_05556_), .B(_05558_), .Y(_05559_));
AND_g _27197_ (.A(_11215_), .B(_05559_), .Y(_05560_));
NAND_g _27198_ (.A(_05555_), .B(_05560_), .Y(_05561_));
NAND_g _27199_ (.A(_05551_), .B(_05561_), .Y(_05562_));
NAND_g _27200_ (.A(_11213_), .B(_05562_), .Y(_05563_));
NAND_g _27201_ (.A(cpuregs_7[6]), .B(_00012_[0]), .Y(_05564_));
NAND_g _27202_ (.A(cpuregs_6[6]), .B(_11212_), .Y(_05565_));
AND_g _27203_ (.A(_00012_[2]), .B(_05565_), .Y(_05566_));
NAND_g _27204_ (.A(_05564_), .B(_05566_), .Y(_05567_));
NAND_g _27205_ (.A(cpuregs_3[6]), .B(_00012_[0]), .Y(_05568_));
NAND_g _27206_ (.A(cpuregs_2[6]), .B(_11212_), .Y(_05569_));
AND_g _27207_ (.A(_11214_), .B(_05569_), .Y(_05570_));
NAND_g _27208_ (.A(_05568_), .B(_05570_), .Y(_05571_));
AND_g _27209_ (.A(_11215_), .B(_05571_), .Y(_05572_));
NAND_g _27210_ (.A(_05567_), .B(_05572_), .Y(_05573_));
NAND_g _27211_ (.A(cpuregs_15[6]), .B(_00012_[0]), .Y(_05574_));
NAND_g _27212_ (.A(cpuregs_14[6]), .B(_11212_), .Y(_05575_));
AND_g _27213_ (.A(_00012_[2]), .B(_05575_), .Y(_05576_));
NAND_g _27214_ (.A(_05574_), .B(_05576_), .Y(_05577_));
NAND_g _27215_ (.A(cpuregs_11[6]), .B(_00012_[0]), .Y(_05578_));
NAND_g _27216_ (.A(cpuregs_10[6]), .B(_11212_), .Y(_05579_));
AND_g _27217_ (.A(_11214_), .B(_05579_), .Y(_05580_));
NAND_g _27218_ (.A(_05578_), .B(_05580_), .Y(_05581_));
AND_g _27219_ (.A(_00012_[3]), .B(_05581_), .Y(_05582_));
NAND_g _27220_ (.A(_05577_), .B(_05582_), .Y(_05583_));
NAND_g _27221_ (.A(_05573_), .B(_05583_), .Y(_05584_));
NAND_g _27222_ (.A(_00012_[1]), .B(_05584_), .Y(_05585_));
AND_g _27223_ (.A(_05563_), .B(_05585_), .Y(_05586_));
NAND_g _27224_ (.A(_11216_), .B(_05586_), .Y(_05587_));
NAND_g _27225_ (.A(_11095_), .B(_00012_[2]), .Y(_05588_));
NOR_g _27226_ (.A(cpuregs_24[6]), .B(_00012_[2]), .Y(_05589_));
NOR_g _27227_ (.A(_00012_[0]), .B(_05589_), .Y(_05590_));
AND_g _27228_ (.A(_05588_), .B(_05590_), .Y(_05591_));
NOR_g _27229_ (.A(cpuregs_25[6]), .B(_00012_[2]), .Y(_05592_));
NAND_g _27230_ (.A(_10925_), .B(_00012_[2]), .Y(_05593_));
NOR_g _27231_ (.A(_11212_), .B(_05592_), .Y(_05594_));
AND_g _27232_ (.A(_05593_), .B(_05594_), .Y(_05595_));
NOR_g _27233_ (.A(_05591_), .B(_05595_), .Y(_05596_));
NAND_g _27234_ (.A(_11194_), .B(_00012_[2]), .Y(_05597_));
NOR_g _27235_ (.A(cpuregs_16[6]), .B(_00012_[2]), .Y(_05598_));
NOR_g _27236_ (.A(_00012_[0]), .B(_05598_), .Y(_05599_));
NAND_g _27237_ (.A(_05597_), .B(_05599_), .Y(_05600_));
NAND_g _27238_ (.A(_11025_), .B(_00012_[2]), .Y(_05601_));
NOR_g _27239_ (.A(cpuregs_17[6]), .B(_00012_[2]), .Y(_05602_));
NOR_g _27240_ (.A(_11212_), .B(_05602_), .Y(_05603_));
NAND_g _27241_ (.A(_05601_), .B(_05603_), .Y(_05604_));
NAND_g _27242_ (.A(_00012_[3]), .B(_05596_), .Y(_05605_));
AND_g _27243_ (.A(_11215_), .B(_05600_), .Y(_05606_));
NAND_g _27244_ (.A(_05604_), .B(_05606_), .Y(_05607_));
AND_g _27245_ (.A(_05605_), .B(_05607_), .Y(_05608_));
NAND_g _27246_ (.A(_11213_), .B(_05608_), .Y(_05609_));
NAND_g _27247_ (.A(cpuregs_23[6]), .B(_11215_), .Y(_05610_));
NAND_g _27248_ (.A(cpuregs_31[6]), .B(_00012_[3]), .Y(_05611_));
AND_g _27249_ (.A(_00012_[2]), .B(_05611_), .Y(_05612_));
NAND_g _27250_ (.A(_05610_), .B(_05612_), .Y(_05613_));
NAND_g _27251_ (.A(cpuregs_19[6]), .B(_11215_), .Y(_05614_));
NAND_g _27252_ (.A(cpuregs_27[6]), .B(_00012_[3]), .Y(_05615_));
AND_g _27253_ (.A(_11214_), .B(_05615_), .Y(_05616_));
NAND_g _27254_ (.A(_05614_), .B(_05616_), .Y(_05617_));
AND_g _27255_ (.A(_00012_[0]), .B(_05617_), .Y(_05618_));
NAND_g _27256_ (.A(_05613_), .B(_05618_), .Y(_05619_));
NAND_g _27257_ (.A(cpuregs_22[6]), .B(_11215_), .Y(_05620_));
NAND_g _27258_ (.A(cpuregs_30[6]), .B(_00012_[3]), .Y(_05621_));
AND_g _27259_ (.A(_00012_[2]), .B(_05621_), .Y(_05622_));
NAND_g _27260_ (.A(_05620_), .B(_05622_), .Y(_05623_));
NAND_g _27261_ (.A(cpuregs_18[6]), .B(_11215_), .Y(_05624_));
NAND_g _27262_ (.A(cpuregs_26[6]), .B(_00012_[3]), .Y(_05625_));
AND_g _27263_ (.A(_11214_), .B(_05625_), .Y(_05626_));
NAND_g _27264_ (.A(_05624_), .B(_05626_), .Y(_05627_));
AND_g _27265_ (.A(_11212_), .B(_05627_), .Y(_05628_));
NAND_g _27266_ (.A(_05623_), .B(_05628_), .Y(_05629_));
NAND_g _27267_ (.A(_05619_), .B(_05629_), .Y(_05630_));
NAND_g _27268_ (.A(_00012_[1]), .B(_05630_), .Y(_05631_));
AND_g _27269_ (.A(_05609_), .B(_05631_), .Y(_05632_));
NAND_g _27270_ (.A(_00012_[4]), .B(_05632_), .Y(_05633_));
AND_g _27271_ (.A(_13409_), .B(_05633_), .Y(_05634_));
AND_g _27272_ (.A(_05587_), .B(_05634_), .Y(_05635_));
AND_g _27273_ (.A(_13613_), .B(_05635_), .Y(_05636_));
NAND_g _27274_ (.A(reg_pc[6]), .B(_13714_), .Y(_05637_));
NAND_g _27275_ (.A(pcpi_rs1[10]), .B(_13419_), .Y(_05638_));
AND_g _27276_ (.A(_13383_), .B(_05638_), .Y(_05639_));
NAND_g _27277_ (.A(_05303_), .B(_05639_), .Y(_05640_));
NAND_g _27278_ (.A(pcpi_rs1[5]), .B(_13420_), .Y(_05641_));
AND_g _27279_ (.A(_13382_), .B(_05641_), .Y(_05642_));
NAND_g _27280_ (.A(_05305_), .B(_05642_), .Y(_05643_));
AND_g _27281_ (.A(_05640_), .B(_05643_), .Y(_05644_));
NAND_g _27282_ (.A(_13389_), .B(_05644_), .Y(_05645_));
NAND_g _27283_ (.A(_05637_), .B(_05645_), .Y(_05646_));
NOR_g _27284_ (.A(_05636_), .B(_05646_), .Y(_05647_));
AND_g _27285_ (.A(_13425_), .B(_05647_), .Y(_05648_));
XOR_g _27286_ (.A(_13481_), .B(_13502_), .Y(_05649_));
NAND_g _27287_ (.A(_13432_), .B(_05649_), .Y(_05650_));
AND_g _27288_ (.A(_05648_), .B(_05650_), .Y(_05651_));
NOR_g _27289_ (.A(pcpi_rs1[6]), .B(_13425_), .Y(_05652_));
NOR_g _27290_ (.A(_05651_), .B(_05652_), .Y(_01213_));
XOR_g _27291_ (.A(decoded_imm[7]), .B(pcpi_rs1[7]), .Y(_05653_));
XNOR_g _27292_ (.A(_13504_), .B(_05653_), .Y(_05654_));
NAND_g _27293_ (.A(_13432_), .B(_05654_), .Y(_05655_));
NAND_g _27294_ (.A(cpuregs_13[7]), .B(_00012_[2]), .Y(_05656_));
NAND_g _27295_ (.A(cpuregs_9[7]), .B(_11214_), .Y(_05657_));
NAND_g _27296_ (.A(_05656_), .B(_05657_), .Y(_05658_));
NAND_g _27297_ (.A(_00012_[0]), .B(_05658_), .Y(_05659_));
NAND_g _27298_ (.A(cpuregs_12[7]), .B(_00012_[2]), .Y(_05660_));
NAND_g _27299_ (.A(cpuregs_8[7]), .B(_11214_), .Y(_05661_));
AND_g _27300_ (.A(_05660_), .B(_05661_), .Y(_05662_));
NOR_g _27301_ (.A(_00012_[0]), .B(_05662_), .Y(_05663_));
NAND_g _27302_ (.A(_10952_), .B(_00012_[2]), .Y(_05664_));
NOR_g _27303_ (.A(cpuregs_0[7]), .B(_00012_[2]), .Y(_05665_));
NOR_g _27304_ (.A(_00012_[0]), .B(_05665_), .Y(_05666_));
NAND_g _27305_ (.A(_05664_), .B(_05666_), .Y(_05667_));
NAND_g _27306_ (.A(_11110_), .B(_00012_[2]), .Y(_05668_));
NOR_g _27307_ (.A(cpuregs_1[7]), .B(_00012_[2]), .Y(_05669_));
NOR_g _27308_ (.A(_11212_), .B(_05669_), .Y(_05670_));
NAND_g _27309_ (.A(_05668_), .B(_05670_), .Y(_05671_));
NAND_g _27310_ (.A(cpuregs_11[7]), .B(_11214_), .Y(_05672_));
NAND_g _27311_ (.A(cpuregs_15[7]), .B(_00012_[2]), .Y(_05673_));
NAND_g _27312_ (.A(_05672_), .B(_05673_), .Y(_05674_));
AND_g _27313_ (.A(_00012_[0]), .B(_05674_), .Y(_05675_));
NAND_g _27314_ (.A(cpuregs_14[7]), .B(_00012_[2]), .Y(_05676_));
NAND_g _27315_ (.A(cpuregs_10[7]), .B(_11214_), .Y(_05677_));
AND_g _27316_ (.A(_05676_), .B(_05677_), .Y(_05678_));
NOR_g _27317_ (.A(_00012_[0]), .B(_05678_), .Y(_05679_));
NOR_g _27318_ (.A(_05675_), .B(_05679_), .Y(_05680_));
NAND_g _27319_ (.A(_10940_), .B(_00012_[2]), .Y(_05681_));
NOR_g _27320_ (.A(cpuregs_2[7]), .B(_00012_[2]), .Y(_05682_));
NOR_g _27321_ (.A(_00012_[0]), .B(_05682_), .Y(_05683_));
NAND_g _27322_ (.A(_05681_), .B(_05683_), .Y(_05684_));
NAND_g _27323_ (.A(_11126_), .B(_00012_[2]), .Y(_05685_));
NOR_g _27324_ (.A(cpuregs_3[7]), .B(_00012_[2]), .Y(_05686_));
NOR_g _27325_ (.A(_11212_), .B(_05686_), .Y(_05687_));
NAND_g _27326_ (.A(_05685_), .B(_05687_), .Y(_05688_));
AND_g _27327_ (.A(_05684_), .B(_05688_), .Y(_05689_));
NAND_g _27328_ (.A(_00012_[1]), .B(_05689_), .Y(_05690_));
AND_g _27329_ (.A(_11213_), .B(_05667_), .Y(_05691_));
NAND_g _27330_ (.A(_05671_), .B(_05691_), .Y(_05692_));
AND_g _27331_ (.A(_05690_), .B(_05692_), .Y(_05693_));
NAND_g _27332_ (.A(_11215_), .B(_05693_), .Y(_05694_));
NAND_g _27333_ (.A(_00012_[1]), .B(_05680_), .Y(_05695_));
NOR_g _27334_ (.A(_00012_[1]), .B(_05663_), .Y(_05696_));
NAND_g _27335_ (.A(_05659_), .B(_05696_), .Y(_05697_));
AND_g _27336_ (.A(_00012_[3]), .B(_05697_), .Y(_05698_));
NAND_g _27337_ (.A(_05695_), .B(_05698_), .Y(_05699_));
AND_g _27338_ (.A(_05694_), .B(_05699_), .Y(_05700_));
NAND_g _27339_ (.A(_11216_), .B(_05700_), .Y(_05701_));
NAND_g _27340_ (.A(cpuregs_20[7]), .B(_11213_), .Y(_05702_));
NAND_g _27341_ (.A(cpuregs_22[7]), .B(_00012_[1]), .Y(_05703_));
AND_g _27342_ (.A(_00012_[2]), .B(_05703_), .Y(_05704_));
NAND_g _27343_ (.A(_05702_), .B(_05704_), .Y(_05705_));
NAND_g _27344_ (.A(cpuregs_16[7]), .B(_11213_), .Y(_05706_));
NAND_g _27345_ (.A(cpuregs_18[7]), .B(_00012_[1]), .Y(_05707_));
AND_g _27346_ (.A(_11214_), .B(_05707_), .Y(_05708_));
NAND_g _27347_ (.A(_05706_), .B(_05708_), .Y(_05709_));
AND_g _27348_ (.A(_11212_), .B(_05709_), .Y(_05710_));
NAND_g _27349_ (.A(_05705_), .B(_05710_), .Y(_05711_));
NAND_g _27350_ (.A(cpuregs_21[7]), .B(_11213_), .Y(_05712_));
NAND_g _27351_ (.A(cpuregs_23[7]), .B(_00012_[1]), .Y(_05713_));
AND_g _27352_ (.A(_00012_[2]), .B(_05713_), .Y(_05714_));
NAND_g _27353_ (.A(_05712_), .B(_05714_), .Y(_05715_));
NAND_g _27354_ (.A(cpuregs_17[7]), .B(_11213_), .Y(_05716_));
NAND_g _27355_ (.A(cpuregs_19[7]), .B(_00012_[1]), .Y(_05717_));
AND_g _27356_ (.A(_11214_), .B(_05717_), .Y(_05718_));
NAND_g _27357_ (.A(_05716_), .B(_05718_), .Y(_05719_));
AND_g _27358_ (.A(_00012_[0]), .B(_05719_), .Y(_05720_));
NAND_g _27359_ (.A(_05715_), .B(_05720_), .Y(_05721_));
NAND_g _27360_ (.A(_05711_), .B(_05721_), .Y(_05722_));
NAND_g _27361_ (.A(_11215_), .B(_05722_), .Y(_05723_));
NAND_g _27362_ (.A(cpuregs_26[7]), .B(_11214_), .Y(_05724_));
NAND_g _27363_ (.A(cpuregs_30[7]), .B(_00012_[2]), .Y(_05725_));
AND_g _27364_ (.A(_00012_[1]), .B(_05725_), .Y(_05726_));
NAND_g _27365_ (.A(_05724_), .B(_05726_), .Y(_05727_));
NAND_g _27366_ (.A(cpuregs_24[7]), .B(_11214_), .Y(_05728_));
NAND_g _27367_ (.A(cpuregs_28[7]), .B(_00012_[2]), .Y(_05729_));
AND_g _27368_ (.A(_11213_), .B(_05729_), .Y(_05730_));
NAND_g _27369_ (.A(_05728_), .B(_05730_), .Y(_05731_));
AND_g _27370_ (.A(_11212_), .B(_05731_), .Y(_05732_));
NAND_g _27371_ (.A(_05727_), .B(_05732_), .Y(_05733_));
NAND_g _27372_ (.A(cpuregs_27[7]), .B(_11214_), .Y(_05734_));
NAND_g _27373_ (.A(cpuregs_31[7]), .B(_00012_[2]), .Y(_05735_));
AND_g _27374_ (.A(_00012_[1]), .B(_05735_), .Y(_05736_));
NAND_g _27375_ (.A(_05734_), .B(_05736_), .Y(_05737_));
NAND_g _27376_ (.A(cpuregs_29[7]), .B(_00012_[2]), .Y(_05738_));
NAND_g _27377_ (.A(cpuregs_25[7]), .B(_11214_), .Y(_05739_));
AND_g _27378_ (.A(_11213_), .B(_05739_), .Y(_05740_));
NAND_g _27379_ (.A(_05738_), .B(_05740_), .Y(_05741_));
AND_g _27380_ (.A(_00012_[0]), .B(_05741_), .Y(_05742_));
NAND_g _27381_ (.A(_05737_), .B(_05742_), .Y(_05743_));
NAND_g _27382_ (.A(_05733_), .B(_05743_), .Y(_05744_));
NAND_g _27383_ (.A(_00012_[3]), .B(_05744_), .Y(_05745_));
AND_g _27384_ (.A(_00012_[4]), .B(_05723_), .Y(_05746_));
NAND_g _27385_ (.A(_05745_), .B(_05746_), .Y(_05747_));
AND_g _27386_ (.A(_13409_), .B(_05747_), .Y(_05748_));
AND_g _27387_ (.A(_05701_), .B(_05748_), .Y(_05749_));
AND_g _27388_ (.A(_13613_), .B(_05749_), .Y(_05750_));
NAND_g _27389_ (.A(reg_pc[7]), .B(_13714_), .Y(_05751_));
NAND_g _27390_ (.A(pcpi_rs1[11]), .B(_13419_), .Y(_05752_));
AND_g _27391_ (.A(_13383_), .B(_05417_), .Y(_05753_));
NAND_g _27392_ (.A(_05752_), .B(_05753_), .Y(_05754_));
NAND_g _27393_ (.A(pcpi_rs1[6]), .B(_13420_), .Y(_05755_));
AND_g _27394_ (.A(_13382_), .B(_05755_), .Y(_05756_));
NAND_g _27395_ (.A(_05420_), .B(_05756_), .Y(_05757_));
AND_g _27396_ (.A(_13389_), .B(_05754_), .Y(_05758_));
AND_g _27397_ (.A(_05757_), .B(_05758_), .Y(_05759_));
NOR_g _27398_ (.A(_05750_), .B(_05759_), .Y(_05760_));
AND_g _27399_ (.A(_13425_), .B(_05760_), .Y(_05761_));
AND_g _27400_ (.A(_05751_), .B(_05761_), .Y(_05762_));
AND_g _27401_ (.A(_05655_), .B(_05762_), .Y(_05763_));
NOR_g _27402_ (.A(pcpi_rs1[7]), .B(_13425_), .Y(_05764_));
NOR_g _27403_ (.A(_05763_), .B(_05764_), .Y(_01214_));
AND_g _27404_ (.A(_13409_), .B(_13612_), .Y(_05765_));
NAND_g _27405_ (.A(_11096_), .B(_00012_[2]), .Y(_05766_));
NOR_g _27406_ (.A(cpuregs_24[8]), .B(_00012_[2]), .Y(_05767_));
NOR_g _27407_ (.A(_00012_[0]), .B(_05767_), .Y(_05768_));
NAND_g _27408_ (.A(_05766_), .B(_05768_), .Y(_05769_));
NAND_g _27409_ (.A(_10926_), .B(_00012_[2]), .Y(_05770_));
NOR_g _27410_ (.A(cpuregs_25[8]), .B(_00012_[2]), .Y(_05771_));
NOR_g _27411_ (.A(_11212_), .B(_05771_), .Y(_05772_));
NAND_g _27412_ (.A(_05770_), .B(_05772_), .Y(_05773_));
NAND_g _27413_ (.A(_05769_), .B(_05773_), .Y(_05774_));
NAND_g _27414_ (.A(_00012_[3]), .B(_05774_), .Y(_05775_));
NAND_g _27415_ (.A(cpuregs_20[8]), .B(_00012_[2]), .Y(_05776_));
NAND_g _27416_ (.A(cpuregs_16[8]), .B(_11214_), .Y(_05777_));
AND_g _27417_ (.A(_05776_), .B(_05777_), .Y(_05778_));
NAND_g _27418_ (.A(_11212_), .B(_05778_), .Y(_05779_));
NAND_g _27419_ (.A(cpuregs_21[8]), .B(_00012_[2]), .Y(_05780_));
NAND_g _27420_ (.A(cpuregs_17[8]), .B(_11214_), .Y(_05781_));
AND_g _27421_ (.A(_00012_[0]), .B(_05781_), .Y(_05782_));
NAND_g _27422_ (.A(_05780_), .B(_05782_), .Y(_05783_));
AND_g _27423_ (.A(_11215_), .B(_05783_), .Y(_05784_));
NAND_g _27424_ (.A(_05779_), .B(_05784_), .Y(_05785_));
AND_g _27425_ (.A(_05775_), .B(_05785_), .Y(_05786_));
NAND_g _27426_ (.A(cpuregs_1[8]), .B(_11214_), .Y(_05787_));
NAND_g _27427_ (.A(cpuregs_5[8]), .B(_00012_[2]), .Y(_05788_));
AND_g _27428_ (.A(_00012_[0]), .B(_05788_), .Y(_05789_));
NAND_g _27429_ (.A(_05787_), .B(_05789_), .Y(_05790_));
NAND_g _27430_ (.A(cpuregs_0[8]), .B(_11214_), .Y(_05791_));
NAND_g _27431_ (.A(cpuregs_4[8]), .B(_00012_[2]), .Y(_05792_));
AND_g _27432_ (.A(_11212_), .B(_05792_), .Y(_05793_));
NAND_g _27433_ (.A(_05791_), .B(_05793_), .Y(_05794_));
AND_g _27434_ (.A(_11215_), .B(_05790_), .Y(_05795_));
NAND_g _27435_ (.A(_05794_), .B(_05795_), .Y(_05796_));
NAND_g _27436_ (.A(cpuregs_9[8]), .B(_11214_), .Y(_05797_));
NAND_g _27437_ (.A(cpuregs_13[8]), .B(_00012_[2]), .Y(_05798_));
AND_g _27438_ (.A(_00012_[0]), .B(_05798_), .Y(_05799_));
NAND_g _27439_ (.A(_05797_), .B(_05799_), .Y(_05800_));
NAND_g _27440_ (.A(cpuregs_8[8]), .B(_11214_), .Y(_05801_));
NAND_g _27441_ (.A(cpuregs_12[8]), .B(_00012_[2]), .Y(_05802_));
AND_g _27442_ (.A(_11212_), .B(_05802_), .Y(_05803_));
NAND_g _27443_ (.A(_05801_), .B(_05803_), .Y(_05804_));
AND_g _27444_ (.A(_00012_[3]), .B(_05804_), .Y(_05805_));
NAND_g _27445_ (.A(_05800_), .B(_05805_), .Y(_05806_));
AND_g _27446_ (.A(_05796_), .B(_05806_), .Y(_05807_));
NAND_g _27447_ (.A(_11173_), .B(_00012_[2]), .Y(_05808_));
NOR_g _27448_ (.A(cpuregs_26[8]), .B(_00012_[2]), .Y(_05809_));
NOR_g _27449_ (.A(_00012_[0]), .B(_05809_), .Y(_05810_));
NAND_g _27450_ (.A(_05808_), .B(_05810_), .Y(_05811_));
NAND_g _27451_ (.A(_11089_), .B(_00012_[2]), .Y(_05812_));
NOR_g _27452_ (.A(cpuregs_27[8]), .B(_00012_[2]), .Y(_05813_));
NOR_g _27453_ (.A(_11212_), .B(_05813_), .Y(_05814_));
NAND_g _27454_ (.A(_05812_), .B(_05814_), .Y(_05815_));
NAND_g _27455_ (.A(_05811_), .B(_05815_), .Y(_05816_));
NAND_g _27456_ (.A(_00012_[3]), .B(_05816_), .Y(_05817_));
NAND_g _27457_ (.A(cpuregs_22[8]), .B(_00012_[2]), .Y(_05818_));
NAND_g _27458_ (.A(cpuregs_18[8]), .B(_11214_), .Y(_05819_));
AND_g _27459_ (.A(_05818_), .B(_05819_), .Y(_05820_));
NAND_g _27460_ (.A(_11212_), .B(_05820_), .Y(_05821_));
NAND_g _27461_ (.A(cpuregs_23[8]), .B(_00012_[2]), .Y(_05822_));
NAND_g _27462_ (.A(cpuregs_19[8]), .B(_11214_), .Y(_05823_));
AND_g _27463_ (.A(_00012_[0]), .B(_05823_), .Y(_05824_));
NAND_g _27464_ (.A(_05822_), .B(_05824_), .Y(_05825_));
AND_g _27465_ (.A(_11215_), .B(_05825_), .Y(_05826_));
NAND_g _27466_ (.A(_05821_), .B(_05826_), .Y(_05827_));
AND_g _27467_ (.A(_05817_), .B(_05827_), .Y(_05828_));
NAND_g _27468_ (.A(_00012_[1]), .B(_05828_), .Y(_05829_));
NAND_g _27469_ (.A(_11213_), .B(_05786_), .Y(_05830_));
AND_g _27470_ (.A(_00012_[4]), .B(_05830_), .Y(_05831_));
NAND_g _27471_ (.A(_05829_), .B(_05831_), .Y(_05832_));
NAND_g _27472_ (.A(_11213_), .B(_05807_), .Y(_05833_));
NAND_g _27473_ (.A(cpuregs_6[8]), .B(_00012_[2]), .Y(_05834_));
NAND_g _27474_ (.A(cpuregs_2[8]), .B(_11214_), .Y(_05835_));
AND_g _27475_ (.A(_05834_), .B(_05835_), .Y(_05836_));
NAND_g _27476_ (.A(_11212_), .B(_05836_), .Y(_05837_));
NAND_g _27477_ (.A(cpuregs_7[8]), .B(_00012_[2]), .Y(_05838_));
NAND_g _27478_ (.A(cpuregs_3[8]), .B(_11214_), .Y(_05839_));
AND_g _27479_ (.A(_00012_[0]), .B(_05839_), .Y(_05840_));
NAND_g _27480_ (.A(_05838_), .B(_05840_), .Y(_05841_));
AND_g _27481_ (.A(_11215_), .B(_05841_), .Y(_05842_));
NAND_g _27482_ (.A(_05837_), .B(_05842_), .Y(_05843_));
NOR_g _27483_ (.A(cpuregs_11[8]), .B(_00012_[2]), .Y(_05844_));
NOT_g _27484_ (.A(_05844_), .Y(_05845_));
NAND_g _27485_ (.A(_11159_), .B(_00012_[2]), .Y(_05846_));
AND_g _27486_ (.A(_00012_[0]), .B(_05846_), .Y(_05847_));
NAND_g _27487_ (.A(_05845_), .B(_05847_), .Y(_05848_));
NOR_g _27488_ (.A(cpuregs_10[8]), .B(_00012_[2]), .Y(_05849_));
AND_g _27489_ (.A(_11102_), .B(_00012_[2]), .Y(_05850_));
NOR_g _27490_ (.A(_05849_), .B(_05850_), .Y(_05851_));
NAND_g _27491_ (.A(_11212_), .B(_05851_), .Y(_05852_));
NAND_g _27492_ (.A(_05848_), .B(_05852_), .Y(_05853_));
NAND_g _27493_ (.A(_00012_[3]), .B(_05853_), .Y(_05854_));
AND_g _27494_ (.A(_05843_), .B(_05854_), .Y(_05855_));
NAND_g _27495_ (.A(_00012_[1]), .B(_05855_), .Y(_05856_));
AND_g _27496_ (.A(_05833_), .B(_05856_), .Y(_05857_));
NAND_g _27497_ (.A(_11216_), .B(_05857_), .Y(_05858_));
NAND_g _27498_ (.A(_05832_), .B(_05858_), .Y(_05859_));
AND_g _27499_ (.A(_13561_), .B(_05859_), .Y(_05860_));
NAND_g _27500_ (.A(_05765_), .B(_05860_), .Y(_05861_));
NAND_g _27501_ (.A(reg_pc[8]), .B(_13714_), .Y(_05862_));
NAND_g _27502_ (.A(pcpi_rs1[7]), .B(_13420_), .Y(_05863_));
AND_g _27503_ (.A(_05529_), .B(_05863_), .Y(_05864_));
NAND_g _27504_ (.A(_13382_), .B(_05864_), .Y(_05865_));
NAND_g _27505_ (.A(pcpi_rs1[12]), .B(_13419_), .Y(_05866_));
AND_g _27506_ (.A(_05528_), .B(_05866_), .Y(_05867_));
NAND_g _27507_ (.A(_13383_), .B(_05867_), .Y(_05868_));
AND_g _27508_ (.A(_05865_), .B(_05868_), .Y(_05869_));
NAND_g _27509_ (.A(_13389_), .B(_05869_), .Y(_05870_));
AND_g _27510_ (.A(_05862_), .B(_05870_), .Y(_05871_));
AND_g _27511_ (.A(_05861_), .B(_05871_), .Y(_05872_));
XOR_g _27512_ (.A(_13477_), .B(_13506_), .Y(_05873_));
NAND_g _27513_ (.A(_13432_), .B(_05873_), .Y(_05874_));
AND_g _27514_ (.A(_05872_), .B(_05874_), .Y(_05875_));
NOR_g _27515_ (.A(pcpi_rs1[8]), .B(_13425_), .Y(_05876_));
AND_g _27516_ (.A(_13425_), .B(_05875_), .Y(_05877_));
NOR_g _27517_ (.A(_05876_), .B(_05877_), .Y(_01215_));
NOR_g _27518_ (.A(pcpi_rs1[9]), .B(_13425_), .Y(_05878_));
XOR_g _27519_ (.A(decoded_imm[9]), .B(pcpi_rs1[9]), .Y(_05879_));
XNOR_g _27520_ (.A(_13508_), .B(_05879_), .Y(_05880_));
NAND_g _27521_ (.A(_13432_), .B(_05880_), .Y(_05881_));
NAND_g _27522_ (.A(cpuregs_7[9]), .B(_00012_[2]), .Y(_05882_));
NAND_g _27523_ (.A(cpuregs_3[9]), .B(_11214_), .Y(_05883_));
NAND_g _27524_ (.A(_05882_), .B(_05883_), .Y(_05884_));
AND_g _27525_ (.A(_00012_[0]), .B(_05884_), .Y(_05885_));
NAND_g _27526_ (.A(cpuregs_6[9]), .B(_00012_[2]), .Y(_05886_));
NAND_g _27527_ (.A(cpuregs_2[9]), .B(_11214_), .Y(_05887_));
AND_g _27528_ (.A(_05886_), .B(_05887_), .Y(_05888_));
NOR_g _27529_ (.A(_00012_[0]), .B(_05888_), .Y(_05889_));
NOR_g _27530_ (.A(_05885_), .B(_05889_), .Y(_05890_));
NAND_g _27531_ (.A(cpuregs_5[9]), .B(_00012_[2]), .Y(_05891_));
NAND_g _27532_ (.A(cpuregs_1[9]), .B(_11214_), .Y(_05892_));
NAND_g _27533_ (.A(_05891_), .B(_05892_), .Y(_05893_));
NAND_g _27534_ (.A(_00012_[0]), .B(_05893_), .Y(_05894_));
NAND_g _27535_ (.A(cpuregs_4[9]), .B(_00012_[2]), .Y(_05895_));
NAND_g _27536_ (.A(cpuregs_0[9]), .B(_11214_), .Y(_05896_));
AND_g _27537_ (.A(_05895_), .B(_05896_), .Y(_05897_));
NOR_g _27538_ (.A(_00012_[0]), .B(_05897_), .Y(_05898_));
NAND_g _27539_ (.A(_00012_[1]), .B(_05890_), .Y(_05899_));
NOR_g _27540_ (.A(_00012_[1]), .B(_05898_), .Y(_05900_));
NAND_g _27541_ (.A(_05894_), .B(_05900_), .Y(_05901_));
AND_g _27542_ (.A(_05899_), .B(_05901_), .Y(_05902_));
NAND_g _27543_ (.A(_11215_), .B(_05902_), .Y(_05903_));
NAND_g _27544_ (.A(cpuregs_13[9]), .B(_00012_[0]), .Y(_05904_));
NAND_g _27545_ (.A(cpuregs_12[9]), .B(_11212_), .Y(_05905_));
AND_g _27546_ (.A(_00012_[2]), .B(_05905_), .Y(_05906_));
NAND_g _27547_ (.A(_05904_), .B(_05906_), .Y(_05907_));
NAND_g _27548_ (.A(cpuregs_9[9]), .B(_00012_[0]), .Y(_05908_));
NAND_g _27549_ (.A(cpuregs_8[9]), .B(_11212_), .Y(_05909_));
AND_g _27550_ (.A(_11214_), .B(_05909_), .Y(_05910_));
NAND_g _27551_ (.A(_05908_), .B(_05910_), .Y(_05911_));
AND_g _27552_ (.A(_11213_), .B(_05911_), .Y(_05912_));
NAND_g _27553_ (.A(_05907_), .B(_05912_), .Y(_05913_));
NAND_g _27554_ (.A(cpuregs_15[9]), .B(_00012_[0]), .Y(_05914_));
NAND_g _27555_ (.A(cpuregs_14[9]), .B(_11212_), .Y(_05915_));
AND_g _27556_ (.A(_00012_[2]), .B(_05915_), .Y(_05916_));
NAND_g _27557_ (.A(_05914_), .B(_05916_), .Y(_05917_));
NAND_g _27558_ (.A(cpuregs_11[9]), .B(_00012_[0]), .Y(_05918_));
NAND_g _27559_ (.A(cpuregs_10[9]), .B(_11212_), .Y(_05919_));
AND_g _27560_ (.A(_11214_), .B(_05919_), .Y(_05920_));
NAND_g _27561_ (.A(_05918_), .B(_05920_), .Y(_05921_));
AND_g _27562_ (.A(_00012_[1]), .B(_05921_), .Y(_05922_));
NAND_g _27563_ (.A(_05917_), .B(_05922_), .Y(_05923_));
NAND_g _27564_ (.A(_05913_), .B(_05923_), .Y(_05924_));
NAND_g _27565_ (.A(_00012_[3]), .B(_05924_), .Y(_05925_));
AND_g _27566_ (.A(_05903_), .B(_05925_), .Y(_05926_));
NAND_g _27567_ (.A(_11216_), .B(_05926_), .Y(_05927_));
NAND_g _27568_ (.A(cpuregs_31[9]), .B(_00012_[2]), .Y(_05928_));
NAND_g _27569_ (.A(cpuregs_27[9]), .B(_11214_), .Y(_05929_));
NAND_g _27570_ (.A(_05928_), .B(_05929_), .Y(_05930_));
AND_g _27571_ (.A(_00012_[0]), .B(_05930_), .Y(_05931_));
NAND_g _27572_ (.A(cpuregs_30[9]), .B(_00012_[2]), .Y(_05932_));
NAND_g _27573_ (.A(cpuregs_26[9]), .B(_11214_), .Y(_05933_));
AND_g _27574_ (.A(_05932_), .B(_05933_), .Y(_05934_));
NOR_g _27575_ (.A(_00012_[0]), .B(_05934_), .Y(_05935_));
NOR_g _27576_ (.A(_05931_), .B(_05935_), .Y(_05936_));
NAND_g _27577_ (.A(cpuregs_25[9]), .B(_11214_), .Y(_05937_));
NAND_g _27578_ (.A(cpuregs_29[9]), .B(_00012_[2]), .Y(_05938_));
NAND_g _27579_ (.A(_05937_), .B(_05938_), .Y(_05939_));
NAND_g _27580_ (.A(_00012_[0]), .B(_05939_), .Y(_05940_));
NAND_g _27581_ (.A(cpuregs_28[9]), .B(_00012_[2]), .Y(_05941_));
NAND_g _27582_ (.A(cpuregs_24[9]), .B(_11214_), .Y(_05942_));
NAND_g _27583_ (.A(_05941_), .B(_05942_), .Y(_05943_));
NAND_g _27584_ (.A(_11212_), .B(_05943_), .Y(_05944_));
AND_g _27585_ (.A(_05940_), .B(_05944_), .Y(_05945_));
NAND_g _27586_ (.A(_11213_), .B(_05945_), .Y(_05946_));
NAND_g _27587_ (.A(_00012_[1]), .B(_05936_), .Y(_05947_));
AND_g _27588_ (.A(_00012_[3]), .B(_05947_), .Y(_05948_));
NAND_g _27589_ (.A(_05946_), .B(_05948_), .Y(_05949_));
NAND_g _27590_ (.A(cpuregs_20[9]), .B(_11212_), .Y(_05950_));
NAND_g _27591_ (.A(cpuregs_21[9]), .B(_00012_[0]), .Y(_05951_));
AND_g _27592_ (.A(_00012_[2]), .B(_05951_), .Y(_05952_));
NAND_g _27593_ (.A(_05950_), .B(_05952_), .Y(_05953_));
NAND_g _27594_ (.A(cpuregs_16[9]), .B(_11212_), .Y(_05954_));
NAND_g _27595_ (.A(cpuregs_17[9]), .B(_00012_[0]), .Y(_05955_));
AND_g _27596_ (.A(_11214_), .B(_05955_), .Y(_05956_));
NAND_g _27597_ (.A(_05954_), .B(_05956_), .Y(_05957_));
AND_g _27598_ (.A(_11213_), .B(_05957_), .Y(_05958_));
NAND_g _27599_ (.A(_05953_), .B(_05958_), .Y(_05959_));
NAND_g _27600_ (.A(cpuregs_22[9]), .B(_00012_[2]), .Y(_05960_));
NAND_g _27601_ (.A(cpuregs_18[9]), .B(_11214_), .Y(_05961_));
AND_g _27602_ (.A(_11212_), .B(_05961_), .Y(_05962_));
NAND_g _27603_ (.A(_05960_), .B(_05962_), .Y(_05963_));
NAND_g _27604_ (.A(cpuregs_19[9]), .B(_11214_), .Y(_05964_));
NAND_g _27605_ (.A(cpuregs_23[9]), .B(_00012_[2]), .Y(_05965_));
AND_g _27606_ (.A(_00012_[0]), .B(_05965_), .Y(_05966_));
NAND_g _27607_ (.A(_05964_), .B(_05966_), .Y(_05967_));
AND_g _27608_ (.A(_00012_[1]), .B(_05967_), .Y(_05968_));
NAND_g _27609_ (.A(_05963_), .B(_05968_), .Y(_05969_));
NAND_g _27610_ (.A(_05959_), .B(_05969_), .Y(_05970_));
NAND_g _27611_ (.A(_11215_), .B(_05970_), .Y(_05971_));
AND_g _27612_ (.A(_00012_[4]), .B(_05971_), .Y(_05972_));
NAND_g _27613_ (.A(_05949_), .B(_05972_), .Y(_05973_));
AND_g _27614_ (.A(_05927_), .B(_05973_), .Y(_05974_));
AND_g _27615_ (.A(_13409_), .B(_05974_), .Y(_05975_));
AND_g _27616_ (.A(_13613_), .B(_05975_), .Y(_05976_));
NAND_g _27617_ (.A(reg_pc[9]), .B(_13714_), .Y(_05977_));
NAND_g _27618_ (.A(pcpi_rs1[8]), .B(_13420_), .Y(_05978_));
AND_g _27619_ (.A(_13382_), .B(_05978_), .Y(_05979_));
NAND_g _27620_ (.A(_05638_), .B(_05979_), .Y(_05980_));
NAND_g _27621_ (.A(pcpi_rs1[13]), .B(_13419_), .Y(_05981_));
AND_g _27622_ (.A(_13383_), .B(_05641_), .Y(_05982_));
NAND_g _27623_ (.A(_05981_), .B(_05982_), .Y(_05983_));
AND_g _27624_ (.A(_05980_), .B(_05983_), .Y(_05984_));
NAND_g _27625_ (.A(_13389_), .B(_05984_), .Y(_05985_));
AND_g _27626_ (.A(_05977_), .B(_05985_), .Y(_05986_));
NAND_g _27627_ (.A(_13425_), .B(_05986_), .Y(_05987_));
NOR_g _27628_ (.A(_05976_), .B(_05987_), .Y(_05988_));
AND_g _27629_ (.A(_05881_), .B(_05988_), .Y(_05989_));
NOR_g _27630_ (.A(_05878_), .B(_05989_), .Y(_01216_));
NOR_g _27631_ (.A(pcpi_rs1[10]), .B(_13425_), .Y(_05990_));
XOR_g _27632_ (.A(_13473_), .B(_13510_), .Y(_05991_));
NAND_g _27633_ (.A(_13432_), .B(_05991_), .Y(_05992_));
NAND_g _27634_ (.A(reg_pc[10]), .B(_13714_), .Y(_05993_));
NAND_g _27635_ (.A(pcpi_rs1[9]), .B(_13420_), .Y(_05994_));
AND_g _27636_ (.A(_05752_), .B(_05994_), .Y(_05995_));
NAND_g _27637_ (.A(_13382_), .B(_05995_), .Y(_05996_));
NAND_g _27638_ (.A(pcpi_rs1[14]), .B(_13419_), .Y(_05997_));
AND_g _27639_ (.A(_05755_), .B(_05997_), .Y(_05998_));
NAND_g _27640_ (.A(_13383_), .B(_05998_), .Y(_05999_));
AND_g _27641_ (.A(_05996_), .B(_05999_), .Y(_06000_));
NAND_g _27642_ (.A(_13389_), .B(_06000_), .Y(_06001_));
AND_g _27643_ (.A(_05993_), .B(_06001_), .Y(_06002_));
AND_g _27644_ (.A(_13425_), .B(_06002_), .Y(_06003_));
NOR_g _27645_ (.A(cpuregs_16[10]), .B(_00012_[2]), .Y(_06004_));
AND_g _27646_ (.A(_11195_), .B(_00012_[2]), .Y(_06005_));
NOR_g _27647_ (.A(_06004_), .B(_06005_), .Y(_06006_));
NOR_g _27648_ (.A(cpuregs_18[10]), .B(_00012_[2]), .Y(_06007_));
AND_g _27649_ (.A(_11015_), .B(_00012_[2]), .Y(_06008_));
NOR_g _27650_ (.A(_06007_), .B(_06008_), .Y(_06009_));
NOR_g _27651_ (.A(cpuregs_17[10]), .B(_00012_[2]), .Y(_06010_));
NAND_g _27652_ (.A(_11026_), .B(_00012_[2]), .Y(_06011_));
NAND_g _27653_ (.A(_11180_), .B(_00012_[2]), .Y(_06012_));
NOR_g _27654_ (.A(cpuregs_19[10]), .B(_00012_[2]), .Y(_06013_));
NOR_g _27655_ (.A(_11212_), .B(_06013_), .Y(_06014_));
NAND_g _27656_ (.A(_06012_), .B(_06014_), .Y(_06015_));
NAND_g _27657_ (.A(_11212_), .B(_06009_), .Y(_06016_));
AND_g _27658_ (.A(_06015_), .B(_06016_), .Y(_06017_));
NAND_g _27659_ (.A(_00012_[1]), .B(_06017_), .Y(_06018_));
NOR_g _27660_ (.A(_11212_), .B(_06010_), .Y(_06019_));
NAND_g _27661_ (.A(_06011_), .B(_06019_), .Y(_06020_));
NAND_g _27662_ (.A(_11212_), .B(_06006_), .Y(_06021_));
AND_g _27663_ (.A(_06020_), .B(_06021_), .Y(_06022_));
NAND_g _27664_ (.A(_11213_), .B(_06022_), .Y(_06023_));
AND_g _27665_ (.A(_06018_), .B(_06023_), .Y(_06024_));
NAND_g _27666_ (.A(_11215_), .B(_06024_), .Y(_06025_));
NAND_g _27667_ (.A(cpuregs_27[10]), .B(_00012_[1]), .Y(_06026_));
NAND_g _27668_ (.A(cpuregs_25[10]), .B(_11213_), .Y(_06027_));
NAND_g _27669_ (.A(_06026_), .B(_06027_), .Y(_06028_));
NAND_g _27670_ (.A(_11214_), .B(_06028_), .Y(_06029_));
NAND_g _27671_ (.A(cpuregs_31[10]), .B(_00012_[1]), .Y(_06030_));
NAND_g _27672_ (.A(cpuregs_29[10]), .B(_11213_), .Y(_06031_));
NAND_g _27673_ (.A(_06030_), .B(_06031_), .Y(_06032_));
NAND_g _27674_ (.A(_00012_[2]), .B(_06032_), .Y(_06033_));
AND_g _27675_ (.A(_00012_[0]), .B(_06033_), .Y(_06034_));
NAND_g _27676_ (.A(_06029_), .B(_06034_), .Y(_06035_));
NAND_g _27677_ (.A(cpuregs_26[10]), .B(_00012_[1]), .Y(_06036_));
NAND_g _27678_ (.A(cpuregs_24[10]), .B(_11213_), .Y(_06037_));
NAND_g _27679_ (.A(_06036_), .B(_06037_), .Y(_06038_));
NAND_g _27680_ (.A(_11214_), .B(_06038_), .Y(_06039_));
NAND_g _27681_ (.A(cpuregs_30[10]), .B(_00012_[1]), .Y(_06040_));
NAND_g _27682_ (.A(cpuregs_28[10]), .B(_11213_), .Y(_06041_));
NAND_g _27683_ (.A(_06040_), .B(_06041_), .Y(_06042_));
NAND_g _27684_ (.A(_00012_[2]), .B(_06042_), .Y(_06043_));
AND_g _27685_ (.A(_11212_), .B(_06043_), .Y(_06044_));
NAND_g _27686_ (.A(_06039_), .B(_06044_), .Y(_06045_));
AND_g _27687_ (.A(_00012_[3]), .B(_06045_), .Y(_06046_));
NAND_g _27688_ (.A(_06035_), .B(_06046_), .Y(_06047_));
AND_g _27689_ (.A(_06025_), .B(_06047_), .Y(_06048_));
NAND_g _27690_ (.A(cpuregs_1[10]), .B(_11214_), .Y(_06049_));
NAND_g _27691_ (.A(cpuregs_5[10]), .B(_00012_[2]), .Y(_06050_));
AND_g _27692_ (.A(_00012_[0]), .B(_06050_), .Y(_06051_));
NAND_g _27693_ (.A(_06049_), .B(_06051_), .Y(_06052_));
NAND_g _27694_ (.A(cpuregs_0[10]), .B(_11214_), .Y(_06053_));
NAND_g _27695_ (.A(cpuregs_4[10]), .B(_00012_[2]), .Y(_06054_));
AND_g _27696_ (.A(_11212_), .B(_06054_), .Y(_06055_));
NAND_g _27697_ (.A(_06053_), .B(_06055_), .Y(_06056_));
AND_g _27698_ (.A(_11213_), .B(_06056_), .Y(_06057_));
NAND_g _27699_ (.A(_06052_), .B(_06057_), .Y(_06058_));
NAND_g _27700_ (.A(cpuregs_3[10]), .B(_11214_), .Y(_06059_));
NAND_g _27701_ (.A(cpuregs_7[10]), .B(_00012_[2]), .Y(_06060_));
AND_g _27702_ (.A(_00012_[0]), .B(_06060_), .Y(_06061_));
NAND_g _27703_ (.A(_06059_), .B(_06061_), .Y(_06062_));
NAND_g _27704_ (.A(cpuregs_2[10]), .B(_11214_), .Y(_06063_));
NAND_g _27705_ (.A(cpuregs_6[10]), .B(_00012_[2]), .Y(_06064_));
AND_g _27706_ (.A(_11212_), .B(_06064_), .Y(_06065_));
NAND_g _27707_ (.A(_06063_), .B(_06065_), .Y(_06066_));
AND_g _27708_ (.A(_00012_[1]), .B(_06066_), .Y(_06067_));
NAND_g _27709_ (.A(_06062_), .B(_06067_), .Y(_06068_));
NAND_g _27710_ (.A(_06058_), .B(_06068_), .Y(_06069_));
NAND_g _27711_ (.A(_11215_), .B(_06069_), .Y(_06070_));
NAND_g _27712_ (.A(cpuregs_14[10]), .B(_11212_), .Y(_06071_));
NAND_g _27713_ (.A(cpuregs_15[10]), .B(_00012_[0]), .Y(_06072_));
NAND_g _27714_ (.A(_06071_), .B(_06072_), .Y(_06073_));
NAND_g _27715_ (.A(_00012_[2]), .B(_06073_), .Y(_06074_));
NAND_g _27716_ (.A(cpuregs_10[10]), .B(_11212_), .Y(_06075_));
NAND_g _27717_ (.A(cpuregs_11[10]), .B(_00012_[0]), .Y(_06076_));
NAND_g _27718_ (.A(_06075_), .B(_06076_), .Y(_06077_));
NAND_g _27719_ (.A(_11214_), .B(_06077_), .Y(_06078_));
AND_g _27720_ (.A(_06074_), .B(_06078_), .Y(_06079_));
NAND_g _27721_ (.A(cpuregs_12[10]), .B(_11212_), .Y(_06080_));
NAND_g _27722_ (.A(cpuregs_13[10]), .B(_00012_[0]), .Y(_06081_));
NAND_g _27723_ (.A(_06080_), .B(_06081_), .Y(_06082_));
NAND_g _27724_ (.A(_00012_[2]), .B(_06082_), .Y(_06083_));
NAND_g _27725_ (.A(cpuregs_8[10]), .B(_11212_), .Y(_06084_));
NAND_g _27726_ (.A(cpuregs_9[10]), .B(_00012_[0]), .Y(_06085_));
NAND_g _27727_ (.A(_06084_), .B(_06085_), .Y(_06086_));
NAND_g _27728_ (.A(_11214_), .B(_06086_), .Y(_06087_));
AND_g _27729_ (.A(_06083_), .B(_06087_), .Y(_06088_));
NAND_g _27730_ (.A(_11213_), .B(_06088_), .Y(_06089_));
NAND_g _27731_ (.A(_00012_[1]), .B(_06079_), .Y(_06090_));
AND_g _27732_ (.A(_00012_[3]), .B(_06089_), .Y(_06091_));
NAND_g _27733_ (.A(_06090_), .B(_06091_), .Y(_06092_));
NAND_g _27734_ (.A(_00012_[4]), .B(_06048_), .Y(_06093_));
AND_g _27735_ (.A(_11216_), .B(_06070_), .Y(_06094_));
NAND_g _27736_ (.A(_06092_), .B(_06094_), .Y(_06095_));
AND_g _27737_ (.A(_13561_), .B(_06095_), .Y(_06096_));
AND_g _27738_ (.A(_06093_), .B(_06096_), .Y(_06097_));
NAND_g _27739_ (.A(_05765_), .B(_06097_), .Y(_06098_));
AND_g _27740_ (.A(_06003_), .B(_06098_), .Y(_06099_));
AND_g _27741_ (.A(_05992_), .B(_06099_), .Y(_06100_));
NOR_g _27742_ (.A(_05990_), .B(_06100_), .Y(_01217_));
NOR_g _27743_ (.A(pcpi_rs1[11]), .B(_13425_), .Y(_06101_));
XNOR_g _27744_ (.A(decoded_imm[11]), .B(pcpi_rs1[11]), .Y(_06102_));
NOR_g _27745_ (.A(_13512_), .B(_06102_), .Y(_06103_));
NAND_g _27746_ (.A(_13512_), .B(_06102_), .Y(_06104_));
NAND_g _27747_ (.A(_13432_), .B(_06104_), .Y(_06105_));
NOR_g _27748_ (.A(_06103_), .B(_06105_), .Y(_06106_));
NAND_g _27749_ (.A(cpuregs_13[11]), .B(_00012_[2]), .Y(_06107_));
NAND_g _27750_ (.A(cpuregs_9[11]), .B(_11214_), .Y(_06108_));
NAND_g _27751_ (.A(_06107_), .B(_06108_), .Y(_06109_));
NAND_g _27752_ (.A(_00012_[0]), .B(_06109_), .Y(_06110_));
NAND_g _27753_ (.A(cpuregs_12[11]), .B(_00012_[2]), .Y(_06111_));
NAND_g _27754_ (.A(cpuregs_8[11]), .B(_11214_), .Y(_06112_));
AND_g _27755_ (.A(_06111_), .B(_06112_), .Y(_06113_));
NOR_g _27756_ (.A(_00012_[0]), .B(_06113_), .Y(_06114_));
NAND_g _27757_ (.A(_10954_), .B(_00012_[2]), .Y(_06115_));
NOR_g _27758_ (.A(cpuregs_0[11]), .B(_00012_[2]), .Y(_06116_));
NOR_g _27759_ (.A(_00012_[0]), .B(_06116_), .Y(_06117_));
NAND_g _27760_ (.A(_06115_), .B(_06117_), .Y(_06118_));
NAND_g _27761_ (.A(_11112_), .B(_00012_[2]), .Y(_06119_));
NOR_g _27762_ (.A(cpuregs_1[11]), .B(_00012_[2]), .Y(_06120_));
NOR_g _27763_ (.A(_11212_), .B(_06120_), .Y(_06121_));
NAND_g _27764_ (.A(_06119_), .B(_06121_), .Y(_06122_));
NAND_g _27765_ (.A(cpuregs_11[11]), .B(_11214_), .Y(_06123_));
NAND_g _27766_ (.A(cpuregs_15[11]), .B(_00012_[2]), .Y(_06124_));
NAND_g _27767_ (.A(_06123_), .B(_06124_), .Y(_06125_));
AND_g _27768_ (.A(_00012_[0]), .B(_06125_), .Y(_06126_));
NAND_g _27769_ (.A(cpuregs_14[11]), .B(_00012_[2]), .Y(_06127_));
NAND_g _27770_ (.A(cpuregs_10[11]), .B(_11214_), .Y(_06128_));
AND_g _27771_ (.A(_06127_), .B(_06128_), .Y(_06129_));
NOR_g _27772_ (.A(_00012_[0]), .B(_06129_), .Y(_06130_));
NOR_g _27773_ (.A(_06126_), .B(_06130_), .Y(_06131_));
NAND_g _27774_ (.A(_10942_), .B(_00012_[2]), .Y(_06132_));
NOR_g _27775_ (.A(cpuregs_2[11]), .B(_00012_[2]), .Y(_06133_));
NOR_g _27776_ (.A(_00012_[0]), .B(_06133_), .Y(_06134_));
NAND_g _27777_ (.A(_06132_), .B(_06134_), .Y(_06135_));
NAND_g _27778_ (.A(_11128_), .B(_00012_[2]), .Y(_06136_));
NOR_g _27779_ (.A(cpuregs_3[11]), .B(_00012_[2]), .Y(_06137_));
NOR_g _27780_ (.A(_11212_), .B(_06137_), .Y(_06138_));
NAND_g _27781_ (.A(_06136_), .B(_06138_), .Y(_06139_));
AND_g _27782_ (.A(_06135_), .B(_06139_), .Y(_06140_));
NAND_g _27783_ (.A(_00012_[1]), .B(_06140_), .Y(_06141_));
AND_g _27784_ (.A(_11213_), .B(_06118_), .Y(_06142_));
NAND_g _27785_ (.A(_06122_), .B(_06142_), .Y(_06143_));
AND_g _27786_ (.A(_06141_), .B(_06143_), .Y(_06144_));
NAND_g _27787_ (.A(_11215_), .B(_06144_), .Y(_06145_));
NAND_g _27788_ (.A(_00012_[1]), .B(_06131_), .Y(_06146_));
NOR_g _27789_ (.A(_00012_[1]), .B(_06114_), .Y(_06147_));
NAND_g _27790_ (.A(_06110_), .B(_06147_), .Y(_06148_));
AND_g _27791_ (.A(_00012_[3]), .B(_06148_), .Y(_06149_));
NAND_g _27792_ (.A(_06146_), .B(_06149_), .Y(_06150_));
AND_g _27793_ (.A(_06145_), .B(_06150_), .Y(_06151_));
NAND_g _27794_ (.A(_11216_), .B(_06151_), .Y(_06152_));
NAND_g _27795_ (.A(_11016_), .B(_00012_[2]), .Y(_06153_));
NOR_g _27796_ (.A(cpuregs_18[11]), .B(_00012_[2]), .Y(_06154_));
NOR_g _27797_ (.A(_00012_[0]), .B(_06154_), .Y(_06155_));
NAND_g _27798_ (.A(_06153_), .B(_06155_), .Y(_06156_));
NAND_g _27799_ (.A(_11181_), .B(_00012_[2]), .Y(_06157_));
NOR_g _27800_ (.A(cpuregs_19[11]), .B(_00012_[2]), .Y(_06158_));
NOR_g _27801_ (.A(_11212_), .B(_06158_), .Y(_06159_));
NAND_g _27802_ (.A(_06157_), .B(_06159_), .Y(_06160_));
AND_g _27803_ (.A(_06156_), .B(_06160_), .Y(_06161_));
NAND_g _27804_ (.A(_11196_), .B(_00012_[2]), .Y(_06162_));
NOR_g _27805_ (.A(cpuregs_16[11]), .B(_00012_[2]), .Y(_06163_));
NOR_g _27806_ (.A(_00012_[0]), .B(_06163_), .Y(_06164_));
NAND_g _27807_ (.A(_06162_), .B(_06164_), .Y(_06165_));
NAND_g _27808_ (.A(_11027_), .B(_00012_[2]), .Y(_06166_));
NOR_g _27809_ (.A(cpuregs_17[11]), .B(_00012_[2]), .Y(_06167_));
NOR_g _27810_ (.A(_11212_), .B(_06167_), .Y(_06168_));
NAND_g _27811_ (.A(_06166_), .B(_06168_), .Y(_06169_));
AND_g _27812_ (.A(_06165_), .B(_06169_), .Y(_06170_));
NAND_g _27813_ (.A(_00012_[1]), .B(_06161_), .Y(_06171_));
NAND_g _27814_ (.A(_11213_), .B(_06170_), .Y(_06172_));
AND_g _27815_ (.A(_06171_), .B(_06172_), .Y(_06173_));
NAND_g _27816_ (.A(_11215_), .B(_06173_), .Y(_06174_));
NAND_g _27817_ (.A(cpuregs_29[11]), .B(_11213_), .Y(_06175_));
NAND_g _27818_ (.A(cpuregs_31[11]), .B(_00012_[1]), .Y(_06176_));
AND_g _27819_ (.A(_00012_[2]), .B(_06176_), .Y(_06177_));
NAND_g _27820_ (.A(_06175_), .B(_06177_), .Y(_06178_));
NAND_g _27821_ (.A(cpuregs_25[11]), .B(_11213_), .Y(_06179_));
NAND_g _27822_ (.A(cpuregs_27[11]), .B(_00012_[1]), .Y(_06180_));
AND_g _27823_ (.A(_11214_), .B(_06180_), .Y(_06181_));
NAND_g _27824_ (.A(_06179_), .B(_06181_), .Y(_06182_));
AND_g _27825_ (.A(_00012_[0]), .B(_06182_), .Y(_06183_));
NAND_g _27826_ (.A(_06178_), .B(_06183_), .Y(_06184_));
NAND_g _27827_ (.A(cpuregs_28[11]), .B(_11213_), .Y(_06185_));
NAND_g _27828_ (.A(cpuregs_30[11]), .B(_00012_[1]), .Y(_06186_));
AND_g _27829_ (.A(_00012_[2]), .B(_06186_), .Y(_06187_));
NAND_g _27830_ (.A(_06185_), .B(_06187_), .Y(_06188_));
NAND_g _27831_ (.A(cpuregs_24[11]), .B(_11213_), .Y(_06189_));
NAND_g _27832_ (.A(cpuregs_26[11]), .B(_00012_[1]), .Y(_06190_));
AND_g _27833_ (.A(_11214_), .B(_06190_), .Y(_06191_));
NAND_g _27834_ (.A(_06189_), .B(_06191_), .Y(_06192_));
AND_g _27835_ (.A(_11212_), .B(_06192_), .Y(_06193_));
NAND_g _27836_ (.A(_06188_), .B(_06193_), .Y(_06194_));
NAND_g _27837_ (.A(_06184_), .B(_06194_), .Y(_06195_));
NAND_g _27838_ (.A(_00012_[3]), .B(_06195_), .Y(_06196_));
AND_g _27839_ (.A(_06174_), .B(_06196_), .Y(_06197_));
NAND_g _27840_ (.A(_00012_[4]), .B(_06197_), .Y(_06198_));
AND_g _27841_ (.A(_13409_), .B(_06198_), .Y(_06199_));
AND_g _27842_ (.A(_06152_), .B(_06199_), .Y(_06200_));
AND_g _27843_ (.A(_13613_), .B(_06200_), .Y(_06201_));
NAND_g _27844_ (.A(_13613_), .B(_06200_), .Y(_06202_));
NAND_g _27845_ (.A(reg_pc[11]), .B(_13714_), .Y(_06203_));
NAND_g _27846_ (.A(pcpi_rs1[15]), .B(_13419_), .Y(_06204_));
AND_g _27847_ (.A(_13383_), .B(_06204_), .Y(_06205_));
NAND_g _27848_ (.A(_05863_), .B(_06205_), .Y(_06206_));
NAND_g _27849_ (.A(pcpi_rs1[10]), .B(_13420_), .Y(_06207_));
AND_g _27850_ (.A(_13382_), .B(_06207_), .Y(_06208_));
NAND_g _27851_ (.A(_05866_), .B(_06208_), .Y(_06209_));
AND_g _27852_ (.A(_06206_), .B(_06209_), .Y(_06210_));
NAND_g _27853_ (.A(_13389_), .B(_06210_), .Y(_06211_));
AND_g _27854_ (.A(_06203_), .B(_06211_), .Y(_06212_));
AND_g _27855_ (.A(_13425_), .B(_06212_), .Y(_06213_));
NAND_g _27856_ (.A(_06202_), .B(_06213_), .Y(_06214_));
NOR_g _27857_ (.A(_06106_), .B(_06214_), .Y(_06215_));
NOR_g _27858_ (.A(_06101_), .B(_06215_), .Y(_01218_));
NOR_g _27859_ (.A(pcpi_rs1[12]), .B(_13425_), .Y(_06216_));
XOR_g _27860_ (.A(_13469_), .B(_13514_), .Y(_06217_));
NAND_g _27861_ (.A(_13432_), .B(_06217_), .Y(_06218_));
NOR_g _27862_ (.A(cpuregs_10[12]), .B(_00012_[2]), .Y(_06219_));
NOR_g _27863_ (.A(cpuregs_14[12]), .B(_11214_), .Y(_06220_));
NOR_g _27864_ (.A(_06219_), .B(_06220_), .Y(_06221_));
NOR_g _27865_ (.A(cpuregs_11[12]), .B(_00012_[2]), .Y(_06222_));
NAND_g _27866_ (.A(_11161_), .B(_00012_[2]), .Y(_06223_));
NAND_g _27867_ (.A(_11212_), .B(_06221_), .Y(_06224_));
NOR_g _27868_ (.A(_11212_), .B(_06222_), .Y(_06225_));
NAND_g _27869_ (.A(_06223_), .B(_06225_), .Y(_06226_));
AND_g _27870_ (.A(_00012_[3]), .B(_06226_), .Y(_06227_));
NAND_g _27871_ (.A(_06224_), .B(_06227_), .Y(_06228_));
NAND_g _27872_ (.A(cpuregs_3[12]), .B(_11214_), .Y(_06229_));
NAND_g _27873_ (.A(cpuregs_7[12]), .B(_00012_[2]), .Y(_06230_));
AND_g _27874_ (.A(_00012_[0]), .B(_06230_), .Y(_06231_));
NAND_g _27875_ (.A(_06229_), .B(_06231_), .Y(_06232_));
NAND_g _27876_ (.A(cpuregs_6[12]), .B(_00012_[2]), .Y(_06233_));
NAND_g _27877_ (.A(cpuregs_2[12]), .B(_11214_), .Y(_06234_));
AND_g _27878_ (.A(_11212_), .B(_06234_), .Y(_06235_));
NAND_g _27879_ (.A(_06233_), .B(_06235_), .Y(_06236_));
NAND_g _27880_ (.A(_06232_), .B(_06236_), .Y(_06237_));
NAND_g _27881_ (.A(_11215_), .B(_06237_), .Y(_06238_));
NAND_g _27882_ (.A(_06228_), .B(_06238_), .Y(_06239_));
NAND_g _27883_ (.A(_00012_[1]), .B(_06239_), .Y(_06240_));
NOR_g _27884_ (.A(cpuregs_9[12]), .B(_00012_[2]), .Y(_06241_));
NAND_g _27885_ (.A(_11146_), .B(_00012_[2]), .Y(_06242_));
NOR_g _27886_ (.A(cpuregs_8[12]), .B(_00012_[2]), .Y(_06243_));
NOR_g _27887_ (.A(cpuregs_12[12]), .B(_11214_), .Y(_06244_));
NOR_g _27888_ (.A(_06243_), .B(_06244_), .Y(_06245_));
NAND_g _27889_ (.A(_11212_), .B(_06245_), .Y(_06246_));
NOR_g _27890_ (.A(_11212_), .B(_06241_), .Y(_06247_));
NAND_g _27891_ (.A(_06242_), .B(_06247_), .Y(_06248_));
AND_g _27892_ (.A(_00012_[3]), .B(_06248_), .Y(_06249_));
NAND_g _27893_ (.A(_06246_), .B(_06249_), .Y(_06250_));
NAND_g _27894_ (.A(cpuregs_1[12]), .B(_11214_), .Y(_06251_));
NAND_g _27895_ (.A(cpuregs_5[12]), .B(_00012_[2]), .Y(_06252_));
AND_g _27896_ (.A(_00012_[0]), .B(_06252_), .Y(_06253_));
NAND_g _27897_ (.A(_06251_), .B(_06253_), .Y(_06254_));
NAND_g _27898_ (.A(cpuregs_4[12]), .B(_00012_[2]), .Y(_06255_));
NAND_g _27899_ (.A(cpuregs_0[12]), .B(_11214_), .Y(_06256_));
AND_g _27900_ (.A(_11212_), .B(_06256_), .Y(_06257_));
NAND_g _27901_ (.A(_06255_), .B(_06257_), .Y(_06258_));
NAND_g _27902_ (.A(_06254_), .B(_06258_), .Y(_06259_));
NAND_g _27903_ (.A(_11215_), .B(_06259_), .Y(_06260_));
NAND_g _27904_ (.A(_06250_), .B(_06260_), .Y(_06261_));
NAND_g _27905_ (.A(_11213_), .B(_06261_), .Y(_06262_));
NAND_g _27906_ (.A(cpuregs_26[12]), .B(_11214_), .Y(_06263_));
NAND_g _27907_ (.A(cpuregs_30[12]), .B(_00012_[2]), .Y(_06264_));
AND_g _27908_ (.A(_11212_), .B(_06264_), .Y(_06265_));
NAND_g _27909_ (.A(_06263_), .B(_06265_), .Y(_06266_));
NAND_g _27910_ (.A(cpuregs_31[12]), .B(_00012_[2]), .Y(_06267_));
NAND_g _27911_ (.A(cpuregs_27[12]), .B(_11214_), .Y(_06268_));
AND_g _27912_ (.A(_00012_[0]), .B(_06268_), .Y(_06269_));
NAND_g _27913_ (.A(_06267_), .B(_06269_), .Y(_06270_));
NAND_g _27914_ (.A(_06266_), .B(_06270_), .Y(_06271_));
NAND_g _27915_ (.A(_00012_[3]), .B(_06271_), .Y(_06272_));
NAND_g _27916_ (.A(cpuregs_22[12]), .B(_00012_[2]), .Y(_06273_));
NAND_g _27917_ (.A(cpuregs_18[12]), .B(_11214_), .Y(_06274_));
AND_g _27918_ (.A(_11212_), .B(_06274_), .Y(_06275_));
NAND_g _27919_ (.A(_06273_), .B(_06275_), .Y(_06276_));
NAND_g _27920_ (.A(cpuregs_23[12]), .B(_00012_[2]), .Y(_06277_));
NAND_g _27921_ (.A(cpuregs_19[12]), .B(_11214_), .Y(_06278_));
AND_g _27922_ (.A(_00012_[0]), .B(_06278_), .Y(_06279_));
NAND_g _27923_ (.A(_06277_), .B(_06279_), .Y(_06280_));
NAND_g _27924_ (.A(_06276_), .B(_06280_), .Y(_06281_));
NAND_g _27925_ (.A(_11215_), .B(_06281_), .Y(_06282_));
NAND_g _27926_ (.A(_06272_), .B(_06282_), .Y(_06283_));
NAND_g _27927_ (.A(_00012_[1]), .B(_06283_), .Y(_06284_));
NAND_g _27928_ (.A(_11028_), .B(_00012_[2]), .Y(_06285_));
NOR_g _27929_ (.A(cpuregs_17[12]), .B(_00012_[2]), .Y(_06286_));
NOR_g _27930_ (.A(_11212_), .B(_06286_), .Y(_06287_));
NAND_g _27931_ (.A(_06285_), .B(_06287_), .Y(_06288_));
NOR_g _27932_ (.A(cpuregs_16[12]), .B(_00012_[2]), .Y(_06289_));
AND_g _27933_ (.A(_11197_), .B(_00012_[2]), .Y(_06290_));
NOR_g _27934_ (.A(_06289_), .B(_06290_), .Y(_06291_));
NAND_g _27935_ (.A(_11212_), .B(_06291_), .Y(_06292_));
AND_g _27936_ (.A(_06288_), .B(_06292_), .Y(_06293_));
NAND_g _27937_ (.A(_11215_), .B(_06293_), .Y(_06294_));
NOR_g _27938_ (.A(cpuregs_24[12]), .B(_00012_[2]), .Y(_06295_));
NOR_g _27939_ (.A(cpuregs_28[12]), .B(_11214_), .Y(_06296_));
NOR_g _27940_ (.A(_06295_), .B(_06296_), .Y(_06297_));
NAND_g _27941_ (.A(_11212_), .B(_06297_), .Y(_06298_));
NAND_g _27942_ (.A(_10927_), .B(_00012_[2]), .Y(_06299_));
NOR_g _27943_ (.A(cpuregs_25[12]), .B(_00012_[2]), .Y(_06300_));
NOR_g _27944_ (.A(_11212_), .B(_06300_), .Y(_06301_));
NAND_g _27945_ (.A(_06299_), .B(_06301_), .Y(_06302_));
AND_g _27946_ (.A(_00012_[3]), .B(_06302_), .Y(_06303_));
NAND_g _27947_ (.A(_06298_), .B(_06303_), .Y(_06304_));
NAND_g _27948_ (.A(_06294_), .B(_06304_), .Y(_06305_));
NAND_g _27949_ (.A(_11213_), .B(_06305_), .Y(_06306_));
AND_g _27950_ (.A(_06284_), .B(_06306_), .Y(_06307_));
NAND_g _27951_ (.A(_00012_[4]), .B(_06307_), .Y(_06308_));
AND_g _27952_ (.A(_11216_), .B(_06262_), .Y(_06309_));
NAND_g _27953_ (.A(_06240_), .B(_06309_), .Y(_06310_));
NAND_g _27954_ (.A(_06308_), .B(_06310_), .Y(_06311_));
AND_g _27955_ (.A(_13561_), .B(_06311_), .Y(_06312_));
NAND_g _27956_ (.A(_05765_), .B(_06312_), .Y(_06313_));
NAND_g _27957_ (.A(reg_pc[12]), .B(_13714_), .Y(_06314_));
NAND_g _27958_ (.A(pcpi_rs1[16]), .B(_13419_), .Y(_06315_));
AND_g _27959_ (.A(_13383_), .B(_05978_), .Y(_06316_));
NAND_g _27960_ (.A(_06315_), .B(_06316_), .Y(_06317_));
NAND_g _27961_ (.A(pcpi_rs1[11]), .B(_13420_), .Y(_06318_));
AND_g _27962_ (.A(_13382_), .B(_06318_), .Y(_06319_));
NAND_g _27963_ (.A(_05981_), .B(_06319_), .Y(_06320_));
AND_g _27964_ (.A(_06317_), .B(_06320_), .Y(_06321_));
NAND_g _27965_ (.A(_13389_), .B(_06321_), .Y(_06322_));
AND_g _27966_ (.A(_06314_), .B(_06322_), .Y(_06323_));
AND_g _27967_ (.A(_13425_), .B(_06323_), .Y(_06324_));
AND_g _27968_ (.A(_06313_), .B(_06324_), .Y(_06325_));
AND_g _27969_ (.A(_06218_), .B(_06325_), .Y(_06326_));
NOR_g _27970_ (.A(_06216_), .B(_06326_), .Y(_01219_));
NOR_g _27971_ (.A(pcpi_rs1[13]), .B(_13425_), .Y(_06327_));
XOR_g _27972_ (.A(decoded_imm[13]), .B(pcpi_rs1[13]), .Y(_06328_));
XNOR_g _27973_ (.A(_13516_), .B(_06328_), .Y(_06329_));
NAND_g _27974_ (.A(_13432_), .B(_06329_), .Y(_06330_));
NAND_g _27975_ (.A(reg_pc[13]), .B(_13714_), .Y(_06331_));
NAND_g _27976_ (.A(pcpi_rs1[12]), .B(_13420_), .Y(_06332_));
AND_g _27977_ (.A(_05997_), .B(_06332_), .Y(_06333_));
NAND_g _27978_ (.A(_13382_), .B(_06333_), .Y(_06334_));
NAND_g _27979_ (.A(pcpi_rs1[17]), .B(_13419_), .Y(_06335_));
AND_g _27980_ (.A(_05994_), .B(_06335_), .Y(_06336_));
NAND_g _27981_ (.A(_13383_), .B(_06336_), .Y(_06337_));
AND_g _27982_ (.A(_06334_), .B(_06337_), .Y(_06338_));
NAND_g _27983_ (.A(_13389_), .B(_06338_), .Y(_06339_));
AND_g _27984_ (.A(_06331_), .B(_06339_), .Y(_06340_));
AND_g _27985_ (.A(_13425_), .B(_06340_), .Y(_06341_));
NAND_g _27986_ (.A(_11097_), .B(_00012_[2]), .Y(_06342_));
NOR_g _27987_ (.A(cpuregs_24[13]), .B(_00012_[2]), .Y(_06343_));
NOR_g _27988_ (.A(_00012_[0]), .B(_06343_), .Y(_06344_));
NAND_g _27989_ (.A(_06342_), .B(_06344_), .Y(_06345_));
NAND_g _27990_ (.A(_10928_), .B(_00012_[2]), .Y(_06346_));
NOR_g _27991_ (.A(cpuregs_25[13]), .B(_00012_[2]), .Y(_06347_));
NOR_g _27992_ (.A(_11212_), .B(_06347_), .Y(_06348_));
NAND_g _27993_ (.A(_06346_), .B(_06348_), .Y(_06349_));
NAND_g _27994_ (.A(_06345_), .B(_06349_), .Y(_06350_));
NAND_g _27995_ (.A(_00012_[3]), .B(_06350_), .Y(_06351_));
NAND_g _27996_ (.A(cpuregs_20[13]), .B(_00012_[2]), .Y(_06352_));
NAND_g _27997_ (.A(cpuregs_16[13]), .B(_11214_), .Y(_06353_));
AND_g _27998_ (.A(_06352_), .B(_06353_), .Y(_06354_));
NAND_g _27999_ (.A(_11212_), .B(_06354_), .Y(_06355_));
NAND_g _28000_ (.A(cpuregs_21[13]), .B(_00012_[2]), .Y(_06356_));
NAND_g _28001_ (.A(cpuregs_17[13]), .B(_11214_), .Y(_06357_));
AND_g _28002_ (.A(_00012_[0]), .B(_06357_), .Y(_06358_));
NAND_g _28003_ (.A(_06356_), .B(_06358_), .Y(_06359_));
AND_g _28004_ (.A(_11215_), .B(_06359_), .Y(_06360_));
NAND_g _28005_ (.A(_06355_), .B(_06360_), .Y(_06361_));
AND_g _28006_ (.A(_06351_), .B(_06361_), .Y(_06362_));
NAND_g _28007_ (.A(cpuregs_4[13]), .B(_00012_[2]), .Y(_06363_));
NAND_g _28008_ (.A(cpuregs_0[13]), .B(_11214_), .Y(_06364_));
AND_g _28009_ (.A(_11212_), .B(_06364_), .Y(_06365_));
NAND_g _28010_ (.A(_06363_), .B(_06365_), .Y(_06366_));
NAND_g _28011_ (.A(cpuregs_1[13]), .B(_11214_), .Y(_06367_));
NAND_g _28012_ (.A(cpuregs_5[13]), .B(_00012_[2]), .Y(_06368_));
AND_g _28013_ (.A(_00012_[0]), .B(_06368_), .Y(_06369_));
NAND_g _28014_ (.A(_06367_), .B(_06369_), .Y(_06370_));
NOR_g _28015_ (.A(cpuregs_8[13]), .B(_00012_[2]), .Y(_06371_));
NOR_g _28016_ (.A(cpuregs_12[13]), .B(_11214_), .Y(_06372_));
NOR_g _28017_ (.A(_06371_), .B(_06372_), .Y(_06373_));
NOR_g _28018_ (.A(cpuregs_9[13]), .B(_00012_[2]), .Y(_06374_));
NAND_g _28019_ (.A(_11147_), .B(_00012_[2]), .Y(_06375_));
NAND_g _28020_ (.A(_06366_), .B(_06370_), .Y(_06376_));
NAND_g _28021_ (.A(_11215_), .B(_06376_), .Y(_06377_));
NAND_g _28022_ (.A(_11212_), .B(_06373_), .Y(_06378_));
NOR_g _28023_ (.A(_11212_), .B(_06374_), .Y(_06379_));
NAND_g _28024_ (.A(_06375_), .B(_06379_), .Y(_06380_));
AND_g _28025_ (.A(_00012_[3]), .B(_06380_), .Y(_06381_));
NAND_g _28026_ (.A(_06378_), .B(_06381_), .Y(_06382_));
NAND_g _28027_ (.A(_06377_), .B(_06382_), .Y(_06383_));
NAND_g _28028_ (.A(_11174_), .B(_00012_[2]), .Y(_06384_));
NOR_g _28029_ (.A(cpuregs_26[13]), .B(_00012_[2]), .Y(_06385_));
NOR_g _28030_ (.A(_00012_[0]), .B(_06385_), .Y(_06386_));
NAND_g _28031_ (.A(_06384_), .B(_06386_), .Y(_06387_));
NAND_g _28032_ (.A(_11090_), .B(_00012_[2]), .Y(_06388_));
NOR_g _28033_ (.A(cpuregs_27[13]), .B(_00012_[2]), .Y(_06389_));
NOR_g _28034_ (.A(_11212_), .B(_06389_), .Y(_06390_));
NAND_g _28035_ (.A(_06388_), .B(_06390_), .Y(_06391_));
NAND_g _28036_ (.A(_06387_), .B(_06391_), .Y(_06392_));
NAND_g _28037_ (.A(_00012_[3]), .B(_06392_), .Y(_06393_));
NAND_g _28038_ (.A(cpuregs_22[13]), .B(_00012_[2]), .Y(_06394_));
NAND_g _28039_ (.A(cpuregs_18[13]), .B(_11214_), .Y(_06395_));
AND_g _28040_ (.A(_06394_), .B(_06395_), .Y(_06396_));
NAND_g _28041_ (.A(_11212_), .B(_06396_), .Y(_06397_));
NAND_g _28042_ (.A(cpuregs_23[13]), .B(_00012_[2]), .Y(_06398_));
NAND_g _28043_ (.A(cpuregs_19[13]), .B(_11214_), .Y(_06399_));
AND_g _28044_ (.A(_00012_[0]), .B(_06399_), .Y(_06400_));
NAND_g _28045_ (.A(_06398_), .B(_06400_), .Y(_06401_));
AND_g _28046_ (.A(_11215_), .B(_06401_), .Y(_06402_));
NAND_g _28047_ (.A(_06397_), .B(_06402_), .Y(_06403_));
AND_g _28048_ (.A(_06393_), .B(_06403_), .Y(_06404_));
NAND_g _28049_ (.A(_00012_[1]), .B(_06404_), .Y(_06405_));
NAND_g _28050_ (.A(_11213_), .B(_06362_), .Y(_06406_));
AND_g _28051_ (.A(_00012_[4]), .B(_06406_), .Y(_06407_));
NAND_g _28052_ (.A(_06405_), .B(_06407_), .Y(_06408_));
NAND_g _28053_ (.A(_11213_), .B(_06383_), .Y(_06409_));
NAND_g _28054_ (.A(cpuregs_6[13]), .B(_00012_[2]), .Y(_06410_));
NAND_g _28055_ (.A(cpuregs_2[13]), .B(_11214_), .Y(_06411_));
AND_g _28056_ (.A(_06410_), .B(_06411_), .Y(_06412_));
NAND_g _28057_ (.A(_11212_), .B(_06412_), .Y(_06413_));
NAND_g _28058_ (.A(cpuregs_7[13]), .B(_00012_[2]), .Y(_06414_));
NAND_g _28059_ (.A(cpuregs_3[13]), .B(_11214_), .Y(_06415_));
AND_g _28060_ (.A(_00012_[0]), .B(_06415_), .Y(_06416_));
NAND_g _28061_ (.A(_06414_), .B(_06416_), .Y(_06417_));
AND_g _28062_ (.A(_11215_), .B(_06417_), .Y(_06418_));
NAND_g _28063_ (.A(_06413_), .B(_06418_), .Y(_06419_));
NOR_g _28064_ (.A(cpuregs_11[13]), .B(_00012_[2]), .Y(_06420_));
NOT_g _28065_ (.A(_06420_), .Y(_06421_));
NAND_g _28066_ (.A(_11162_), .B(_00012_[2]), .Y(_06422_));
AND_g _28067_ (.A(_00012_[0]), .B(_06422_), .Y(_06423_));
NAND_g _28068_ (.A(_06421_), .B(_06423_), .Y(_06424_));
NOR_g _28069_ (.A(cpuregs_10[13]), .B(_00012_[2]), .Y(_06425_));
NOR_g _28070_ (.A(cpuregs_14[13]), .B(_11214_), .Y(_06426_));
NOR_g _28071_ (.A(_06425_), .B(_06426_), .Y(_06427_));
NAND_g _28072_ (.A(_11212_), .B(_06427_), .Y(_06428_));
NAND_g _28073_ (.A(_06424_), .B(_06428_), .Y(_06429_));
NAND_g _28074_ (.A(_00012_[3]), .B(_06429_), .Y(_06430_));
AND_g _28075_ (.A(_06419_), .B(_06430_), .Y(_06431_));
NAND_g _28076_ (.A(_00012_[1]), .B(_06431_), .Y(_06432_));
AND_g _28077_ (.A(_06409_), .B(_06432_), .Y(_06433_));
NAND_g _28078_ (.A(_11216_), .B(_06433_), .Y(_06434_));
NAND_g _28079_ (.A(_06408_), .B(_06434_), .Y(_06435_));
AND_g _28080_ (.A(_13561_), .B(_06435_), .Y(_06436_));
NAND_g _28081_ (.A(_05765_), .B(_06436_), .Y(_06437_));
AND_g _28082_ (.A(_06341_), .B(_06437_), .Y(_06438_));
AND_g _28083_ (.A(_06330_), .B(_06438_), .Y(_06439_));
NOR_g _28084_ (.A(_06327_), .B(_06439_), .Y(_01220_));
NOR_g _28085_ (.A(pcpi_rs1[14]), .B(_13425_), .Y(_06440_));
NAND_g _28086_ (.A(_11129_), .B(_00012_[2]), .Y(_06441_));
NOR_g _28087_ (.A(cpuregs_3[14]), .B(_00012_[2]), .Y(_06442_));
NOR_g _28088_ (.A(_11212_), .B(_06442_), .Y(_06443_));
NAND_g _28089_ (.A(_06441_), .B(_06443_), .Y(_06444_));
NOR_g _28090_ (.A(cpuregs_2[14]), .B(_00012_[2]), .Y(_06445_));
AND_g _28091_ (.A(_10943_), .B(_00012_[2]), .Y(_06446_));
NOR_g _28092_ (.A(_06445_), .B(_06446_), .Y(_06447_));
NAND_g _28093_ (.A(_11212_), .B(_06447_), .Y(_06448_));
AND_g _28094_ (.A(_06444_), .B(_06448_), .Y(_06449_));
NAND_g _28095_ (.A(_11113_), .B(_00012_[2]), .Y(_06450_));
NOR_g _28096_ (.A(cpuregs_1[14]), .B(_00012_[2]), .Y(_06451_));
NOR_g _28097_ (.A(_11212_), .B(_06451_), .Y(_06452_));
NAND_g _28098_ (.A(_06450_), .B(_06452_), .Y(_06453_));
NOR_g _28099_ (.A(cpuregs_0[14]), .B(_00012_[2]), .Y(_06454_));
AND_g _28100_ (.A(_10955_), .B(_00012_[2]), .Y(_06455_));
NOR_g _28101_ (.A(_06454_), .B(_06455_), .Y(_06456_));
NAND_g _28102_ (.A(_11212_), .B(_06456_), .Y(_06457_));
AND_g _28103_ (.A(_06453_), .B(_06457_), .Y(_06458_));
NAND_g _28104_ (.A(_00012_[1]), .B(_06449_), .Y(_06459_));
NAND_g _28105_ (.A(_11213_), .B(_06458_), .Y(_06460_));
AND_g _28106_ (.A(_06459_), .B(_06460_), .Y(_06461_));
NAND_g _28107_ (.A(_11215_), .B(_06461_), .Y(_06462_));
NAND_g _28108_ (.A(cpuregs_13[14]), .B(_00012_[0]), .Y(_06463_));
NAND_g _28109_ (.A(cpuregs_12[14]), .B(_11212_), .Y(_06464_));
AND_g _28110_ (.A(_00012_[2]), .B(_06464_), .Y(_06465_));
NAND_g _28111_ (.A(_06463_), .B(_06465_), .Y(_06466_));
NAND_g _28112_ (.A(cpuregs_9[14]), .B(_00012_[0]), .Y(_06467_));
NAND_g _28113_ (.A(cpuregs_8[14]), .B(_11212_), .Y(_06468_));
AND_g _28114_ (.A(_11214_), .B(_06468_), .Y(_06469_));
NAND_g _28115_ (.A(_06467_), .B(_06469_), .Y(_06470_));
AND_g _28116_ (.A(_11213_), .B(_06470_), .Y(_06471_));
NAND_g _28117_ (.A(_06466_), .B(_06471_), .Y(_06472_));
NAND_g _28118_ (.A(cpuregs_15[14]), .B(_00012_[0]), .Y(_06473_));
NAND_g _28119_ (.A(cpuregs_14[14]), .B(_11212_), .Y(_06474_));
AND_g _28120_ (.A(_00012_[2]), .B(_06474_), .Y(_06475_));
NAND_g _28121_ (.A(_06473_), .B(_06475_), .Y(_06476_));
NAND_g _28122_ (.A(cpuregs_11[14]), .B(_00012_[0]), .Y(_06477_));
NAND_g _28123_ (.A(cpuregs_10[14]), .B(_11212_), .Y(_06478_));
AND_g _28124_ (.A(_11214_), .B(_06478_), .Y(_06479_));
NAND_g _28125_ (.A(_06477_), .B(_06479_), .Y(_06480_));
AND_g _28126_ (.A(_00012_[1]), .B(_06480_), .Y(_06481_));
NAND_g _28127_ (.A(_06476_), .B(_06481_), .Y(_06482_));
NAND_g _28128_ (.A(_06472_), .B(_06482_), .Y(_06483_));
NAND_g _28129_ (.A(_00012_[3]), .B(_06483_), .Y(_06484_));
AND_g _28130_ (.A(_06462_), .B(_06484_), .Y(_06485_));
NAND_g _28131_ (.A(_11216_), .B(_06485_), .Y(_06486_));
NAND_g _28132_ (.A(cpuregs_20[14]), .B(_11213_), .Y(_06487_));
NAND_g _28133_ (.A(cpuregs_22[14]), .B(_00012_[1]), .Y(_06488_));
AND_g _28134_ (.A(_00012_[2]), .B(_06488_), .Y(_06489_));
NAND_g _28135_ (.A(_06487_), .B(_06489_), .Y(_06490_));
NAND_g _28136_ (.A(cpuregs_16[14]), .B(_11213_), .Y(_06491_));
NAND_g _28137_ (.A(cpuregs_18[14]), .B(_00012_[1]), .Y(_06492_));
AND_g _28138_ (.A(_11214_), .B(_06492_), .Y(_06493_));
NAND_g _28139_ (.A(_06491_), .B(_06493_), .Y(_06494_));
AND_g _28140_ (.A(_11212_), .B(_06494_), .Y(_06495_));
NAND_g _28141_ (.A(_06490_), .B(_06495_), .Y(_06496_));
NAND_g _28142_ (.A(cpuregs_21[14]), .B(_11213_), .Y(_06497_));
NAND_g _28143_ (.A(cpuregs_23[14]), .B(_00012_[1]), .Y(_06498_));
AND_g _28144_ (.A(_00012_[2]), .B(_06498_), .Y(_06499_));
NAND_g _28145_ (.A(_06497_), .B(_06499_), .Y(_06500_));
NAND_g _28146_ (.A(cpuregs_17[14]), .B(_11213_), .Y(_06501_));
NAND_g _28147_ (.A(cpuregs_19[14]), .B(_00012_[1]), .Y(_06502_));
AND_g _28148_ (.A(_11214_), .B(_06502_), .Y(_06503_));
NAND_g _28149_ (.A(_06501_), .B(_06503_), .Y(_06504_));
AND_g _28150_ (.A(_00012_[0]), .B(_06504_), .Y(_06505_));
NAND_g _28151_ (.A(_06500_), .B(_06505_), .Y(_06506_));
NAND_g _28152_ (.A(_06496_), .B(_06506_), .Y(_06507_));
NAND_g _28153_ (.A(_11215_), .B(_06507_), .Y(_06508_));
NAND_g _28154_ (.A(cpuregs_26[14]), .B(_11214_), .Y(_06509_));
NAND_g _28155_ (.A(cpuregs_30[14]), .B(_00012_[2]), .Y(_06510_));
AND_g _28156_ (.A(_00012_[1]), .B(_06510_), .Y(_06511_));
NAND_g _28157_ (.A(_06509_), .B(_06511_), .Y(_06512_));
NAND_g _28158_ (.A(cpuregs_24[14]), .B(_11214_), .Y(_06513_));
NAND_g _28159_ (.A(cpuregs_28[14]), .B(_00012_[2]), .Y(_06514_));
AND_g _28160_ (.A(_11213_), .B(_06514_), .Y(_06515_));
NAND_g _28161_ (.A(_06513_), .B(_06515_), .Y(_06516_));
AND_g _28162_ (.A(_11212_), .B(_06516_), .Y(_06517_));
NAND_g _28163_ (.A(_06512_), .B(_06517_), .Y(_06518_));
NAND_g _28164_ (.A(cpuregs_27[14]), .B(_11214_), .Y(_06519_));
NAND_g _28165_ (.A(cpuregs_31[14]), .B(_00012_[2]), .Y(_06520_));
AND_g _28166_ (.A(_00012_[1]), .B(_06520_), .Y(_06521_));
NAND_g _28167_ (.A(_06519_), .B(_06521_), .Y(_06522_));
NAND_g _28168_ (.A(cpuregs_29[14]), .B(_00012_[2]), .Y(_06523_));
NAND_g _28169_ (.A(cpuregs_25[14]), .B(_11214_), .Y(_06524_));
AND_g _28170_ (.A(_11213_), .B(_06524_), .Y(_06525_));
NAND_g _28171_ (.A(_06523_), .B(_06525_), .Y(_06526_));
AND_g _28172_ (.A(_00012_[0]), .B(_06526_), .Y(_06527_));
NAND_g _28173_ (.A(_06522_), .B(_06527_), .Y(_06528_));
NAND_g _28174_ (.A(_06518_), .B(_06528_), .Y(_06529_));
NAND_g _28175_ (.A(_00012_[3]), .B(_06529_), .Y(_06530_));
AND_g _28176_ (.A(_00012_[4]), .B(_06508_), .Y(_06531_));
NAND_g _28177_ (.A(_06530_), .B(_06531_), .Y(_06532_));
AND_g _28178_ (.A(_13409_), .B(_06532_), .Y(_06533_));
AND_g _28179_ (.A(_06486_), .B(_06533_), .Y(_06534_));
AND_g _28180_ (.A(_13613_), .B(_06534_), .Y(_06535_));
NAND_g _28181_ (.A(reg_pc[14]), .B(_13714_), .Y(_06536_));
NAND_g _28182_ (.A(pcpi_rs1[18]), .B(_13419_), .Y(_06537_));
AND_g _28183_ (.A(_13383_), .B(_06207_), .Y(_06538_));
NAND_g _28184_ (.A(_06537_), .B(_06538_), .Y(_06539_));
NAND_g _28185_ (.A(pcpi_rs1[13]), .B(_13420_), .Y(_06540_));
AND_g _28186_ (.A(_13382_), .B(_06540_), .Y(_06541_));
NAND_g _28187_ (.A(_06204_), .B(_06541_), .Y(_06542_));
AND_g _28188_ (.A(_06539_), .B(_06542_), .Y(_06543_));
NAND_g _28189_ (.A(_13389_), .B(_06543_), .Y(_06544_));
AND_g _28190_ (.A(_06536_), .B(_06544_), .Y(_06545_));
NAND_g _28191_ (.A(_13425_), .B(_06545_), .Y(_06546_));
NOR_g _28192_ (.A(_06535_), .B(_06546_), .Y(_06547_));
XOR_g _28193_ (.A(_13465_), .B(_13518_), .Y(_06548_));
NAND_g _28194_ (.A(_13432_), .B(_06548_), .Y(_06549_));
AND_g _28195_ (.A(_06547_), .B(_06549_), .Y(_06550_));
NOR_g _28196_ (.A(_06440_), .B(_06550_), .Y(_01221_));
NOR_g _28197_ (.A(pcpi_rs1[15]), .B(_13425_), .Y(_06551_));
XOR_g _28198_ (.A(decoded_imm[15]), .B(pcpi_rs1[15]), .Y(_06552_));
XNOR_g _28199_ (.A(_13520_), .B(_06552_), .Y(_06553_));
NAND_g _28200_ (.A(_13432_), .B(_06553_), .Y(_06554_));
NAND_g _28201_ (.A(reg_pc[15]), .B(_13714_), .Y(_06555_));
NAND_g _28202_ (.A(pcpi_rs1[19]), .B(_13419_), .Y(_06556_));
AND_g _28203_ (.A(_13383_), .B(_06318_), .Y(_06557_));
NAND_g _28204_ (.A(_06556_), .B(_06557_), .Y(_06558_));
NAND_g _28205_ (.A(pcpi_rs1[14]), .B(_13420_), .Y(_06559_));
AND_g _28206_ (.A(_13382_), .B(_06559_), .Y(_06560_));
NAND_g _28207_ (.A(_06315_), .B(_06560_), .Y(_06561_));
AND_g _28208_ (.A(_06558_), .B(_06561_), .Y(_06562_));
NAND_g _28209_ (.A(_13389_), .B(_06562_), .Y(_06563_));
AND_g _28210_ (.A(_06555_), .B(_06563_), .Y(_06564_));
AND_g _28211_ (.A(_13425_), .B(_06564_), .Y(_06565_));
NAND_g _28212_ (.A(cpuregs_23[15]), .B(_00012_[0]), .Y(_06566_));
NAND_g _28213_ (.A(cpuregs_22[15]), .B(_11212_), .Y(_06567_));
AND_g _28214_ (.A(_00012_[2]), .B(_06567_), .Y(_06568_));
NAND_g _28215_ (.A(_06566_), .B(_06568_), .Y(_06569_));
NAND_g _28216_ (.A(cpuregs_19[15]), .B(_00012_[0]), .Y(_06570_));
NAND_g _28217_ (.A(cpuregs_18[15]), .B(_11212_), .Y(_06571_));
AND_g _28218_ (.A(_11214_), .B(_06571_), .Y(_06572_));
NAND_g _28219_ (.A(_06570_), .B(_06572_), .Y(_06573_));
AND_g _28220_ (.A(_11215_), .B(_06573_), .Y(_06574_));
NAND_g _28221_ (.A(_06569_), .B(_06574_), .Y(_06575_));
NAND_g _28222_ (.A(cpuregs_31[15]), .B(_00012_[0]), .Y(_06576_));
NAND_g _28223_ (.A(cpuregs_30[15]), .B(_11212_), .Y(_06577_));
AND_g _28224_ (.A(_00012_[2]), .B(_06577_), .Y(_06578_));
NAND_g _28225_ (.A(_06576_), .B(_06578_), .Y(_06579_));
NAND_g _28226_ (.A(cpuregs_27[15]), .B(_00012_[0]), .Y(_06580_));
NAND_g _28227_ (.A(cpuregs_26[15]), .B(_11212_), .Y(_06581_));
AND_g _28228_ (.A(_11214_), .B(_06581_), .Y(_06582_));
NAND_g _28229_ (.A(_06580_), .B(_06582_), .Y(_06583_));
AND_g _28230_ (.A(_00012_[3]), .B(_06583_), .Y(_06584_));
NAND_g _28231_ (.A(_06579_), .B(_06584_), .Y(_06585_));
NAND_g _28232_ (.A(_06575_), .B(_06585_), .Y(_06586_));
NAND_g _28233_ (.A(_00012_[4]), .B(_06586_), .Y(_06587_));
NAND_g _28234_ (.A(cpuregs_6[15]), .B(_00012_[2]), .Y(_06588_));
NAND_g _28235_ (.A(cpuregs_2[15]), .B(_11214_), .Y(_06589_));
AND_g _28236_ (.A(_11212_), .B(_06589_), .Y(_06590_));
NAND_g _28237_ (.A(_06588_), .B(_06590_), .Y(_06591_));
NAND_g _28238_ (.A(cpuregs_3[15]), .B(_11214_), .Y(_06592_));
NAND_g _28239_ (.A(cpuregs_7[15]), .B(_00012_[2]), .Y(_06593_));
AND_g _28240_ (.A(_00012_[0]), .B(_06593_), .Y(_06594_));
NAND_g _28241_ (.A(_06592_), .B(_06594_), .Y(_06595_));
NOR_g _28242_ (.A(cpuregs_10[15]), .B(_00012_[2]), .Y(_06596_));
NOR_g _28243_ (.A(cpuregs_14[15]), .B(_11214_), .Y(_06597_));
NOR_g _28244_ (.A(_06596_), .B(_06597_), .Y(_06598_));
NOR_g _28245_ (.A(cpuregs_11[15]), .B(_00012_[2]), .Y(_06599_));
NAND_g _28246_ (.A(_11163_), .B(_00012_[2]), .Y(_06600_));
NAND_g _28247_ (.A(_06591_), .B(_06595_), .Y(_06601_));
NAND_g _28248_ (.A(_11215_), .B(_06601_), .Y(_06602_));
NAND_g _28249_ (.A(_11212_), .B(_06598_), .Y(_06603_));
NOR_g _28250_ (.A(_11212_), .B(_06599_), .Y(_06604_));
NAND_g _28251_ (.A(_06600_), .B(_06604_), .Y(_06605_));
AND_g _28252_ (.A(_00012_[3]), .B(_06605_), .Y(_06606_));
NAND_g _28253_ (.A(_06603_), .B(_06606_), .Y(_06607_));
AND_g _28254_ (.A(_06602_), .B(_06607_), .Y(_06608_));
NAND_g _28255_ (.A(_11216_), .B(_06608_), .Y(_06609_));
NAND_g _28256_ (.A(_06587_), .B(_06609_), .Y(_06610_));
NAND_g _28257_ (.A(_00012_[1]), .B(_06610_), .Y(_06611_));
NAND_g _28258_ (.A(cpuregs_4[15]), .B(_00012_[2]), .Y(_06612_));
NAND_g _28259_ (.A(cpuregs_0[15]), .B(_11214_), .Y(_06613_));
AND_g _28260_ (.A(_11212_), .B(_06613_), .Y(_06614_));
NAND_g _28261_ (.A(_06612_), .B(_06614_), .Y(_06615_));
NAND_g _28262_ (.A(cpuregs_1[15]), .B(_11214_), .Y(_06616_));
NAND_g _28263_ (.A(cpuregs_5[15]), .B(_00012_[2]), .Y(_06617_));
AND_g _28264_ (.A(_00012_[0]), .B(_06617_), .Y(_06618_));
NAND_g _28265_ (.A(_06616_), .B(_06618_), .Y(_06619_));
NOR_g _28266_ (.A(cpuregs_8[15]), .B(_00012_[2]), .Y(_06620_));
AND_g _28267_ (.A(_11119_), .B(_00012_[2]), .Y(_06621_));
NOR_g _28268_ (.A(_06620_), .B(_06621_), .Y(_06622_));
NOR_g _28269_ (.A(cpuregs_9[15]), .B(_00012_[2]), .Y(_06623_));
NAND_g _28270_ (.A(_11148_), .B(_00012_[2]), .Y(_06624_));
NAND_g _28271_ (.A(_06615_), .B(_06619_), .Y(_06625_));
NAND_g _28272_ (.A(_11215_), .B(_06625_), .Y(_06626_));
NAND_g _28273_ (.A(_11212_), .B(_06622_), .Y(_06627_));
NOR_g _28274_ (.A(_11212_), .B(_06623_), .Y(_06628_));
NAND_g _28275_ (.A(_06624_), .B(_06628_), .Y(_06629_));
AND_g _28276_ (.A(_00012_[3]), .B(_06629_), .Y(_06630_));
NAND_g _28277_ (.A(_06627_), .B(_06630_), .Y(_06631_));
AND_g _28278_ (.A(_06626_), .B(_06631_), .Y(_06632_));
NAND_g _28279_ (.A(_11216_), .B(_06632_), .Y(_06633_));
NAND_g _28280_ (.A(cpuregs_25[15]), .B(_00012_[3]), .Y(_06634_));
NAND_g _28281_ (.A(cpuregs_17[15]), .B(_11215_), .Y(_06635_));
NAND_g _28282_ (.A(_06634_), .B(_06635_), .Y(_06636_));
NAND_g _28283_ (.A(_11214_), .B(_06636_), .Y(_06637_));
NAND_g _28284_ (.A(cpuregs_29[15]), .B(_00012_[3]), .Y(_06638_));
NAND_g _28285_ (.A(cpuregs_21[15]), .B(_11215_), .Y(_06639_));
NAND_g _28286_ (.A(_06638_), .B(_06639_), .Y(_06640_));
NAND_g _28287_ (.A(_00012_[2]), .B(_06640_), .Y(_06641_));
AND_g _28288_ (.A(_00012_[0]), .B(_06641_), .Y(_06642_));
NAND_g _28289_ (.A(_06637_), .B(_06642_), .Y(_06643_));
NAND_g _28290_ (.A(cpuregs_24[15]), .B(_00012_[3]), .Y(_06644_));
NAND_g _28291_ (.A(cpuregs_16[15]), .B(_11215_), .Y(_06645_));
NAND_g _28292_ (.A(_06644_), .B(_06645_), .Y(_06646_));
NAND_g _28293_ (.A(_11214_), .B(_06646_), .Y(_06647_));
NAND_g _28294_ (.A(cpuregs_28[15]), .B(_00012_[3]), .Y(_06648_));
NAND_g _28295_ (.A(cpuregs_20[15]), .B(_11215_), .Y(_06649_));
NAND_g _28296_ (.A(_06648_), .B(_06649_), .Y(_06650_));
NAND_g _28297_ (.A(_00012_[2]), .B(_06650_), .Y(_06651_));
AND_g _28298_ (.A(_11212_), .B(_06651_), .Y(_06652_));
NAND_g _28299_ (.A(_06647_), .B(_06652_), .Y(_06653_));
AND_g _28300_ (.A(_00012_[4]), .B(_06653_), .Y(_06654_));
NAND_g _28301_ (.A(_06643_), .B(_06654_), .Y(_06655_));
NAND_g _28302_ (.A(_06633_), .B(_06655_), .Y(_06656_));
NAND_g _28303_ (.A(_11213_), .B(_06656_), .Y(_06657_));
NAND_g _28304_ (.A(_06611_), .B(_06657_), .Y(_06658_));
AND_g _28305_ (.A(_13561_), .B(_06658_), .Y(_06659_));
NAND_g _28306_ (.A(_05765_), .B(_06659_), .Y(_06660_));
AND_g _28307_ (.A(_06565_), .B(_06660_), .Y(_06661_));
AND_g _28308_ (.A(_06554_), .B(_06661_), .Y(_06662_));
NOR_g _28309_ (.A(_06551_), .B(_06662_), .Y(_01222_));
NOR_g _28310_ (.A(pcpi_rs1[16]), .B(_13425_), .Y(_06663_));
XOR_g _28311_ (.A(_13461_), .B(_13522_), .Y(_06664_));
NAND_g _28312_ (.A(_13432_), .B(_06664_), .Y(_06665_));
NAND_g _28313_ (.A(reg_pc[16]), .B(_13714_), .Y(_06666_));
NAND_g _28314_ (.A(pcpi_rs1[15]), .B(_13420_), .Y(_06667_));
AND_g _28315_ (.A(_06335_), .B(_06667_), .Y(_06668_));
NAND_g _28316_ (.A(_13382_), .B(_06668_), .Y(_06669_));
NAND_g _28317_ (.A(pcpi_rs1[20]), .B(_13419_), .Y(_06670_));
AND_g _28318_ (.A(_06332_), .B(_06670_), .Y(_06671_));
NAND_g _28319_ (.A(_13383_), .B(_06671_), .Y(_06672_));
AND_g _28320_ (.A(_06669_), .B(_06672_), .Y(_06673_));
NAND_g _28321_ (.A(_13389_), .B(_06673_), .Y(_06674_));
AND_g _28322_ (.A(_06666_), .B(_06674_), .Y(_06675_));
AND_g _28323_ (.A(_13425_), .B(_06675_), .Y(_06676_));
NAND_g _28324_ (.A(cpuregs_19[16]), .B(_11214_), .Y(_06677_));
NAND_g _28325_ (.A(cpuregs_23[16]), .B(_00012_[2]), .Y(_06678_));
AND_g _28326_ (.A(_00012_[0]), .B(_06678_), .Y(_06679_));
NAND_g _28327_ (.A(_06677_), .B(_06679_), .Y(_06680_));
NAND_g _28328_ (.A(cpuregs_18[16]), .B(_11214_), .Y(_06681_));
NAND_g _28329_ (.A(cpuregs_22[16]), .B(_00012_[2]), .Y(_06682_));
AND_g _28330_ (.A(_11212_), .B(_06682_), .Y(_06683_));
NAND_g _28331_ (.A(_06681_), .B(_06683_), .Y(_06684_));
AND_g _28332_ (.A(_11215_), .B(_06684_), .Y(_06685_));
NAND_g _28333_ (.A(_06680_), .B(_06685_), .Y(_06686_));
NAND_g _28334_ (.A(cpuregs_27[16]), .B(_11214_), .Y(_06687_));
NAND_g _28335_ (.A(cpuregs_31[16]), .B(_00012_[2]), .Y(_06688_));
AND_g _28336_ (.A(_00012_[0]), .B(_06688_), .Y(_06689_));
NAND_g _28337_ (.A(_06687_), .B(_06689_), .Y(_06690_));
NAND_g _28338_ (.A(cpuregs_26[16]), .B(_11214_), .Y(_06691_));
NAND_g _28339_ (.A(cpuregs_30[16]), .B(_00012_[2]), .Y(_06692_));
AND_g _28340_ (.A(_11212_), .B(_06692_), .Y(_06693_));
NAND_g _28341_ (.A(_06691_), .B(_06693_), .Y(_06694_));
AND_g _28342_ (.A(_00012_[3]), .B(_06694_), .Y(_06695_));
NAND_g _28343_ (.A(_06690_), .B(_06695_), .Y(_06696_));
NAND_g _28344_ (.A(_06686_), .B(_06696_), .Y(_06697_));
NAND_g _28345_ (.A(_00012_[1]), .B(_06697_), .Y(_06698_));
NAND_g _28346_ (.A(cpuregs_21[16]), .B(_00012_[2]), .Y(_06699_));
NAND_g _28347_ (.A(cpuregs_17[16]), .B(_11214_), .Y(_06700_));
AND_g _28348_ (.A(_00012_[0]), .B(_06700_), .Y(_06701_));
NAND_g _28349_ (.A(_06699_), .B(_06701_), .Y(_06702_));
NAND_g _28350_ (.A(cpuregs_20[16]), .B(_00012_[2]), .Y(_06703_));
NAND_g _28351_ (.A(cpuregs_16[16]), .B(_11214_), .Y(_06704_));
AND_g _28352_ (.A(_11212_), .B(_06704_), .Y(_06705_));
NAND_g _28353_ (.A(_06703_), .B(_06705_), .Y(_06706_));
AND_g _28354_ (.A(_11215_), .B(_06706_), .Y(_06707_));
NAND_g _28355_ (.A(_06702_), .B(_06707_), .Y(_06708_));
NAND_g _28356_ (.A(cpuregs_25[16]), .B(_11214_), .Y(_06709_));
NAND_g _28357_ (.A(cpuregs_29[16]), .B(_00012_[2]), .Y(_06710_));
AND_g _28358_ (.A(_00012_[0]), .B(_06710_), .Y(_06711_));
NAND_g _28359_ (.A(_06709_), .B(_06711_), .Y(_06712_));
NAND_g _28360_ (.A(cpuregs_24[16]), .B(_11214_), .Y(_06713_));
NAND_g _28361_ (.A(cpuregs_28[16]), .B(_00012_[2]), .Y(_06714_));
AND_g _28362_ (.A(_11212_), .B(_06714_), .Y(_06715_));
NAND_g _28363_ (.A(_06713_), .B(_06715_), .Y(_06716_));
AND_g _28364_ (.A(_00012_[3]), .B(_06716_), .Y(_06717_));
NAND_g _28365_ (.A(_06712_), .B(_06717_), .Y(_06718_));
NAND_g _28366_ (.A(_06708_), .B(_06718_), .Y(_06719_));
NAND_g _28367_ (.A(_11213_), .B(_06719_), .Y(_06720_));
AND_g _28368_ (.A(_06698_), .B(_06720_), .Y(_06721_));
NAND_g _28369_ (.A(cpuregs_6[16]), .B(_00012_[2]), .Y(_06722_));
NAND_g _28370_ (.A(cpuregs_2[16]), .B(_11214_), .Y(_06723_));
AND_g _28371_ (.A(_11212_), .B(_06723_), .Y(_06724_));
NAND_g _28372_ (.A(_06722_), .B(_06724_), .Y(_06725_));
NAND_g _28373_ (.A(cpuregs_3[16]), .B(_11214_), .Y(_06726_));
NAND_g _28374_ (.A(cpuregs_7[16]), .B(_00012_[2]), .Y(_06727_));
AND_g _28375_ (.A(_00012_[0]), .B(_06727_), .Y(_06728_));
NAND_g _28376_ (.A(_06726_), .B(_06728_), .Y(_06729_));
NAND_g _28377_ (.A(_06725_), .B(_06729_), .Y(_06730_));
NAND_g _28378_ (.A(_11103_), .B(_00012_[2]), .Y(_06731_));
NOR_g _28379_ (.A(cpuregs_10[16]), .B(_00012_[2]), .Y(_06732_));
NOR_g _28380_ (.A(_00012_[0]), .B(_06732_), .Y(_06733_));
AND_g _28381_ (.A(_06731_), .B(_06733_), .Y(_06734_));
NOR_g _28382_ (.A(cpuregs_11[16]), .B(_00012_[2]), .Y(_06735_));
NAND_g _28383_ (.A(_11164_), .B(_00012_[2]), .Y(_06736_));
NOR_g _28384_ (.A(_11212_), .B(_06735_), .Y(_06737_));
AND_g _28385_ (.A(_06736_), .B(_06737_), .Y(_06738_));
NOR_g _28386_ (.A(_06734_), .B(_06738_), .Y(_06739_));
NAND_g _28387_ (.A(_11215_), .B(_06730_), .Y(_06740_));
NAND_g _28388_ (.A(_00012_[3]), .B(_06739_), .Y(_06741_));
AND_g _28389_ (.A(_06740_), .B(_06741_), .Y(_06742_));
NAND_g _28390_ (.A(_00012_[1]), .B(_06742_), .Y(_06743_));
NAND_g _28391_ (.A(cpuregs_5[16]), .B(_00012_[2]), .Y(_06744_));
NAND_g _28392_ (.A(cpuregs_1[16]), .B(_11214_), .Y(_06745_));
NAND_g _28393_ (.A(_06744_), .B(_06745_), .Y(_06746_));
NAND_g _28394_ (.A(_00012_[0]), .B(_06746_), .Y(_06747_));
NAND_g _28395_ (.A(cpuregs_4[16]), .B(_00012_[2]), .Y(_06748_));
NAND_g _28396_ (.A(cpuregs_0[16]), .B(_11214_), .Y(_06749_));
NAND_g _28397_ (.A(_06748_), .B(_06749_), .Y(_06750_));
NAND_g _28398_ (.A(_11212_), .B(_06750_), .Y(_06751_));
NAND_g _28399_ (.A(_06747_), .B(_06751_), .Y(_06752_));
NAND_g _28400_ (.A(_11215_), .B(_06752_), .Y(_06753_));
NAND_g _28401_ (.A(cpuregs_13[16]), .B(_00012_[2]), .Y(_06754_));
NAND_g _28402_ (.A(cpuregs_9[16]), .B(_11214_), .Y(_06755_));
NAND_g _28403_ (.A(_06754_), .B(_06755_), .Y(_06756_));
NAND_g _28404_ (.A(_00012_[0]), .B(_06756_), .Y(_06757_));
NAND_g _28405_ (.A(cpuregs_12[16]), .B(_00012_[2]), .Y(_06758_));
NAND_g _28406_ (.A(cpuregs_8[16]), .B(_11214_), .Y(_06759_));
NAND_g _28407_ (.A(_06758_), .B(_06759_), .Y(_06760_));
NAND_g _28408_ (.A(_11212_), .B(_06760_), .Y(_06761_));
NAND_g _28409_ (.A(_06757_), .B(_06761_), .Y(_06762_));
NAND_g _28410_ (.A(_00012_[3]), .B(_06762_), .Y(_06763_));
NAND_g _28411_ (.A(_06753_), .B(_06763_), .Y(_06764_));
NAND_g _28412_ (.A(_11213_), .B(_06764_), .Y(_06765_));
AND_g _28413_ (.A(_06743_), .B(_06765_), .Y(_06766_));
NAND_g _28414_ (.A(_00012_[4]), .B(_06721_), .Y(_06767_));
NAND_g _28415_ (.A(_11216_), .B(_06766_), .Y(_06768_));
AND_g _28416_ (.A(_06767_), .B(_06768_), .Y(_06769_));
AND_g _28417_ (.A(_13561_), .B(_06769_), .Y(_06770_));
NAND_g _28418_ (.A(_05765_), .B(_06770_), .Y(_06771_));
AND_g _28419_ (.A(_06676_), .B(_06771_), .Y(_06772_));
AND_g _28420_ (.A(_06665_), .B(_06772_), .Y(_06773_));
NOR_g _28421_ (.A(_06663_), .B(_06773_), .Y(_01223_));
NOR_g _28422_ (.A(pcpi_rs1[17]), .B(_13425_), .Y(_06774_));
NAND_g _28423_ (.A(cpuregs_7[17]), .B(_00012_[2]), .Y(_06775_));
NAND_g _28424_ (.A(cpuregs_3[17]), .B(_11214_), .Y(_06776_));
NAND_g _28425_ (.A(_06775_), .B(_06776_), .Y(_06777_));
AND_g _28426_ (.A(_00012_[0]), .B(_06777_), .Y(_06778_));
NAND_g _28427_ (.A(cpuregs_6[17]), .B(_00012_[2]), .Y(_06779_));
NAND_g _28428_ (.A(cpuregs_2[17]), .B(_11214_), .Y(_06780_));
AND_g _28429_ (.A(_06779_), .B(_06780_), .Y(_06781_));
NOR_g _28430_ (.A(_00012_[0]), .B(_06781_), .Y(_06782_));
NOR_g _28431_ (.A(_06778_), .B(_06782_), .Y(_06783_));
NAND_g _28432_ (.A(cpuregs_5[17]), .B(_00012_[2]), .Y(_06784_));
NAND_g _28433_ (.A(cpuregs_1[17]), .B(_11214_), .Y(_06785_));
NAND_g _28434_ (.A(_06784_), .B(_06785_), .Y(_06786_));
NAND_g _28435_ (.A(_00012_[0]), .B(_06786_), .Y(_06787_));
NAND_g _28436_ (.A(cpuregs_4[17]), .B(_00012_[2]), .Y(_06788_));
NAND_g _28437_ (.A(cpuregs_0[17]), .B(_11214_), .Y(_06789_));
AND_g _28438_ (.A(_06788_), .B(_06789_), .Y(_06790_));
NOR_g _28439_ (.A(_00012_[0]), .B(_06790_), .Y(_06791_));
NAND_g _28440_ (.A(_00012_[1]), .B(_06783_), .Y(_06792_));
NOR_g _28441_ (.A(_00012_[1]), .B(_06791_), .Y(_06793_));
NAND_g _28442_ (.A(_06787_), .B(_06793_), .Y(_06794_));
AND_g _28443_ (.A(_06792_), .B(_06794_), .Y(_06795_));
NAND_g _28444_ (.A(_11215_), .B(_06795_), .Y(_06796_));
NAND_g _28445_ (.A(cpuregs_13[17]), .B(_00012_[0]), .Y(_06797_));
NAND_g _28446_ (.A(cpuregs_12[17]), .B(_11212_), .Y(_06798_));
AND_g _28447_ (.A(_00012_[2]), .B(_06798_), .Y(_06799_));
NAND_g _28448_ (.A(_06797_), .B(_06799_), .Y(_06800_));
NAND_g _28449_ (.A(cpuregs_9[17]), .B(_00012_[0]), .Y(_06801_));
NAND_g _28450_ (.A(cpuregs_8[17]), .B(_11212_), .Y(_06802_));
AND_g _28451_ (.A(_11214_), .B(_06802_), .Y(_06803_));
NAND_g _28452_ (.A(_06801_), .B(_06803_), .Y(_06804_));
AND_g _28453_ (.A(_11213_), .B(_06804_), .Y(_06805_));
NAND_g _28454_ (.A(_06800_), .B(_06805_), .Y(_06806_));
NAND_g _28455_ (.A(cpuregs_15[17]), .B(_00012_[0]), .Y(_06807_));
NAND_g _28456_ (.A(cpuregs_14[17]), .B(_11212_), .Y(_06808_));
AND_g _28457_ (.A(_00012_[2]), .B(_06808_), .Y(_06809_));
NAND_g _28458_ (.A(_06807_), .B(_06809_), .Y(_06810_));
NAND_g _28459_ (.A(cpuregs_11[17]), .B(_00012_[0]), .Y(_06811_));
NAND_g _28460_ (.A(cpuregs_10[17]), .B(_11212_), .Y(_06812_));
AND_g _28461_ (.A(_11214_), .B(_06812_), .Y(_06813_));
NAND_g _28462_ (.A(_06811_), .B(_06813_), .Y(_06814_));
AND_g _28463_ (.A(_00012_[1]), .B(_06814_), .Y(_06815_));
NAND_g _28464_ (.A(_06810_), .B(_06815_), .Y(_06816_));
NAND_g _28465_ (.A(_06806_), .B(_06816_), .Y(_06817_));
NAND_g _28466_ (.A(_00012_[3]), .B(_06817_), .Y(_06818_));
AND_g _28467_ (.A(_06796_), .B(_06818_), .Y(_06819_));
NAND_g _28468_ (.A(_11216_), .B(_06819_), .Y(_06820_));
NAND_g _28469_ (.A(_11017_), .B(_00012_[2]), .Y(_06821_));
NOR_g _28470_ (.A(cpuregs_18[17]), .B(_00012_[2]), .Y(_06822_));
NOR_g _28471_ (.A(_00012_[0]), .B(_06822_), .Y(_06823_));
NAND_g _28472_ (.A(_06821_), .B(_06823_), .Y(_06824_));
NAND_g _28473_ (.A(_11184_), .B(_00012_[2]), .Y(_06825_));
NOR_g _28474_ (.A(cpuregs_19[17]), .B(_00012_[2]), .Y(_06826_));
NOR_g _28475_ (.A(_11212_), .B(_06826_), .Y(_06827_));
NAND_g _28476_ (.A(_06825_), .B(_06827_), .Y(_06828_));
AND_g _28477_ (.A(_06824_), .B(_06828_), .Y(_06829_));
NAND_g _28478_ (.A(_11198_), .B(_00012_[2]), .Y(_06830_));
NOR_g _28479_ (.A(cpuregs_16[17]), .B(_00012_[2]), .Y(_06831_));
NOR_g _28480_ (.A(_00012_[0]), .B(_06831_), .Y(_06832_));
NAND_g _28481_ (.A(_06830_), .B(_06832_), .Y(_06833_));
NAND_g _28482_ (.A(_11031_), .B(_00012_[2]), .Y(_06834_));
NOR_g _28483_ (.A(cpuregs_17[17]), .B(_00012_[2]), .Y(_06835_));
NOR_g _28484_ (.A(_11212_), .B(_06835_), .Y(_06836_));
NAND_g _28485_ (.A(_06834_), .B(_06836_), .Y(_06837_));
AND_g _28486_ (.A(_06833_), .B(_06837_), .Y(_06838_));
NAND_g _28487_ (.A(_00012_[1]), .B(_06829_), .Y(_06839_));
NAND_g _28488_ (.A(_11213_), .B(_06838_), .Y(_06840_));
AND_g _28489_ (.A(_06839_), .B(_06840_), .Y(_06841_));
NAND_g _28490_ (.A(_11215_), .B(_06841_), .Y(_06842_));
NAND_g _28491_ (.A(cpuregs_29[17]), .B(_11213_), .Y(_06843_));
NAND_g _28492_ (.A(cpuregs_31[17]), .B(_00012_[1]), .Y(_06844_));
AND_g _28493_ (.A(_00012_[2]), .B(_06844_), .Y(_06845_));
NAND_g _28494_ (.A(_06843_), .B(_06845_), .Y(_06846_));
NAND_g _28495_ (.A(cpuregs_25[17]), .B(_11213_), .Y(_06847_));
NAND_g _28496_ (.A(cpuregs_27[17]), .B(_00012_[1]), .Y(_06848_));
AND_g _28497_ (.A(_11214_), .B(_06848_), .Y(_06849_));
NAND_g _28498_ (.A(_06847_), .B(_06849_), .Y(_06850_));
AND_g _28499_ (.A(_00012_[0]), .B(_06850_), .Y(_06851_));
NAND_g _28500_ (.A(_06846_), .B(_06851_), .Y(_06852_));
NAND_g _28501_ (.A(cpuregs_28[17]), .B(_11213_), .Y(_06853_));
NAND_g _28502_ (.A(cpuregs_30[17]), .B(_00012_[1]), .Y(_06854_));
AND_g _28503_ (.A(_00012_[2]), .B(_06854_), .Y(_06855_));
NAND_g _28504_ (.A(_06853_), .B(_06855_), .Y(_06856_));
NAND_g _28505_ (.A(cpuregs_24[17]), .B(_11213_), .Y(_06857_));
NAND_g _28506_ (.A(cpuregs_26[17]), .B(_00012_[1]), .Y(_06858_));
AND_g _28507_ (.A(_11214_), .B(_06858_), .Y(_06859_));
NAND_g _28508_ (.A(_06857_), .B(_06859_), .Y(_06860_));
AND_g _28509_ (.A(_11212_), .B(_06860_), .Y(_06861_));
NAND_g _28510_ (.A(_06856_), .B(_06861_), .Y(_06862_));
NAND_g _28511_ (.A(_06852_), .B(_06862_), .Y(_06863_));
NAND_g _28512_ (.A(_00012_[3]), .B(_06863_), .Y(_06864_));
AND_g _28513_ (.A(_06842_), .B(_06864_), .Y(_06865_));
NAND_g _28514_ (.A(_00012_[4]), .B(_06865_), .Y(_06866_));
AND_g _28515_ (.A(_13409_), .B(_06866_), .Y(_06867_));
AND_g _28516_ (.A(_06820_), .B(_06867_), .Y(_06868_));
AND_g _28517_ (.A(_13613_), .B(_06868_), .Y(_06869_));
NAND_g _28518_ (.A(reg_pc[17]), .B(_13714_), .Y(_06870_));
NAND_g _28519_ (.A(pcpi_rs1[21]), .B(_13419_), .Y(_06871_));
AND_g _28520_ (.A(_13383_), .B(_06540_), .Y(_06872_));
NAND_g _28521_ (.A(_06871_), .B(_06872_), .Y(_06873_));
NAND_g _28522_ (.A(pcpi_rs1[16]), .B(_13420_), .Y(_06874_));
AND_g _28523_ (.A(_13382_), .B(_06874_), .Y(_06875_));
NAND_g _28524_ (.A(_06537_), .B(_06875_), .Y(_06876_));
AND_g _28525_ (.A(_06873_), .B(_06876_), .Y(_06877_));
NAND_g _28526_ (.A(_13389_), .B(_06877_), .Y(_06878_));
AND_g _28527_ (.A(_06870_), .B(_06878_), .Y(_06879_));
NAND_g _28528_ (.A(_13425_), .B(_06879_), .Y(_06880_));
NOR_g _28529_ (.A(_06869_), .B(_06880_), .Y(_06881_));
XOR_g _28530_ (.A(decoded_imm[17]), .B(pcpi_rs1[17]), .Y(_06882_));
XNOR_g _28531_ (.A(_13524_), .B(_06882_), .Y(_06883_));
NAND_g _28532_ (.A(_13432_), .B(_06883_), .Y(_06884_));
AND_g _28533_ (.A(_06881_), .B(_06884_), .Y(_06885_));
NOR_g _28534_ (.A(_06774_), .B(_06885_), .Y(_01224_));
NOR_g _28535_ (.A(pcpi_rs1[18]), .B(_13425_), .Y(_06886_));
NAND_g _28536_ (.A(reg_pc[18]), .B(_13714_), .Y(_06887_));
NAND_g _28537_ (.A(pcpi_rs1[22]), .B(_13419_), .Y(_06888_));
AND_g _28538_ (.A(_13383_), .B(_06559_), .Y(_06889_));
NAND_g _28539_ (.A(_06888_), .B(_06889_), .Y(_06890_));
NAND_g _28540_ (.A(pcpi_rs1[17]), .B(_13420_), .Y(_06891_));
AND_g _28541_ (.A(_13382_), .B(_06891_), .Y(_06892_));
NAND_g _28542_ (.A(_06556_), .B(_06892_), .Y(_06893_));
AND_g _28543_ (.A(_06890_), .B(_06893_), .Y(_06894_));
NAND_g _28544_ (.A(_13389_), .B(_06894_), .Y(_06895_));
AND_g _28545_ (.A(_06887_), .B(_06895_), .Y(_06896_));
AND_g _28546_ (.A(_13425_), .B(_06896_), .Y(_06897_));
NAND_g _28547_ (.A(_11175_), .B(_00012_[2]), .Y(_06898_));
NOR_g _28548_ (.A(cpuregs_26[18]), .B(_00012_[2]), .Y(_06899_));
NOR_g _28549_ (.A(_00012_[0]), .B(_06899_), .Y(_06900_));
NAND_g _28550_ (.A(_06898_), .B(_06900_), .Y(_06901_));
NOR_g _28551_ (.A(cpuregs_27[18]), .B(_00012_[2]), .Y(_06902_));
NAND_g _28552_ (.A(_11091_), .B(_00012_[2]), .Y(_06903_));
NOR_g _28553_ (.A(_11212_), .B(_06902_), .Y(_06904_));
NAND_g _28554_ (.A(_06903_), .B(_06904_), .Y(_06905_));
NAND_g _28555_ (.A(_06901_), .B(_06905_), .Y(_06906_));
NAND_g _28556_ (.A(_00012_[3]), .B(_06906_), .Y(_06907_));
NAND_g _28557_ (.A(_11018_), .B(_00012_[2]), .Y(_06908_));
NOR_g _28558_ (.A(cpuregs_18[18]), .B(_00012_[2]), .Y(_06909_));
NOR_g _28559_ (.A(_00012_[0]), .B(_06909_), .Y(_06910_));
NAND_g _28560_ (.A(_06908_), .B(_06910_), .Y(_06911_));
NAND_g _28561_ (.A(_11185_), .B(_00012_[2]), .Y(_06912_));
NOR_g _28562_ (.A(cpuregs_19[18]), .B(_00012_[2]), .Y(_06913_));
NOR_g _28563_ (.A(_11212_), .B(_06913_), .Y(_06914_));
NAND_g _28564_ (.A(_06912_), .B(_06914_), .Y(_06915_));
NAND_g _28565_ (.A(_06911_), .B(_06915_), .Y(_06916_));
NAND_g _28566_ (.A(_11215_), .B(_06916_), .Y(_06917_));
NAND_g _28567_ (.A(_06907_), .B(_06917_), .Y(_06918_));
NAND_g _28568_ (.A(_00012_[1]), .B(_06918_), .Y(_06919_));
NAND_g _28569_ (.A(_11099_), .B(_00012_[2]), .Y(_06920_));
NOR_g _28570_ (.A(cpuregs_24[18]), .B(_00012_[2]), .Y(_06921_));
NOR_g _28571_ (.A(_00012_[0]), .B(_06921_), .Y(_06922_));
NAND_g _28572_ (.A(_06920_), .B(_06922_), .Y(_06923_));
NAND_g _28573_ (.A(_10931_), .B(_00012_[2]), .Y(_06924_));
NOR_g _28574_ (.A(cpuregs_25[18]), .B(_00012_[2]), .Y(_06925_));
NOR_g _28575_ (.A(_11212_), .B(_06925_), .Y(_06926_));
NAND_g _28576_ (.A(_06924_), .B(_06926_), .Y(_06927_));
NAND_g _28577_ (.A(_06923_), .B(_06927_), .Y(_06928_));
NAND_g _28578_ (.A(_00012_[3]), .B(_06928_), .Y(_06929_));
NAND_g _28579_ (.A(_11199_), .B(_00012_[2]), .Y(_06930_));
NOR_g _28580_ (.A(cpuregs_16[18]), .B(_00012_[2]), .Y(_06931_));
NOR_g _28581_ (.A(_00012_[0]), .B(_06931_), .Y(_06932_));
NAND_g _28582_ (.A(_06930_), .B(_06932_), .Y(_06933_));
NAND_g _28583_ (.A(_11032_), .B(_00012_[2]), .Y(_06934_));
NOR_g _28584_ (.A(cpuregs_17[18]), .B(_00012_[2]), .Y(_06935_));
NOR_g _28585_ (.A(_11212_), .B(_06935_), .Y(_06936_));
NAND_g _28586_ (.A(_06934_), .B(_06936_), .Y(_06937_));
NAND_g _28587_ (.A(_06933_), .B(_06937_), .Y(_06938_));
NAND_g _28588_ (.A(_11215_), .B(_06938_), .Y(_06939_));
NAND_g _28589_ (.A(_06929_), .B(_06939_), .Y(_06940_));
NAND_g _28590_ (.A(_11213_), .B(_06940_), .Y(_06941_));
NAND_g _28591_ (.A(_06919_), .B(_06941_), .Y(_06942_));
NAND_g _28592_ (.A(_00012_[4]), .B(_06942_), .Y(_06943_));
NAND_g _28593_ (.A(_10944_), .B(_00012_[2]), .Y(_06944_));
NOR_g _28594_ (.A(cpuregs_2[18]), .B(_00012_[2]), .Y(_06945_));
NOR_g _28595_ (.A(_00012_[0]), .B(_06945_), .Y(_06946_));
NAND_g _28596_ (.A(_06944_), .B(_06946_), .Y(_06947_));
NAND_g _28597_ (.A(_11130_), .B(_00012_[2]), .Y(_06948_));
NOR_g _28598_ (.A(cpuregs_3[18]), .B(_00012_[2]), .Y(_06949_));
NOR_g _28599_ (.A(_11212_), .B(_06949_), .Y(_06950_));
NAND_g _28600_ (.A(_06948_), .B(_06950_), .Y(_06951_));
NAND_g _28601_ (.A(_06947_), .B(_06951_), .Y(_06952_));
NAND_g _28602_ (.A(_11104_), .B(_00012_[2]), .Y(_06953_));
NOR_g _28603_ (.A(cpuregs_10[18]), .B(_00012_[2]), .Y(_06954_));
NOR_g _28604_ (.A(_00012_[0]), .B(_06954_), .Y(_06955_));
AND_g _28605_ (.A(_06953_), .B(_06955_), .Y(_06956_));
NOR_g _28606_ (.A(cpuregs_11[18]), .B(_00012_[2]), .Y(_06957_));
NAND_g _28607_ (.A(_11166_), .B(_00012_[2]), .Y(_06958_));
NOR_g _28608_ (.A(_11212_), .B(_06957_), .Y(_06959_));
AND_g _28609_ (.A(_06958_), .B(_06959_), .Y(_06960_));
NOR_g _28610_ (.A(_06956_), .B(_06960_), .Y(_06961_));
NOR_g _28611_ (.A(_00012_[3]), .B(_06952_), .Y(_06962_));
AND_g _28612_ (.A(_00012_[3]), .B(_06961_), .Y(_06963_));
NOR_g _28613_ (.A(_06962_), .B(_06963_), .Y(_06964_));
NAND_g _28614_ (.A(_00012_[1]), .B(_06964_), .Y(_06965_));
NAND_g _28615_ (.A(_11120_), .B(_00012_[2]), .Y(_06966_));
NOR_g _28616_ (.A(cpuregs_8[18]), .B(_00012_[2]), .Y(_06967_));
NOR_g _28617_ (.A(_00012_[0]), .B(_06967_), .Y(_06968_));
AND_g _28618_ (.A(_06966_), .B(_06968_), .Y(_06969_));
NOR_g _28619_ (.A(cpuregs_9[18]), .B(_00012_[2]), .Y(_06970_));
NAND_g _28620_ (.A(_11150_), .B(_00012_[2]), .Y(_06971_));
NOR_g _28621_ (.A(_11212_), .B(_06970_), .Y(_06972_));
AND_g _28622_ (.A(_06971_), .B(_06972_), .Y(_06973_));
NOR_g _28623_ (.A(_06969_), .B(_06973_), .Y(_06974_));
NAND_g _28624_ (.A(_10956_), .B(_00012_[2]), .Y(_06975_));
NOR_g _28625_ (.A(cpuregs_0[18]), .B(_00012_[2]), .Y(_06976_));
NOR_g _28626_ (.A(_00012_[0]), .B(_06976_), .Y(_06977_));
NAND_g _28627_ (.A(_06975_), .B(_06977_), .Y(_06978_));
NAND_g _28628_ (.A(_11114_), .B(_00012_[2]), .Y(_06979_));
NOR_g _28629_ (.A(cpuregs_1[18]), .B(_00012_[2]), .Y(_06980_));
NOR_g _28630_ (.A(_11212_), .B(_06980_), .Y(_06981_));
NAND_g _28631_ (.A(_06979_), .B(_06981_), .Y(_06982_));
NAND_g _28632_ (.A(_06978_), .B(_06982_), .Y(_06983_));
NOR_g _28633_ (.A(_00012_[3]), .B(_06983_), .Y(_06984_));
AND_g _28634_ (.A(_00012_[3]), .B(_06974_), .Y(_06985_));
NOR_g _28635_ (.A(_06984_), .B(_06985_), .Y(_06986_));
NAND_g _28636_ (.A(_11213_), .B(_06986_), .Y(_06987_));
NAND_g _28637_ (.A(_06965_), .B(_06987_), .Y(_06988_));
NAND_g _28638_ (.A(_11216_), .B(_06988_), .Y(_06989_));
NAND_g _28639_ (.A(_06943_), .B(_06989_), .Y(_06990_));
AND_g _28640_ (.A(_13561_), .B(_06990_), .Y(_06991_));
NAND_g _28641_ (.A(_05765_), .B(_06991_), .Y(_06992_));
AND_g _28642_ (.A(_06897_), .B(_06992_), .Y(_06993_));
XOR_g _28643_ (.A(_13457_), .B(_13526_), .Y(_06994_));
NAND_g _28644_ (.A(_13432_), .B(_06994_), .Y(_06995_));
AND_g _28645_ (.A(_06993_), .B(_06995_), .Y(_06996_));
NOR_g _28646_ (.A(_06886_), .B(_06996_), .Y(_01225_));
NOR_g _28647_ (.A(pcpi_rs1[19]), .B(_13425_), .Y(_06997_));
XOR_g _28648_ (.A(decoded_imm[19]), .B(pcpi_rs1[19]), .Y(_06998_));
XNOR_g _28649_ (.A(_13528_), .B(_06998_), .Y(_06999_));
NAND_g _28650_ (.A(_13432_), .B(_06999_), .Y(_07000_));
NOR_g _28651_ (.A(cpuregs_11[19]), .B(_00012_[2]), .Y(_07001_));
AND_g _28652_ (.A(_11167_), .B(_00012_[2]), .Y(_07002_));
NOR_g _28653_ (.A(_07001_), .B(_07002_), .Y(_07003_));
NOR_g _28654_ (.A(_11212_), .B(_07003_), .Y(_07004_));
NOR_g _28655_ (.A(cpuregs_10[19]), .B(_00012_[2]), .Y(_07005_));
AND_g _28656_ (.A(_11105_), .B(_00012_[2]), .Y(_07006_));
NOR_g _28657_ (.A(_07005_), .B(_07006_), .Y(_07007_));
NOR_g _28658_ (.A(_00012_[0]), .B(_07007_), .Y(_07008_));
NOR_g _28659_ (.A(_07004_), .B(_07008_), .Y(_07009_));
NAND_g _28660_ (.A(cpuregs_6[19]), .B(_00012_[2]), .Y(_07010_));
NAND_g _28661_ (.A(cpuregs_2[19]), .B(_11214_), .Y(_07011_));
AND_g _28662_ (.A(_07010_), .B(_07011_), .Y(_07012_));
NAND_g _28663_ (.A(_11212_), .B(_07012_), .Y(_07013_));
NAND_g _28664_ (.A(cpuregs_7[19]), .B(_00012_[2]), .Y(_07014_));
NAND_g _28665_ (.A(cpuregs_3[19]), .B(_11214_), .Y(_07015_));
AND_g _28666_ (.A(_00012_[0]), .B(_07015_), .Y(_07016_));
NAND_g _28667_ (.A(_07014_), .B(_07016_), .Y(_07017_));
AND_g _28668_ (.A(_11215_), .B(_07017_), .Y(_07018_));
NAND_g _28669_ (.A(_07013_), .B(_07018_), .Y(_07019_));
NAND_g _28670_ (.A(_00012_[3]), .B(_07009_), .Y(_07020_));
AND_g _28671_ (.A(_07019_), .B(_07020_), .Y(_07021_));
NAND_g _28672_ (.A(_00012_[1]), .B(_07021_), .Y(_07022_));
NOR_g _28673_ (.A(cpuregs_8[19]), .B(_00012_[2]), .Y(_07023_));
AND_g _28674_ (.A(_11121_), .B(_00012_[2]), .Y(_07024_));
NOR_g _28675_ (.A(_07023_), .B(_07024_), .Y(_07025_));
NOR_g _28676_ (.A(cpuregs_9[19]), .B(_00012_[2]), .Y(_07026_));
NAND_g _28677_ (.A(_11151_), .B(_00012_[2]), .Y(_07027_));
NAND_g _28678_ (.A(_11212_), .B(_07025_), .Y(_07028_));
NOR_g _28679_ (.A(_11212_), .B(_07026_), .Y(_07029_));
NAND_g _28680_ (.A(_07027_), .B(_07029_), .Y(_07030_));
AND_g _28681_ (.A(_00012_[3]), .B(_07030_), .Y(_07031_));
NAND_g _28682_ (.A(_07028_), .B(_07031_), .Y(_07032_));
NAND_g _28683_ (.A(cpuregs_1[19]), .B(_11214_), .Y(_07033_));
NAND_g _28684_ (.A(cpuregs_5[19]), .B(_00012_[2]), .Y(_07034_));
AND_g _28685_ (.A(_00012_[0]), .B(_07034_), .Y(_07035_));
NAND_g _28686_ (.A(_07033_), .B(_07035_), .Y(_07036_));
NAND_g _28687_ (.A(cpuregs_4[19]), .B(_00012_[2]), .Y(_07037_));
NAND_g _28688_ (.A(cpuregs_0[19]), .B(_11214_), .Y(_07038_));
AND_g _28689_ (.A(_11212_), .B(_07038_), .Y(_07039_));
NAND_g _28690_ (.A(_07037_), .B(_07039_), .Y(_07040_));
NAND_g _28691_ (.A(_07036_), .B(_07040_), .Y(_07041_));
NAND_g _28692_ (.A(_11215_), .B(_07041_), .Y(_07042_));
NAND_g _28693_ (.A(_07032_), .B(_07042_), .Y(_07043_));
NAND_g _28694_ (.A(_11213_), .B(_07043_), .Y(_07044_));
NAND_g _28695_ (.A(_07022_), .B(_07044_), .Y(_07045_));
NAND_g _28696_ (.A(_11216_), .B(_07045_), .Y(_07046_));
NAND_g _28697_ (.A(cpuregs_18[19]), .B(_11214_), .Y(_07047_));
NAND_g _28698_ (.A(cpuregs_22[19]), .B(_00012_[2]), .Y(_07048_));
AND_g _28699_ (.A(_11212_), .B(_07048_), .Y(_07049_));
NAND_g _28700_ (.A(_07047_), .B(_07049_), .Y(_07050_));
NAND_g _28701_ (.A(cpuregs_19[19]), .B(_11214_), .Y(_07051_));
NAND_g _28702_ (.A(cpuregs_23[19]), .B(_00012_[2]), .Y(_07052_));
AND_g _28703_ (.A(_00012_[0]), .B(_07052_), .Y(_07053_));
NAND_g _28704_ (.A(_07051_), .B(_07053_), .Y(_07054_));
NAND_g _28705_ (.A(_07050_), .B(_07054_), .Y(_07055_));
NAND_g _28706_ (.A(_11215_), .B(_07055_), .Y(_07056_));
NAND_g _28707_ (.A(cpuregs_26[19]), .B(_11214_), .Y(_07057_));
NAND_g _28708_ (.A(cpuregs_30[19]), .B(_00012_[2]), .Y(_07058_));
AND_g _28709_ (.A(_11212_), .B(_07058_), .Y(_07059_));
NAND_g _28710_ (.A(_07057_), .B(_07059_), .Y(_07060_));
NAND_g _28711_ (.A(cpuregs_27[19]), .B(_11214_), .Y(_07061_));
NAND_g _28712_ (.A(cpuregs_31[19]), .B(_00012_[2]), .Y(_07062_));
AND_g _28713_ (.A(_00012_[0]), .B(_07062_), .Y(_07063_));
NAND_g _28714_ (.A(_07061_), .B(_07063_), .Y(_07064_));
NAND_g _28715_ (.A(_07060_), .B(_07064_), .Y(_07065_));
NAND_g _28716_ (.A(_00012_[3]), .B(_07065_), .Y(_07066_));
NAND_g _28717_ (.A(_07056_), .B(_07066_), .Y(_07067_));
NAND_g _28718_ (.A(_00012_[1]), .B(_07067_), .Y(_07068_));
NAND_g _28719_ (.A(cpuregs_24[19]), .B(_11214_), .Y(_07069_));
NAND_g _28720_ (.A(cpuregs_28[19]), .B(_00012_[2]), .Y(_07070_));
AND_g _28721_ (.A(_11212_), .B(_07070_), .Y(_07071_));
NAND_g _28722_ (.A(_07069_), .B(_07071_), .Y(_07072_));
NAND_g _28723_ (.A(cpuregs_25[19]), .B(_11214_), .Y(_07073_));
NAND_g _28724_ (.A(cpuregs_29[19]), .B(_00012_[2]), .Y(_07074_));
AND_g _28725_ (.A(_00012_[0]), .B(_07074_), .Y(_07075_));
NAND_g _28726_ (.A(_07073_), .B(_07075_), .Y(_07076_));
NAND_g _28727_ (.A(_07072_), .B(_07076_), .Y(_07077_));
NAND_g _28728_ (.A(_00012_[3]), .B(_07077_), .Y(_07078_));
NAND_g _28729_ (.A(cpuregs_20[19]), .B(_00012_[2]), .Y(_07079_));
NAND_g _28730_ (.A(cpuregs_16[19]), .B(_11214_), .Y(_07080_));
AND_g _28731_ (.A(_11212_), .B(_07080_), .Y(_07081_));
NAND_g _28732_ (.A(_07079_), .B(_07081_), .Y(_07082_));
NAND_g _28733_ (.A(cpuregs_21[19]), .B(_00012_[2]), .Y(_07083_));
NAND_g _28734_ (.A(cpuregs_17[19]), .B(_11214_), .Y(_07084_));
AND_g _28735_ (.A(_00012_[0]), .B(_07084_), .Y(_07085_));
NAND_g _28736_ (.A(_07083_), .B(_07085_), .Y(_07086_));
NAND_g _28737_ (.A(_07082_), .B(_07086_), .Y(_07087_));
NAND_g _28738_ (.A(_11215_), .B(_07087_), .Y(_07088_));
NAND_g _28739_ (.A(_07078_), .B(_07088_), .Y(_07089_));
NAND_g _28740_ (.A(_11213_), .B(_07089_), .Y(_07090_));
NAND_g _28741_ (.A(_07068_), .B(_07090_), .Y(_07091_));
NAND_g _28742_ (.A(_00012_[4]), .B(_07091_), .Y(_07092_));
AND_g _28743_ (.A(_07046_), .B(_07092_), .Y(_07093_));
AND_g _28744_ (.A(_13613_), .B(_07093_), .Y(_07094_));
NAND_g _28745_ (.A(_13409_), .B(_07094_), .Y(_07095_));
NAND_g _28746_ (.A(reg_pc[19]), .B(_13714_), .Y(_07096_));
NAND_g _28747_ (.A(pcpi_rs1[18]), .B(_13420_), .Y(_07097_));
AND_g _28748_ (.A(_06670_), .B(_07097_), .Y(_07098_));
NAND_g _28749_ (.A(_13382_), .B(_07098_), .Y(_07099_));
NAND_g _28750_ (.A(pcpi_rs1[23]), .B(_13419_), .Y(_07100_));
AND_g _28751_ (.A(_06667_), .B(_07100_), .Y(_07101_));
NAND_g _28752_ (.A(_13383_), .B(_07101_), .Y(_07102_));
AND_g _28753_ (.A(_07099_), .B(_07102_), .Y(_07103_));
NAND_g _28754_ (.A(_13389_), .B(_07103_), .Y(_07104_));
AND_g _28755_ (.A(_07096_), .B(_07104_), .Y(_07105_));
AND_g _28756_ (.A(_13425_), .B(_07105_), .Y(_07106_));
AND_g _28757_ (.A(_07095_), .B(_07106_), .Y(_07107_));
AND_g _28758_ (.A(_07000_), .B(_07107_), .Y(_07108_));
NOR_g _28759_ (.A(_06997_), .B(_07108_), .Y(_01226_));
NOR_g _28760_ (.A(pcpi_rs1[20]), .B(_13425_), .Y(_07109_));
NAND_g _28761_ (.A(reg_pc[20]), .B(_13714_), .Y(_07110_));
NAND_g _28762_ (.A(pcpi_rs1[24]), .B(_13419_), .Y(_07111_));
AND_g _28763_ (.A(_13383_), .B(_06874_), .Y(_07112_));
NAND_g _28764_ (.A(_07111_), .B(_07112_), .Y(_07113_));
NAND_g _28765_ (.A(pcpi_rs1[19]), .B(_13420_), .Y(_07114_));
AND_g _28766_ (.A(_13382_), .B(_07114_), .Y(_07115_));
NAND_g _28767_ (.A(_06871_), .B(_07115_), .Y(_07116_));
AND_g _28768_ (.A(_07113_), .B(_07116_), .Y(_07117_));
NAND_g _28769_ (.A(_13389_), .B(_07117_), .Y(_07118_));
AND_g _28770_ (.A(_07110_), .B(_07118_), .Y(_07119_));
AND_g _28771_ (.A(_13425_), .B(_07119_), .Y(_07120_));
NAND_g _28772_ (.A(_11176_), .B(_00012_[2]), .Y(_07121_));
NOR_g _28773_ (.A(cpuregs_26[20]), .B(_00012_[2]), .Y(_07122_));
NOR_g _28774_ (.A(_00012_[0]), .B(_07122_), .Y(_07123_));
AND_g _28775_ (.A(_07121_), .B(_07123_), .Y(_07124_));
NOR_g _28776_ (.A(cpuregs_27[20]), .B(_00012_[2]), .Y(_07125_));
NAND_g _28777_ (.A(_11092_), .B(_00012_[2]), .Y(_07126_));
NOR_g _28778_ (.A(_11212_), .B(_07125_), .Y(_07127_));
AND_g _28779_ (.A(_07126_), .B(_07127_), .Y(_07128_));
NOR_g _28780_ (.A(_07124_), .B(_07128_), .Y(_07129_));
NAND_g _28781_ (.A(cpuregs_22[20]), .B(_00012_[2]), .Y(_07130_));
NAND_g _28782_ (.A(cpuregs_18[20]), .B(_11214_), .Y(_07131_));
AND_g _28783_ (.A(_11212_), .B(_07131_), .Y(_07132_));
NAND_g _28784_ (.A(_07130_), .B(_07132_), .Y(_07133_));
NAND_g _28785_ (.A(cpuregs_19[20]), .B(_11214_), .Y(_07134_));
NAND_g _28786_ (.A(cpuregs_23[20]), .B(_00012_[2]), .Y(_07135_));
AND_g _28787_ (.A(_00012_[0]), .B(_07135_), .Y(_07136_));
NAND_g _28788_ (.A(_07134_), .B(_07136_), .Y(_07137_));
NAND_g _28789_ (.A(_07133_), .B(_07137_), .Y(_07138_));
NAND_g _28790_ (.A(_11215_), .B(_07138_), .Y(_07139_));
NAND_g _28791_ (.A(_00012_[3]), .B(_07129_), .Y(_07140_));
AND_g _28792_ (.A(_07139_), .B(_07140_), .Y(_07141_));
NAND_g _28793_ (.A(_00012_[4]), .B(_07141_), .Y(_07142_));
NAND_g _28794_ (.A(cpuregs_6[20]), .B(_00012_[2]), .Y(_07143_));
NAND_g _28795_ (.A(cpuregs_2[20]), .B(_11214_), .Y(_07144_));
AND_g _28796_ (.A(_11212_), .B(_07144_), .Y(_07145_));
NAND_g _28797_ (.A(_07143_), .B(_07145_), .Y(_07146_));
NAND_g _28798_ (.A(cpuregs_3[20]), .B(_11214_), .Y(_07147_));
NAND_g _28799_ (.A(cpuregs_7[20]), .B(_00012_[2]), .Y(_07148_));
AND_g _28800_ (.A(_00012_[0]), .B(_07148_), .Y(_07149_));
NAND_g _28801_ (.A(_07147_), .B(_07149_), .Y(_07150_));
NOR_g _28802_ (.A(cpuregs_11[20]), .B(_00012_[2]), .Y(_07151_));
NAND_g _28803_ (.A(_11168_), .B(_00012_[2]), .Y(_07152_));
NOR_g _28804_ (.A(cpuregs_10[20]), .B(_00012_[2]), .Y(_07153_));
NOR_g _28805_ (.A(cpuregs_14[20]), .B(_11214_), .Y(_07154_));
NOR_g _28806_ (.A(_07153_), .B(_07154_), .Y(_07155_));
NAND_g _28807_ (.A(_07146_), .B(_07150_), .Y(_07156_));
NAND_g _28808_ (.A(_11215_), .B(_07156_), .Y(_07157_));
NAND_g _28809_ (.A(_11212_), .B(_07155_), .Y(_07158_));
NOR_g _28810_ (.A(_11212_), .B(_07151_), .Y(_07159_));
NAND_g _28811_ (.A(_07152_), .B(_07159_), .Y(_07160_));
AND_g _28812_ (.A(_00012_[3]), .B(_07160_), .Y(_07161_));
NAND_g _28813_ (.A(_07158_), .B(_07161_), .Y(_07162_));
AND_g _28814_ (.A(_07157_), .B(_07162_), .Y(_07163_));
NAND_g _28815_ (.A(_11216_), .B(_07163_), .Y(_07164_));
NAND_g _28816_ (.A(_07142_), .B(_07164_), .Y(_07165_));
NAND_g _28817_ (.A(_00012_[1]), .B(_07165_), .Y(_07166_));
NAND_g _28818_ (.A(_11100_), .B(_00012_[2]), .Y(_07167_));
NOR_g _28819_ (.A(cpuregs_24[20]), .B(_00012_[2]), .Y(_07168_));
NOR_g _28820_ (.A(_00012_[0]), .B(_07168_), .Y(_07169_));
NAND_g _28821_ (.A(_07167_), .B(_07169_), .Y(_07170_));
NAND_g _28822_ (.A(_10932_), .B(_00012_[2]), .Y(_07171_));
NOR_g _28823_ (.A(cpuregs_25[20]), .B(_00012_[2]), .Y(_07172_));
NOR_g _28824_ (.A(_11212_), .B(_07172_), .Y(_07173_));
NAND_g _28825_ (.A(_07171_), .B(_07173_), .Y(_07174_));
NAND_g _28826_ (.A(_07170_), .B(_07174_), .Y(_07175_));
NAND_g _28827_ (.A(_00012_[3]), .B(_07175_), .Y(_07176_));
NAND_g _28828_ (.A(cpuregs_20[20]), .B(_00012_[2]), .Y(_07177_));
NAND_g _28829_ (.A(cpuregs_16[20]), .B(_11214_), .Y(_07178_));
AND_g _28830_ (.A(_07177_), .B(_07178_), .Y(_07179_));
NAND_g _28831_ (.A(_11212_), .B(_07179_), .Y(_07180_));
NAND_g _28832_ (.A(cpuregs_21[20]), .B(_00012_[2]), .Y(_07181_));
NAND_g _28833_ (.A(cpuregs_17[20]), .B(_11214_), .Y(_07182_));
AND_g _28834_ (.A(_00012_[0]), .B(_07182_), .Y(_07183_));
NAND_g _28835_ (.A(_07181_), .B(_07183_), .Y(_07184_));
AND_g _28836_ (.A(_11215_), .B(_07184_), .Y(_07185_));
NAND_g _28837_ (.A(_07180_), .B(_07185_), .Y(_07186_));
NAND_g _28838_ (.A(_07176_), .B(_07186_), .Y(_07187_));
NAND_g _28839_ (.A(_00012_[4]), .B(_07187_), .Y(_07188_));
NAND_g _28840_ (.A(cpuregs_4[20]), .B(_00012_[2]), .Y(_07189_));
NAND_g _28841_ (.A(cpuregs_0[20]), .B(_11214_), .Y(_07190_));
AND_g _28842_ (.A(_07189_), .B(_07190_), .Y(_07191_));
NAND_g _28843_ (.A(_11212_), .B(_07191_), .Y(_07192_));
NAND_g _28844_ (.A(cpuregs_5[20]), .B(_00012_[2]), .Y(_07193_));
NAND_g _28845_ (.A(cpuregs_1[20]), .B(_11214_), .Y(_07194_));
AND_g _28846_ (.A(_00012_[0]), .B(_07194_), .Y(_07195_));
NAND_g _28847_ (.A(_07193_), .B(_07195_), .Y(_07196_));
AND_g _28848_ (.A(_11215_), .B(_07196_), .Y(_07197_));
NAND_g _28849_ (.A(_07192_), .B(_07197_), .Y(_07198_));
NOR_g _28850_ (.A(cpuregs_8[20]), .B(_00012_[2]), .Y(_07199_));
NOR_g _28851_ (.A(cpuregs_12[20]), .B(_11214_), .Y(_07200_));
NOR_g _28852_ (.A(_07199_), .B(_07200_), .Y(_07201_));
NOR_g _28853_ (.A(cpuregs_9[20]), .B(_00012_[2]), .Y(_07202_));
NOT_g _28854_ (.A(_07202_), .Y(_07203_));
NAND_g _28855_ (.A(_11152_), .B(_00012_[2]), .Y(_07204_));
AND_g _28856_ (.A(_00012_[0]), .B(_07204_), .Y(_07205_));
NAND_g _28857_ (.A(_07203_), .B(_07205_), .Y(_07206_));
NAND_g _28858_ (.A(_11212_), .B(_07201_), .Y(_07207_));
NAND_g _28859_ (.A(_07206_), .B(_07207_), .Y(_07208_));
NAND_g _28860_ (.A(_00012_[3]), .B(_07208_), .Y(_07209_));
NAND_g _28861_ (.A(_07198_), .B(_07209_), .Y(_07210_));
NAND_g _28862_ (.A(_11216_), .B(_07210_), .Y(_07211_));
NAND_g _28863_ (.A(_07188_), .B(_07211_), .Y(_07212_));
NAND_g _28864_ (.A(_11213_), .B(_07212_), .Y(_07213_));
NAND_g _28865_ (.A(_07166_), .B(_07213_), .Y(_07214_));
AND_g _28866_ (.A(_13561_), .B(_07214_), .Y(_07215_));
NAND_g _28867_ (.A(_05765_), .B(_07215_), .Y(_07216_));
AND_g _28868_ (.A(_07120_), .B(_07216_), .Y(_07217_));
XOR_g _28869_ (.A(_13453_), .B(_13530_), .Y(_07218_));
NAND_g _28870_ (.A(_13432_), .B(_07218_), .Y(_07219_));
AND_g _28871_ (.A(_07217_), .B(_07219_), .Y(_07220_));
NOR_g _28872_ (.A(_07109_), .B(_07220_), .Y(_01227_));
NOR_g _28873_ (.A(pcpi_rs1[21]), .B(_13425_), .Y(_07221_));
XOR_g _28874_ (.A(decoded_imm[21]), .B(pcpi_rs1[21]), .Y(_07222_));
XNOR_g _28875_ (.A(_13532_), .B(_07222_), .Y(_07223_));
NAND_g _28876_ (.A(_13432_), .B(_07223_), .Y(_07224_));
NAND_g _28877_ (.A(reg_pc[21]), .B(_13714_), .Y(_07225_));
NAND_g _28878_ (.A(pcpi_rs1[20]), .B(_13420_), .Y(_07226_));
AND_g _28879_ (.A(_06888_), .B(_07226_), .Y(_07227_));
NAND_g _28880_ (.A(_13382_), .B(_07227_), .Y(_07228_));
NAND_g _28881_ (.A(pcpi_rs1[25]), .B(_13419_), .Y(_07229_));
AND_g _28882_ (.A(_06891_), .B(_07229_), .Y(_07230_));
NAND_g _28883_ (.A(_13383_), .B(_07230_), .Y(_07231_));
NOR_g _28884_ (.A(cpuregs_16[21]), .B(_00012_[2]), .Y(_07232_));
AND_g _28885_ (.A(_11200_), .B(_00012_[2]), .Y(_07233_));
NOR_g _28886_ (.A(_07232_), .B(_07233_), .Y(_07234_));
NOR_g _28887_ (.A(cpuregs_18[21]), .B(_00012_[2]), .Y(_07235_));
AND_g _28888_ (.A(_11019_), .B(_00012_[2]), .Y(_07236_));
NOR_g _28889_ (.A(_07235_), .B(_07236_), .Y(_07237_));
NOR_g _28890_ (.A(cpuregs_17[21]), .B(_00012_[2]), .Y(_07238_));
NAND_g _28891_ (.A(_11033_), .B(_00012_[2]), .Y(_07239_));
NAND_g _28892_ (.A(_11186_), .B(_00012_[2]), .Y(_07240_));
NOR_g _28893_ (.A(cpuregs_19[21]), .B(_00012_[2]), .Y(_07241_));
NOR_g _28894_ (.A(_11212_), .B(_07241_), .Y(_07242_));
NAND_g _28895_ (.A(_07240_), .B(_07242_), .Y(_07243_));
NAND_g _28896_ (.A(_11212_), .B(_07237_), .Y(_07244_));
AND_g _28897_ (.A(_07243_), .B(_07244_), .Y(_07245_));
NAND_g _28898_ (.A(_00012_[1]), .B(_07245_), .Y(_07246_));
NOR_g _28899_ (.A(_11212_), .B(_07238_), .Y(_07247_));
NAND_g _28900_ (.A(_07239_), .B(_07247_), .Y(_07248_));
NAND_g _28901_ (.A(_11212_), .B(_07234_), .Y(_07249_));
AND_g _28902_ (.A(_07248_), .B(_07249_), .Y(_07250_));
NAND_g _28903_ (.A(_11213_), .B(_07250_), .Y(_07251_));
AND_g _28904_ (.A(_07246_), .B(_07251_), .Y(_07252_));
NAND_g _28905_ (.A(_11215_), .B(_07252_), .Y(_07253_));
NAND_g _28906_ (.A(cpuregs_27[21]), .B(_00012_[1]), .Y(_07254_));
NAND_g _28907_ (.A(cpuregs_25[21]), .B(_11213_), .Y(_07255_));
NAND_g _28908_ (.A(_07254_), .B(_07255_), .Y(_07256_));
NAND_g _28909_ (.A(_11214_), .B(_07256_), .Y(_07257_));
NAND_g _28910_ (.A(cpuregs_31[21]), .B(_00012_[1]), .Y(_07258_));
NAND_g _28911_ (.A(cpuregs_29[21]), .B(_11213_), .Y(_07259_));
NAND_g _28912_ (.A(_07258_), .B(_07259_), .Y(_07260_));
NAND_g _28913_ (.A(_00012_[2]), .B(_07260_), .Y(_07261_));
AND_g _28914_ (.A(_00012_[0]), .B(_07261_), .Y(_07262_));
NAND_g _28915_ (.A(_07257_), .B(_07262_), .Y(_07263_));
NAND_g _28916_ (.A(cpuregs_26[21]), .B(_00012_[1]), .Y(_07264_));
NAND_g _28917_ (.A(cpuregs_24[21]), .B(_11213_), .Y(_07265_));
NAND_g _28918_ (.A(_07264_), .B(_07265_), .Y(_07266_));
NAND_g _28919_ (.A(_11214_), .B(_07266_), .Y(_07267_));
NAND_g _28920_ (.A(cpuregs_30[21]), .B(_00012_[1]), .Y(_07268_));
NAND_g _28921_ (.A(cpuregs_28[21]), .B(_11213_), .Y(_07269_));
NAND_g _28922_ (.A(_07268_), .B(_07269_), .Y(_07270_));
NAND_g _28923_ (.A(_00012_[2]), .B(_07270_), .Y(_07271_));
AND_g _28924_ (.A(_11212_), .B(_07271_), .Y(_07272_));
NAND_g _28925_ (.A(_07267_), .B(_07272_), .Y(_07273_));
AND_g _28926_ (.A(_00012_[3]), .B(_07273_), .Y(_07274_));
NAND_g _28927_ (.A(_07263_), .B(_07274_), .Y(_07275_));
AND_g _28928_ (.A(_07253_), .B(_07275_), .Y(_07276_));
NAND_g _28929_ (.A(cpuregs_1[21]), .B(_11214_), .Y(_07277_));
NAND_g _28930_ (.A(cpuregs_5[21]), .B(_00012_[2]), .Y(_07278_));
AND_g _28931_ (.A(_00012_[0]), .B(_07278_), .Y(_07279_));
NAND_g _28932_ (.A(_07277_), .B(_07279_), .Y(_07280_));
NAND_g _28933_ (.A(cpuregs_0[21]), .B(_11214_), .Y(_07281_));
NAND_g _28934_ (.A(cpuregs_4[21]), .B(_00012_[2]), .Y(_07282_));
AND_g _28935_ (.A(_11212_), .B(_07282_), .Y(_07283_));
NAND_g _28936_ (.A(_07281_), .B(_07283_), .Y(_07284_));
AND_g _28937_ (.A(_11213_), .B(_07284_), .Y(_07285_));
NAND_g _28938_ (.A(_07280_), .B(_07285_), .Y(_07286_));
NAND_g _28939_ (.A(cpuregs_3[21]), .B(_11214_), .Y(_07287_));
NAND_g _28940_ (.A(cpuregs_7[21]), .B(_00012_[2]), .Y(_07288_));
AND_g _28941_ (.A(_00012_[0]), .B(_07288_), .Y(_07289_));
NAND_g _28942_ (.A(_07287_), .B(_07289_), .Y(_07290_));
NAND_g _28943_ (.A(cpuregs_2[21]), .B(_11214_), .Y(_07291_));
NAND_g _28944_ (.A(cpuregs_6[21]), .B(_00012_[2]), .Y(_07292_));
AND_g _28945_ (.A(_11212_), .B(_07292_), .Y(_07293_));
NAND_g _28946_ (.A(_07291_), .B(_07293_), .Y(_07294_));
AND_g _28947_ (.A(_00012_[1]), .B(_07294_), .Y(_07295_));
NAND_g _28948_ (.A(_07290_), .B(_07295_), .Y(_07296_));
NAND_g _28949_ (.A(_07286_), .B(_07296_), .Y(_07297_));
NAND_g _28950_ (.A(_11215_), .B(_07297_), .Y(_07298_));
NAND_g _28951_ (.A(cpuregs_14[21]), .B(_11212_), .Y(_07299_));
NAND_g _28952_ (.A(cpuregs_15[21]), .B(_00012_[0]), .Y(_07300_));
NAND_g _28953_ (.A(_07299_), .B(_07300_), .Y(_07301_));
NAND_g _28954_ (.A(_00012_[2]), .B(_07301_), .Y(_07302_));
NAND_g _28955_ (.A(cpuregs_10[21]), .B(_11212_), .Y(_07303_));
NAND_g _28956_ (.A(cpuregs_11[21]), .B(_00012_[0]), .Y(_07304_));
NAND_g _28957_ (.A(_07303_), .B(_07304_), .Y(_07305_));
NAND_g _28958_ (.A(_11214_), .B(_07305_), .Y(_07306_));
AND_g _28959_ (.A(_07302_), .B(_07306_), .Y(_07307_));
NAND_g _28960_ (.A(cpuregs_12[21]), .B(_11212_), .Y(_07308_));
NAND_g _28961_ (.A(cpuregs_13[21]), .B(_00012_[0]), .Y(_07309_));
NAND_g _28962_ (.A(_07308_), .B(_07309_), .Y(_07310_));
NAND_g _28963_ (.A(_00012_[2]), .B(_07310_), .Y(_07311_));
NAND_g _28964_ (.A(cpuregs_8[21]), .B(_11212_), .Y(_07312_));
NAND_g _28965_ (.A(cpuregs_9[21]), .B(_00012_[0]), .Y(_07313_));
NAND_g _28966_ (.A(_07312_), .B(_07313_), .Y(_07314_));
NAND_g _28967_ (.A(_11214_), .B(_07314_), .Y(_07315_));
AND_g _28968_ (.A(_07311_), .B(_07315_), .Y(_07316_));
NAND_g _28969_ (.A(_11213_), .B(_07316_), .Y(_07317_));
NAND_g _28970_ (.A(_00012_[1]), .B(_07307_), .Y(_07318_));
AND_g _28971_ (.A(_00012_[3]), .B(_07317_), .Y(_07319_));
NAND_g _28972_ (.A(_07318_), .B(_07319_), .Y(_07320_));
AND_g _28973_ (.A(_13389_), .B(_07228_), .Y(_07321_));
NAND_g _28974_ (.A(_07231_), .B(_07321_), .Y(_07322_));
NAND_g _28975_ (.A(_00012_[4]), .B(_07276_), .Y(_07323_));
AND_g _28976_ (.A(_11216_), .B(_07298_), .Y(_07324_));
NAND_g _28977_ (.A(_07320_), .B(_07324_), .Y(_07325_));
AND_g _28978_ (.A(_13561_), .B(_07325_), .Y(_07326_));
AND_g _28979_ (.A(_07323_), .B(_07326_), .Y(_07327_));
NAND_g _28980_ (.A(_05765_), .B(_07327_), .Y(_07328_));
AND_g _28981_ (.A(_07225_), .B(_07328_), .Y(_07329_));
AND_g _28982_ (.A(_13425_), .B(_07329_), .Y(_07330_));
AND_g _28983_ (.A(_07322_), .B(_07330_), .Y(_07331_));
AND_g _28984_ (.A(_07224_), .B(_07331_), .Y(_07332_));
NOR_g _28985_ (.A(_07221_), .B(_07332_), .Y(_01228_));
NOR_g _28986_ (.A(pcpi_rs1[22]), .B(_13425_), .Y(_07333_));
XOR_g _28987_ (.A(_13449_), .B(_13534_), .Y(_07334_));
NAND_g _28988_ (.A(_13432_), .B(_07334_), .Y(_07335_));
NAND_g _28989_ (.A(_10946_), .B(_00012_[2]), .Y(_07336_));
NOR_g _28990_ (.A(cpuregs_2[22]), .B(_00012_[2]), .Y(_07337_));
NOR_g _28991_ (.A(_00012_[0]), .B(_07337_), .Y(_07338_));
NAND_g _28992_ (.A(_07336_), .B(_07338_), .Y(_07339_));
NAND_g _28993_ (.A(_11132_), .B(_00012_[2]), .Y(_07340_));
NOR_g _28994_ (.A(cpuregs_3[22]), .B(_00012_[2]), .Y(_07341_));
NOR_g _28995_ (.A(_11212_), .B(_07341_), .Y(_07342_));
NAND_g _28996_ (.A(_07340_), .B(_07342_), .Y(_07343_));
AND_g _28997_ (.A(_07339_), .B(_07343_), .Y(_07344_));
NAND_g _28998_ (.A(_10958_), .B(_00012_[2]), .Y(_07345_));
NOR_g _28999_ (.A(cpuregs_0[22]), .B(_00012_[2]), .Y(_07346_));
NOR_g _29000_ (.A(_00012_[0]), .B(_07346_), .Y(_07347_));
NAND_g _29001_ (.A(_07345_), .B(_07347_), .Y(_07348_));
NAND_g _29002_ (.A(_11116_), .B(_00012_[2]), .Y(_07349_));
NOR_g _29003_ (.A(cpuregs_1[22]), .B(_00012_[2]), .Y(_07350_));
NOR_g _29004_ (.A(_11212_), .B(_07350_), .Y(_07351_));
NAND_g _29005_ (.A(_07349_), .B(_07351_), .Y(_07352_));
NAND_g _29006_ (.A(_00012_[1]), .B(_07344_), .Y(_07353_));
AND_g _29007_ (.A(_11213_), .B(_07348_), .Y(_07354_));
NAND_g _29008_ (.A(_07352_), .B(_07354_), .Y(_07355_));
AND_g _29009_ (.A(_07353_), .B(_07355_), .Y(_07356_));
NAND_g _29010_ (.A(_11215_), .B(_07356_), .Y(_07357_));
NAND_g _29011_ (.A(cpuregs_13[22]), .B(_11213_), .Y(_07358_));
NAND_g _29012_ (.A(cpuregs_15[22]), .B(_00012_[1]), .Y(_07359_));
AND_g _29013_ (.A(_00012_[2]), .B(_07359_), .Y(_07360_));
NAND_g _29014_ (.A(_07358_), .B(_07360_), .Y(_07361_));
NAND_g _29015_ (.A(cpuregs_9[22]), .B(_11213_), .Y(_07362_));
NAND_g _29016_ (.A(cpuregs_11[22]), .B(_00012_[1]), .Y(_07363_));
AND_g _29017_ (.A(_11214_), .B(_07363_), .Y(_07364_));
NAND_g _29018_ (.A(_07362_), .B(_07364_), .Y(_07365_));
AND_g _29019_ (.A(_00012_[0]), .B(_07365_), .Y(_07366_));
NAND_g _29020_ (.A(_07361_), .B(_07366_), .Y(_07367_));
NAND_g _29021_ (.A(cpuregs_12[22]), .B(_11213_), .Y(_07368_));
NAND_g _29022_ (.A(cpuregs_14[22]), .B(_00012_[1]), .Y(_07369_));
AND_g _29023_ (.A(_00012_[2]), .B(_07369_), .Y(_07370_));
NAND_g _29024_ (.A(_07368_), .B(_07370_), .Y(_07371_));
NAND_g _29025_ (.A(cpuregs_8[22]), .B(_11213_), .Y(_07372_));
NAND_g _29026_ (.A(cpuregs_10[22]), .B(_00012_[1]), .Y(_07373_));
AND_g _29027_ (.A(_11214_), .B(_07373_), .Y(_07374_));
NAND_g _29028_ (.A(_07372_), .B(_07374_), .Y(_07375_));
AND_g _29029_ (.A(_11212_), .B(_07375_), .Y(_07376_));
NAND_g _29030_ (.A(_07371_), .B(_07376_), .Y(_07377_));
NAND_g _29031_ (.A(_07367_), .B(_07377_), .Y(_07378_));
NAND_g _29032_ (.A(_00012_[3]), .B(_07378_), .Y(_07379_));
AND_g _29033_ (.A(_11216_), .B(_07379_), .Y(_07380_));
NAND_g _29034_ (.A(_07357_), .B(_07380_), .Y(_07381_));
NAND_g _29035_ (.A(cpuregs_18[22]), .B(_00012_[1]), .Y(_07382_));
NAND_g _29036_ (.A(cpuregs_16[22]), .B(_11213_), .Y(_07383_));
NAND_g _29037_ (.A(_07382_), .B(_07383_), .Y(_07384_));
NAND_g _29038_ (.A(_11214_), .B(_07384_), .Y(_07385_));
NAND_g _29039_ (.A(cpuregs_22[22]), .B(_00012_[1]), .Y(_07386_));
NAND_g _29040_ (.A(cpuregs_20[22]), .B(_11213_), .Y(_07387_));
NAND_g _29041_ (.A(_07386_), .B(_07387_), .Y(_07388_));
NAND_g _29042_ (.A(_00012_[2]), .B(_07388_), .Y(_07389_));
AND_g _29043_ (.A(_11212_), .B(_07389_), .Y(_07390_));
NAND_g _29044_ (.A(_07385_), .B(_07390_), .Y(_07391_));
NAND_g _29045_ (.A(cpuregs_19[22]), .B(_00012_[1]), .Y(_07392_));
NAND_g _29046_ (.A(cpuregs_17[22]), .B(_11213_), .Y(_07393_));
NAND_g _29047_ (.A(_07392_), .B(_07393_), .Y(_07394_));
NAND_g _29048_ (.A(_11214_), .B(_07394_), .Y(_07395_));
NAND_g _29049_ (.A(cpuregs_23[22]), .B(_00012_[1]), .Y(_07396_));
NAND_g _29050_ (.A(cpuregs_21[22]), .B(_11213_), .Y(_07397_));
NAND_g _29051_ (.A(_07396_), .B(_07397_), .Y(_07398_));
NAND_g _29052_ (.A(_00012_[2]), .B(_07398_), .Y(_07399_));
AND_g _29053_ (.A(_00012_[0]), .B(_07399_), .Y(_07400_));
NAND_g _29054_ (.A(_07395_), .B(_07400_), .Y(_07401_));
AND_g _29055_ (.A(_07391_), .B(_07401_), .Y(_07402_));
NAND_g _29056_ (.A(cpuregs_24[22]), .B(_11214_), .Y(_07403_));
NAND_g _29057_ (.A(cpuregs_28[22]), .B(_00012_[2]), .Y(_07404_));
AND_g _29058_ (.A(_11212_), .B(_07404_), .Y(_07405_));
NAND_g _29059_ (.A(_07403_), .B(_07405_), .Y(_07406_));
NAND_g _29060_ (.A(cpuregs_29[22]), .B(_00012_[2]), .Y(_07407_));
NAND_g _29061_ (.A(cpuregs_25[22]), .B(_11214_), .Y(_07408_));
AND_g _29062_ (.A(_00012_[0]), .B(_07408_), .Y(_07409_));
NAND_g _29063_ (.A(_07407_), .B(_07409_), .Y(_07410_));
NAND_g _29064_ (.A(_07406_), .B(_07410_), .Y(_07411_));
NAND_g _29065_ (.A(_11213_), .B(_07411_), .Y(_07412_));
NAND_g _29066_ (.A(cpuregs_26[22]), .B(_11214_), .Y(_07413_));
NAND_g _29067_ (.A(cpuregs_30[22]), .B(_00012_[2]), .Y(_07414_));
AND_g _29068_ (.A(_11212_), .B(_07414_), .Y(_07415_));
NAND_g _29069_ (.A(_07413_), .B(_07415_), .Y(_07416_));
NAND_g _29070_ (.A(cpuregs_27[22]), .B(_11214_), .Y(_07417_));
NAND_g _29071_ (.A(cpuregs_31[22]), .B(_00012_[2]), .Y(_07418_));
AND_g _29072_ (.A(_00012_[0]), .B(_07418_), .Y(_07419_));
NAND_g _29073_ (.A(_07417_), .B(_07419_), .Y(_07420_));
NAND_g _29074_ (.A(_07416_), .B(_07420_), .Y(_07421_));
NAND_g _29075_ (.A(_00012_[1]), .B(_07421_), .Y(_07422_));
AND_g _29076_ (.A(_00012_[3]), .B(_07422_), .Y(_07423_));
NAND_g _29077_ (.A(_07412_), .B(_07423_), .Y(_07424_));
NAND_g _29078_ (.A(_11215_), .B(_07402_), .Y(_07425_));
AND_g _29079_ (.A(_07424_), .B(_07425_), .Y(_07426_));
NAND_g _29080_ (.A(_00012_[4]), .B(_07426_), .Y(_07427_));
AND_g _29081_ (.A(_13561_), .B(_07381_), .Y(_07428_));
AND_g _29082_ (.A(_07427_), .B(_07428_), .Y(_07429_));
NAND_g _29083_ (.A(_05765_), .B(_07429_), .Y(_07430_));
NAND_g _29084_ (.A(reg_pc[22]), .B(_13714_), .Y(_07431_));
NAND_g _29085_ (.A(pcpi_rs1[21]), .B(_13420_), .Y(_07432_));
AND_g _29086_ (.A(_07100_), .B(_07432_), .Y(_07433_));
NAND_g _29087_ (.A(_13382_), .B(_07433_), .Y(_07434_));
NAND_g _29088_ (.A(pcpi_rs1[26]), .B(_13419_), .Y(_07435_));
AND_g _29089_ (.A(_07097_), .B(_07435_), .Y(_07436_));
NAND_g _29090_ (.A(_13383_), .B(_07436_), .Y(_07437_));
AND_g _29091_ (.A(_07434_), .B(_07437_), .Y(_07438_));
NAND_g _29092_ (.A(_13389_), .B(_07438_), .Y(_07439_));
AND_g _29093_ (.A(_07431_), .B(_07439_), .Y(_07440_));
AND_g _29094_ (.A(_13425_), .B(_07440_), .Y(_07441_));
AND_g _29095_ (.A(_07430_), .B(_07441_), .Y(_07442_));
AND_g _29096_ (.A(_07335_), .B(_07442_), .Y(_07443_));
NOR_g _29097_ (.A(_07333_), .B(_07443_), .Y(_01229_));
NOR_g _29098_ (.A(pcpi_rs1[23]), .B(_13425_), .Y(_07444_));
NAND_g _29099_ (.A(cpuregs_13[23]), .B(_00012_[2]), .Y(_07445_));
NAND_g _29100_ (.A(cpuregs_9[23]), .B(_11214_), .Y(_07446_));
NAND_g _29101_ (.A(_07445_), .B(_07446_), .Y(_07447_));
NAND_g _29102_ (.A(_00012_[0]), .B(_07447_), .Y(_07448_));
NAND_g _29103_ (.A(cpuregs_12[23]), .B(_00012_[2]), .Y(_07449_));
NAND_g _29104_ (.A(cpuregs_8[23]), .B(_11214_), .Y(_07450_));
AND_g _29105_ (.A(_07449_), .B(_07450_), .Y(_07451_));
NOR_g _29106_ (.A(_00012_[0]), .B(_07451_), .Y(_07452_));
NAND_g _29107_ (.A(_10959_), .B(_00012_[2]), .Y(_07453_));
NOR_g _29108_ (.A(cpuregs_0[23]), .B(_00012_[2]), .Y(_07454_));
NOR_g _29109_ (.A(_00012_[0]), .B(_07454_), .Y(_07455_));
NAND_g _29110_ (.A(_07453_), .B(_07455_), .Y(_07456_));
NAND_g _29111_ (.A(_11117_), .B(_00012_[2]), .Y(_07457_));
NOR_g _29112_ (.A(cpuregs_1[23]), .B(_00012_[2]), .Y(_07458_));
NOR_g _29113_ (.A(_11212_), .B(_07458_), .Y(_07459_));
NAND_g _29114_ (.A(_07457_), .B(_07459_), .Y(_07460_));
NAND_g _29115_ (.A(cpuregs_11[23]), .B(_11214_), .Y(_07461_));
NAND_g _29116_ (.A(cpuregs_15[23]), .B(_00012_[2]), .Y(_07462_));
NAND_g _29117_ (.A(_07461_), .B(_07462_), .Y(_07463_));
AND_g _29118_ (.A(_00012_[0]), .B(_07463_), .Y(_07464_));
NAND_g _29119_ (.A(cpuregs_14[23]), .B(_00012_[2]), .Y(_07465_));
NAND_g _29120_ (.A(cpuregs_10[23]), .B(_11214_), .Y(_07466_));
AND_g _29121_ (.A(_07465_), .B(_07466_), .Y(_07467_));
NOR_g _29122_ (.A(_00012_[0]), .B(_07467_), .Y(_07468_));
NOR_g _29123_ (.A(_07464_), .B(_07468_), .Y(_07469_));
NAND_g _29124_ (.A(_10947_), .B(_00012_[2]), .Y(_07470_));
NOR_g _29125_ (.A(cpuregs_2[23]), .B(_00012_[2]), .Y(_07471_));
NOR_g _29126_ (.A(_00012_[0]), .B(_07471_), .Y(_07472_));
NAND_g _29127_ (.A(_07470_), .B(_07472_), .Y(_07473_));
NAND_g _29128_ (.A(_11133_), .B(_00012_[2]), .Y(_07474_));
NOR_g _29129_ (.A(cpuregs_3[23]), .B(_00012_[2]), .Y(_07475_));
NOR_g _29130_ (.A(_11212_), .B(_07475_), .Y(_07476_));
NAND_g _29131_ (.A(_07474_), .B(_07476_), .Y(_07477_));
AND_g _29132_ (.A(_07473_), .B(_07477_), .Y(_07478_));
NAND_g _29133_ (.A(_00012_[1]), .B(_07478_), .Y(_07479_));
AND_g _29134_ (.A(_11213_), .B(_07456_), .Y(_07480_));
NAND_g _29135_ (.A(_07460_), .B(_07480_), .Y(_07481_));
AND_g _29136_ (.A(_07479_), .B(_07481_), .Y(_07482_));
NAND_g _29137_ (.A(_11215_), .B(_07482_), .Y(_07483_));
NAND_g _29138_ (.A(_00012_[1]), .B(_07469_), .Y(_07484_));
NOR_g _29139_ (.A(_00012_[1]), .B(_07452_), .Y(_07485_));
NAND_g _29140_ (.A(_07448_), .B(_07485_), .Y(_07486_));
AND_g _29141_ (.A(_00012_[3]), .B(_07486_), .Y(_07487_));
NAND_g _29142_ (.A(_07484_), .B(_07487_), .Y(_07488_));
AND_g _29143_ (.A(_07483_), .B(_07488_), .Y(_07489_));
NAND_g _29144_ (.A(_11216_), .B(_07489_), .Y(_07490_));
NAND_g _29145_ (.A(cpuregs_31[23]), .B(_00012_[2]), .Y(_07491_));
NAND_g _29146_ (.A(cpuregs_27[23]), .B(_11214_), .Y(_07492_));
NAND_g _29147_ (.A(_07491_), .B(_07492_), .Y(_07493_));
AND_g _29148_ (.A(_00012_[0]), .B(_07493_), .Y(_07494_));
NAND_g _29149_ (.A(cpuregs_30[23]), .B(_00012_[2]), .Y(_07495_));
NAND_g _29150_ (.A(cpuregs_26[23]), .B(_11214_), .Y(_07496_));
AND_g _29151_ (.A(_07495_), .B(_07496_), .Y(_07497_));
NOR_g _29152_ (.A(_00012_[0]), .B(_07497_), .Y(_07498_));
NOR_g _29153_ (.A(_07494_), .B(_07498_), .Y(_07499_));
NAND_g _29154_ (.A(cpuregs_25[23]), .B(_11214_), .Y(_07500_));
NAND_g _29155_ (.A(cpuregs_29[23]), .B(_00012_[2]), .Y(_07501_));
NAND_g _29156_ (.A(_07500_), .B(_07501_), .Y(_07502_));
NAND_g _29157_ (.A(_00012_[0]), .B(_07502_), .Y(_07503_));
NAND_g _29158_ (.A(cpuregs_28[23]), .B(_00012_[2]), .Y(_07504_));
NAND_g _29159_ (.A(cpuregs_24[23]), .B(_11214_), .Y(_07505_));
NAND_g _29160_ (.A(_07504_), .B(_07505_), .Y(_07506_));
NAND_g _29161_ (.A(_11212_), .B(_07506_), .Y(_07507_));
AND_g _29162_ (.A(_07503_), .B(_07507_), .Y(_07508_));
NAND_g _29163_ (.A(_11213_), .B(_07508_), .Y(_07509_));
NAND_g _29164_ (.A(_00012_[1]), .B(_07499_), .Y(_07510_));
AND_g _29165_ (.A(_00012_[3]), .B(_07510_), .Y(_07511_));
NAND_g _29166_ (.A(_07509_), .B(_07511_), .Y(_07512_));
NAND_g _29167_ (.A(cpuregs_20[23]), .B(_11212_), .Y(_07513_));
NAND_g _29168_ (.A(cpuregs_21[23]), .B(_00012_[0]), .Y(_07514_));
AND_g _29169_ (.A(_00012_[2]), .B(_07514_), .Y(_07515_));
NAND_g _29170_ (.A(_07513_), .B(_07515_), .Y(_07516_));
NAND_g _29171_ (.A(cpuregs_16[23]), .B(_11212_), .Y(_07517_));
NAND_g _29172_ (.A(cpuregs_17[23]), .B(_00012_[0]), .Y(_07518_));
AND_g _29173_ (.A(_11214_), .B(_07518_), .Y(_07519_));
NAND_g _29174_ (.A(_07517_), .B(_07519_), .Y(_07520_));
AND_g _29175_ (.A(_11213_), .B(_07520_), .Y(_07521_));
NAND_g _29176_ (.A(_07516_), .B(_07521_), .Y(_07522_));
NAND_g _29177_ (.A(cpuregs_22[23]), .B(_00012_[2]), .Y(_07523_));
NAND_g _29178_ (.A(cpuregs_18[23]), .B(_11214_), .Y(_07524_));
AND_g _29179_ (.A(_11212_), .B(_07524_), .Y(_07525_));
NAND_g _29180_ (.A(_07523_), .B(_07525_), .Y(_07526_));
NAND_g _29181_ (.A(cpuregs_19[23]), .B(_11214_), .Y(_07527_));
NAND_g _29182_ (.A(cpuregs_23[23]), .B(_00012_[2]), .Y(_07528_));
AND_g _29183_ (.A(_00012_[0]), .B(_07528_), .Y(_07529_));
NAND_g _29184_ (.A(_07527_), .B(_07529_), .Y(_07530_));
AND_g _29185_ (.A(_00012_[1]), .B(_07530_), .Y(_07531_));
NAND_g _29186_ (.A(_07526_), .B(_07531_), .Y(_07532_));
NAND_g _29187_ (.A(_07522_), .B(_07532_), .Y(_07533_));
NAND_g _29188_ (.A(_11215_), .B(_07533_), .Y(_07534_));
AND_g _29189_ (.A(_00012_[4]), .B(_07534_), .Y(_07535_));
NAND_g _29190_ (.A(_07512_), .B(_07535_), .Y(_07536_));
AND_g _29191_ (.A(_07490_), .B(_07536_), .Y(_07537_));
AND_g _29192_ (.A(_13409_), .B(_07537_), .Y(_07538_));
AND_g _29193_ (.A(_13613_), .B(_07538_), .Y(_07539_));
NAND_g _29194_ (.A(reg_pc[23]), .B(_13714_), .Y(_07540_));
NAND_g _29195_ (.A(pcpi_rs1[27]), .B(_13419_), .Y(_07541_));
AND_g _29196_ (.A(_13383_), .B(_07114_), .Y(_07542_));
NAND_g _29197_ (.A(_07541_), .B(_07542_), .Y(_07543_));
NAND_g _29198_ (.A(pcpi_rs1[22]), .B(_13420_), .Y(_07544_));
AND_g _29199_ (.A(_13382_), .B(_07544_), .Y(_07545_));
NAND_g _29200_ (.A(_07111_), .B(_07545_), .Y(_07546_));
AND_g _29201_ (.A(_07543_), .B(_07546_), .Y(_07547_));
NAND_g _29202_ (.A(_13389_), .B(_07547_), .Y(_07548_));
AND_g _29203_ (.A(_07540_), .B(_07548_), .Y(_07549_));
NAND_g _29204_ (.A(_13425_), .B(_07549_), .Y(_07550_));
NOR_g _29205_ (.A(_07539_), .B(_07550_), .Y(_07551_));
XOR_g _29206_ (.A(decoded_imm[23]), .B(pcpi_rs1[23]), .Y(_07552_));
XNOR_g _29207_ (.A(_13536_), .B(_07552_), .Y(_07553_));
NAND_g _29208_ (.A(_13432_), .B(_07553_), .Y(_07554_));
AND_g _29209_ (.A(_07551_), .B(_07554_), .Y(_07555_));
NOR_g _29210_ (.A(_07444_), .B(_07555_), .Y(_01230_));
NOR_g _29211_ (.A(pcpi_rs1[24]), .B(_13425_), .Y(_07556_));
NAND_g _29212_ (.A(cpuregs_7[24]), .B(_00012_[2]), .Y(_07557_));
NAND_g _29213_ (.A(cpuregs_3[24]), .B(_11214_), .Y(_07558_));
NAND_g _29214_ (.A(_07557_), .B(_07558_), .Y(_07559_));
AND_g _29215_ (.A(_00012_[0]), .B(_07559_), .Y(_07560_));
NAND_g _29216_ (.A(cpuregs_6[24]), .B(_00012_[2]), .Y(_07561_));
NAND_g _29217_ (.A(cpuregs_2[24]), .B(_11214_), .Y(_07562_));
AND_g _29218_ (.A(_07561_), .B(_07562_), .Y(_07563_));
NOR_g _29219_ (.A(_00012_[0]), .B(_07563_), .Y(_07564_));
NOR_g _29220_ (.A(_07560_), .B(_07564_), .Y(_07565_));
NAND_g _29221_ (.A(cpuregs_5[24]), .B(_00012_[2]), .Y(_07566_));
NAND_g _29222_ (.A(cpuregs_1[24]), .B(_11214_), .Y(_07567_));
NAND_g _29223_ (.A(_07566_), .B(_07567_), .Y(_07568_));
NAND_g _29224_ (.A(_00012_[0]), .B(_07568_), .Y(_07569_));
NAND_g _29225_ (.A(cpuregs_4[24]), .B(_00012_[2]), .Y(_07570_));
NAND_g _29226_ (.A(cpuregs_0[24]), .B(_11214_), .Y(_07571_));
AND_g _29227_ (.A(_07570_), .B(_07571_), .Y(_07572_));
NOR_g _29228_ (.A(_00012_[0]), .B(_07572_), .Y(_07573_));
NAND_g _29229_ (.A(_00012_[1]), .B(_07565_), .Y(_07574_));
NOR_g _29230_ (.A(_00012_[1]), .B(_07573_), .Y(_07575_));
NAND_g _29231_ (.A(_07569_), .B(_07575_), .Y(_07576_));
AND_g _29232_ (.A(_07574_), .B(_07576_), .Y(_07577_));
NAND_g _29233_ (.A(_11215_), .B(_07577_), .Y(_07578_));
NAND_g _29234_ (.A(cpuregs_13[24]), .B(_00012_[0]), .Y(_07579_));
NAND_g _29235_ (.A(cpuregs_12[24]), .B(_11212_), .Y(_07580_));
AND_g _29236_ (.A(_00012_[2]), .B(_07580_), .Y(_07581_));
NAND_g _29237_ (.A(_07579_), .B(_07581_), .Y(_07582_));
NAND_g _29238_ (.A(cpuregs_9[24]), .B(_00012_[0]), .Y(_07583_));
NAND_g _29239_ (.A(cpuregs_8[24]), .B(_11212_), .Y(_07584_));
AND_g _29240_ (.A(_11214_), .B(_07584_), .Y(_07585_));
NAND_g _29241_ (.A(_07583_), .B(_07585_), .Y(_07586_));
AND_g _29242_ (.A(_11213_), .B(_07586_), .Y(_07587_));
NAND_g _29243_ (.A(_07582_), .B(_07587_), .Y(_07588_));
NAND_g _29244_ (.A(cpuregs_15[24]), .B(_00012_[0]), .Y(_07589_));
NAND_g _29245_ (.A(cpuregs_14[24]), .B(_11212_), .Y(_07590_));
AND_g _29246_ (.A(_00012_[2]), .B(_07590_), .Y(_07591_));
NAND_g _29247_ (.A(_07589_), .B(_07591_), .Y(_07592_));
NAND_g _29248_ (.A(cpuregs_11[24]), .B(_00012_[0]), .Y(_07593_));
NAND_g _29249_ (.A(cpuregs_10[24]), .B(_11212_), .Y(_07594_));
AND_g _29250_ (.A(_11214_), .B(_07594_), .Y(_07595_));
NAND_g _29251_ (.A(_07593_), .B(_07595_), .Y(_07596_));
AND_g _29252_ (.A(_00012_[1]), .B(_07596_), .Y(_07597_));
NAND_g _29253_ (.A(_07592_), .B(_07597_), .Y(_07598_));
NAND_g _29254_ (.A(_07588_), .B(_07598_), .Y(_07599_));
NAND_g _29255_ (.A(_00012_[3]), .B(_07599_), .Y(_07600_));
AND_g _29256_ (.A(_07578_), .B(_07600_), .Y(_07601_));
NAND_g _29257_ (.A(_11216_), .B(_07601_), .Y(_07602_));
NAND_g _29258_ (.A(cpuregs_23[24]), .B(_00012_[0]), .Y(_07603_));
NAND_g _29259_ (.A(cpuregs_22[24]), .B(_11212_), .Y(_07604_));
NAND_g _29260_ (.A(_07603_), .B(_07604_), .Y(_07605_));
NAND_g _29261_ (.A(_00012_[2]), .B(_07605_), .Y(_07606_));
NAND_g _29262_ (.A(cpuregs_19[24]), .B(_00012_[0]), .Y(_07607_));
NAND_g _29263_ (.A(cpuregs_18[24]), .B(_11212_), .Y(_07608_));
NAND_g _29264_ (.A(_07607_), .B(_07608_), .Y(_07609_));
NAND_g _29265_ (.A(_11214_), .B(_07609_), .Y(_07610_));
NAND_g _29266_ (.A(_07606_), .B(_07610_), .Y(_07611_));
NAND_g _29267_ (.A(_00012_[1]), .B(_07611_), .Y(_07612_));
NAND_g _29268_ (.A(cpuregs_20[24]), .B(_00012_[2]), .Y(_07613_));
NAND_g _29269_ (.A(cpuregs_16[24]), .B(_11214_), .Y(_07614_));
AND_g _29270_ (.A(_07613_), .B(_07614_), .Y(_07615_));
NAND_g _29271_ (.A(_11212_), .B(_07615_), .Y(_07616_));
NAND_g _29272_ (.A(cpuregs_21[24]), .B(_00012_[2]), .Y(_07617_));
NAND_g _29273_ (.A(cpuregs_17[24]), .B(_11214_), .Y(_07618_));
AND_g _29274_ (.A(_00012_[0]), .B(_07618_), .Y(_07619_));
NAND_g _29275_ (.A(_07617_), .B(_07619_), .Y(_07620_));
AND_g _29276_ (.A(_07616_), .B(_07620_), .Y(_07621_));
NAND_g _29277_ (.A(_11213_), .B(_07621_), .Y(_07622_));
NAND_g _29278_ (.A(_07612_), .B(_07622_), .Y(_07623_));
NAND_g _29279_ (.A(_11215_), .B(_07623_), .Y(_07624_));
NAND_g _29280_ (.A(cpuregs_29[24]), .B(_11213_), .Y(_07625_));
NAND_g _29281_ (.A(cpuregs_31[24]), .B(_00012_[1]), .Y(_07626_));
AND_g _29282_ (.A(_00012_[2]), .B(_07626_), .Y(_07627_));
NAND_g _29283_ (.A(_07625_), .B(_07627_), .Y(_07628_));
NAND_g _29284_ (.A(cpuregs_25[24]), .B(_11213_), .Y(_07629_));
NAND_g _29285_ (.A(cpuregs_27[24]), .B(_00012_[1]), .Y(_07630_));
AND_g _29286_ (.A(_11214_), .B(_07630_), .Y(_07631_));
NAND_g _29287_ (.A(_07629_), .B(_07631_), .Y(_07632_));
AND_g _29288_ (.A(_00012_[0]), .B(_07632_), .Y(_07633_));
NAND_g _29289_ (.A(_07628_), .B(_07633_), .Y(_07634_));
NAND_g _29290_ (.A(cpuregs_28[24]), .B(_11213_), .Y(_07635_));
NAND_g _29291_ (.A(cpuregs_30[24]), .B(_00012_[1]), .Y(_07636_));
AND_g _29292_ (.A(_00012_[2]), .B(_07636_), .Y(_07637_));
NAND_g _29293_ (.A(_07635_), .B(_07637_), .Y(_07638_));
NAND_g _29294_ (.A(cpuregs_24[24]), .B(_11213_), .Y(_07639_));
NAND_g _29295_ (.A(cpuregs_26[24]), .B(_00012_[1]), .Y(_07640_));
AND_g _29296_ (.A(_11214_), .B(_07640_), .Y(_07641_));
NAND_g _29297_ (.A(_07639_), .B(_07641_), .Y(_07642_));
AND_g _29298_ (.A(_11212_), .B(_07642_), .Y(_07643_));
NAND_g _29299_ (.A(_07638_), .B(_07643_), .Y(_07644_));
NAND_g _29300_ (.A(_07634_), .B(_07644_), .Y(_07645_));
NAND_g _29301_ (.A(_00012_[3]), .B(_07645_), .Y(_07646_));
AND_g _29302_ (.A(_00012_[4]), .B(_07646_), .Y(_07647_));
NAND_g _29303_ (.A(_07624_), .B(_07647_), .Y(_07648_));
AND_g _29304_ (.A(_07602_), .B(_07648_), .Y(_07649_));
AND_g _29305_ (.A(_13409_), .B(_07649_), .Y(_07650_));
AND_g _29306_ (.A(_13613_), .B(_07650_), .Y(_07651_));
NAND_g _29307_ (.A(reg_pc[24]), .B(_13714_), .Y(_07652_));
NAND_g _29308_ (.A(pcpi_rs1[28]), .B(_13419_), .Y(_07653_));
AND_g _29309_ (.A(_13383_), .B(_07653_), .Y(_07654_));
NAND_g _29310_ (.A(_07226_), .B(_07654_), .Y(_07655_));
NAND_g _29311_ (.A(pcpi_rs1[23]), .B(_13420_), .Y(_07656_));
AND_g _29312_ (.A(_13382_), .B(_07656_), .Y(_07657_));
NAND_g _29313_ (.A(_07229_), .B(_07657_), .Y(_07658_));
AND_g _29314_ (.A(_07655_), .B(_07658_), .Y(_07659_));
NAND_g _29315_ (.A(_13389_), .B(_07659_), .Y(_07660_));
AND_g _29316_ (.A(_07652_), .B(_07660_), .Y(_07661_));
NAND_g _29317_ (.A(_13425_), .B(_07661_), .Y(_07662_));
NOR_g _29318_ (.A(_07651_), .B(_07662_), .Y(_07663_));
XOR_g _29319_ (.A(_13445_), .B(_13538_), .Y(_07664_));
NAND_g _29320_ (.A(_13432_), .B(_07664_), .Y(_07665_));
AND_g _29321_ (.A(_07663_), .B(_07665_), .Y(_07666_));
NOR_g _29322_ (.A(_07556_), .B(_07666_), .Y(_01231_));
NOR_g _29323_ (.A(pcpi_rs1[25]), .B(_13425_), .Y(_07667_));
XOR_g _29324_ (.A(_13540_), .B(_13541_), .Y(_07668_));
NAND_g _29325_ (.A(_13432_), .B(_07668_), .Y(_07669_));
NAND_g _29326_ (.A(cpuregs_23[25]), .B(_00012_[0]), .Y(_07670_));
NAND_g _29327_ (.A(cpuregs_22[25]), .B(_11212_), .Y(_07671_));
AND_g _29328_ (.A(_00012_[2]), .B(_07671_), .Y(_07672_));
NAND_g _29329_ (.A(_07670_), .B(_07672_), .Y(_07673_));
NAND_g _29330_ (.A(cpuregs_19[25]), .B(_00012_[0]), .Y(_07674_));
NAND_g _29331_ (.A(cpuregs_18[25]), .B(_11212_), .Y(_07675_));
AND_g _29332_ (.A(_11214_), .B(_07675_), .Y(_07676_));
NAND_g _29333_ (.A(_07674_), .B(_07676_), .Y(_07677_));
AND_g _29334_ (.A(_11215_), .B(_07677_), .Y(_07678_));
NAND_g _29335_ (.A(_07673_), .B(_07678_), .Y(_07679_));
NAND_g _29336_ (.A(cpuregs_31[25]), .B(_00012_[0]), .Y(_07680_));
NAND_g _29337_ (.A(cpuregs_30[25]), .B(_11212_), .Y(_07681_));
AND_g _29338_ (.A(_00012_[2]), .B(_07681_), .Y(_07682_));
NAND_g _29339_ (.A(_07680_), .B(_07682_), .Y(_07683_));
NAND_g _29340_ (.A(cpuregs_27[25]), .B(_00012_[0]), .Y(_07684_));
NAND_g _29341_ (.A(cpuregs_26[25]), .B(_11212_), .Y(_07685_));
AND_g _29342_ (.A(_11214_), .B(_07685_), .Y(_07686_));
NAND_g _29343_ (.A(_07684_), .B(_07686_), .Y(_07687_));
AND_g _29344_ (.A(_00012_[3]), .B(_07687_), .Y(_07688_));
NAND_g _29345_ (.A(_07683_), .B(_07688_), .Y(_07689_));
NAND_g _29346_ (.A(_07679_), .B(_07689_), .Y(_07690_));
NAND_g _29347_ (.A(_00012_[4]), .B(_07690_), .Y(_07691_));
NAND_g _29348_ (.A(cpuregs_6[25]), .B(_00012_[2]), .Y(_07692_));
NAND_g _29349_ (.A(cpuregs_2[25]), .B(_11214_), .Y(_07693_));
AND_g _29350_ (.A(_07692_), .B(_07693_), .Y(_07694_));
NAND_g _29351_ (.A(_11212_), .B(_07694_), .Y(_07695_));
NAND_g _29352_ (.A(cpuregs_7[25]), .B(_00012_[2]), .Y(_07696_));
NAND_g _29353_ (.A(cpuregs_3[25]), .B(_11214_), .Y(_07697_));
AND_g _29354_ (.A(_00012_[0]), .B(_07697_), .Y(_07698_));
NAND_g _29355_ (.A(_07696_), .B(_07698_), .Y(_07699_));
AND_g _29356_ (.A(_07695_), .B(_07699_), .Y(_07700_));
NAND_g _29357_ (.A(_11215_), .B(_07700_), .Y(_07701_));
NOR_g _29358_ (.A(cpuregs_10[25]), .B(_00012_[2]), .Y(_07702_));
NOR_g _29359_ (.A(cpuregs_14[25]), .B(_11214_), .Y(_07703_));
NOR_g _29360_ (.A(_07702_), .B(_07703_), .Y(_07704_));
NOR_g _29361_ (.A(cpuregs_11[25]), .B(_00012_[2]), .Y(_07705_));
NOT_g _29362_ (.A(_07705_), .Y(_07706_));
NAND_g _29363_ (.A(_11169_), .B(_00012_[2]), .Y(_07707_));
AND_g _29364_ (.A(_00012_[0]), .B(_07707_), .Y(_07708_));
NAND_g _29365_ (.A(_07706_), .B(_07708_), .Y(_07709_));
NAND_g _29366_ (.A(_11212_), .B(_07704_), .Y(_07710_));
NAND_g _29367_ (.A(_07709_), .B(_07710_), .Y(_07711_));
NAND_g _29368_ (.A(_00012_[3]), .B(_07711_), .Y(_07712_));
NAND_g _29369_ (.A(_07701_), .B(_07712_), .Y(_07713_));
AND_g _29370_ (.A(_11216_), .B(_07713_), .Y(_07714_));
NOT_g _29371_ (.A(_07714_), .Y(_07715_));
NAND_g _29372_ (.A(_07691_), .B(_07715_), .Y(_07716_));
NAND_g _29373_ (.A(_00012_[1]), .B(_07716_), .Y(_07717_));
NAND_g _29374_ (.A(cpuregs_4[25]), .B(_00012_[2]), .Y(_07718_));
NAND_g _29375_ (.A(cpuregs_0[25]), .B(_11214_), .Y(_07719_));
AND_g _29376_ (.A(_07718_), .B(_07719_), .Y(_07720_));
NAND_g _29377_ (.A(_11212_), .B(_07720_), .Y(_07721_));
NAND_g _29378_ (.A(cpuregs_5[25]), .B(_00012_[2]), .Y(_07722_));
NAND_g _29379_ (.A(cpuregs_1[25]), .B(_11214_), .Y(_07723_));
AND_g _29380_ (.A(_00012_[0]), .B(_07723_), .Y(_07724_));
NAND_g _29381_ (.A(_07722_), .B(_07724_), .Y(_07725_));
AND_g _29382_ (.A(_11215_), .B(_07725_), .Y(_07726_));
NAND_g _29383_ (.A(_07721_), .B(_07726_), .Y(_07727_));
NAND_g _29384_ (.A(_10935_), .B(_11214_), .Y(_07728_));
NAND_g _29385_ (.A(_11153_), .B(_00012_[2]), .Y(_07729_));
NOR_g _29386_ (.A(cpuregs_8[25]), .B(_00012_[2]), .Y(_07730_));
NOR_g _29387_ (.A(cpuregs_12[25]), .B(_11214_), .Y(_07731_));
NOR_g _29388_ (.A(_07730_), .B(_07731_), .Y(_07732_));
AND_g _29389_ (.A(_00012_[0]), .B(_07729_), .Y(_07733_));
NAND_g _29390_ (.A(_07728_), .B(_07733_), .Y(_07734_));
NAND_g _29391_ (.A(_11212_), .B(_07732_), .Y(_07735_));
NAND_g _29392_ (.A(_07734_), .B(_07735_), .Y(_07736_));
NAND_g _29393_ (.A(_00012_[3]), .B(_07736_), .Y(_07737_));
NAND_g _29394_ (.A(_07727_), .B(_07737_), .Y(_07738_));
NAND_g _29395_ (.A(_11216_), .B(_07738_), .Y(_07739_));
NAND_g _29396_ (.A(cpuregs_25[25]), .B(_00012_[3]), .Y(_07740_));
NAND_g _29397_ (.A(cpuregs_17[25]), .B(_11215_), .Y(_07741_));
NAND_g _29398_ (.A(_07740_), .B(_07741_), .Y(_07742_));
NAND_g _29399_ (.A(_11214_), .B(_07742_), .Y(_07743_));
NAND_g _29400_ (.A(cpuregs_29[25]), .B(_00012_[3]), .Y(_07744_));
NAND_g _29401_ (.A(cpuregs_21[25]), .B(_11215_), .Y(_07745_));
NAND_g _29402_ (.A(_07744_), .B(_07745_), .Y(_07746_));
NAND_g _29403_ (.A(_00012_[2]), .B(_07746_), .Y(_07747_));
AND_g _29404_ (.A(_00012_[0]), .B(_07747_), .Y(_07748_));
NAND_g _29405_ (.A(_07743_), .B(_07748_), .Y(_07749_));
NAND_g _29406_ (.A(cpuregs_24[25]), .B(_00012_[3]), .Y(_07750_));
NAND_g _29407_ (.A(cpuregs_16[25]), .B(_11215_), .Y(_07751_));
NAND_g _29408_ (.A(_07750_), .B(_07751_), .Y(_07752_));
NAND_g _29409_ (.A(_11214_), .B(_07752_), .Y(_07753_));
NAND_g _29410_ (.A(cpuregs_28[25]), .B(_00012_[3]), .Y(_07754_));
NAND_g _29411_ (.A(cpuregs_20[25]), .B(_11215_), .Y(_07755_));
NAND_g _29412_ (.A(_07754_), .B(_07755_), .Y(_07756_));
NAND_g _29413_ (.A(_00012_[2]), .B(_07756_), .Y(_07757_));
AND_g _29414_ (.A(_11212_), .B(_07757_), .Y(_07758_));
NAND_g _29415_ (.A(_07753_), .B(_07758_), .Y(_07759_));
AND_g _29416_ (.A(_00012_[4]), .B(_07759_), .Y(_07760_));
NAND_g _29417_ (.A(_07749_), .B(_07760_), .Y(_07761_));
NAND_g _29418_ (.A(_07739_), .B(_07761_), .Y(_07762_));
NAND_g _29419_ (.A(_11213_), .B(_07762_), .Y(_07763_));
NAND_g _29420_ (.A(_07717_), .B(_07763_), .Y(_07764_));
NAND_g _29421_ (.A(reg_pc[25]), .B(_13714_), .Y(_07765_));
NAND_g _29422_ (.A(pcpi_rs1[29]), .B(_13419_), .Y(_07766_));
AND_g _29423_ (.A(_13383_), .B(_07766_), .Y(_07767_));
NAND_g _29424_ (.A(_07432_), .B(_07767_), .Y(_07768_));
NAND_g _29425_ (.A(pcpi_rs1[24]), .B(_13420_), .Y(_07769_));
AND_g _29426_ (.A(_13382_), .B(_07769_), .Y(_07770_));
NAND_g _29427_ (.A(_07435_), .B(_07770_), .Y(_07771_));
AND_g _29428_ (.A(_13561_), .B(_07764_), .Y(_07772_));
NAND_g _29429_ (.A(_05765_), .B(_07772_), .Y(_07773_));
AND_g _29430_ (.A(_13389_), .B(_07768_), .Y(_07774_));
NAND_g _29431_ (.A(_07771_), .B(_07774_), .Y(_07775_));
AND_g _29432_ (.A(_07773_), .B(_07775_), .Y(_07776_));
AND_g _29433_ (.A(_13425_), .B(_07776_), .Y(_07777_));
AND_g _29434_ (.A(_07765_), .B(_07777_), .Y(_07778_));
AND_g _29435_ (.A(_07669_), .B(_07778_), .Y(_07779_));
NOR_g _29436_ (.A(_07667_), .B(_07779_), .Y(_01232_));
NOR_g _29437_ (.A(pcpi_rs1[26]), .B(_13425_), .Y(_07780_));
XOR_g _29438_ (.A(_13442_), .B(_13543_), .Y(_07781_));
NAND_g _29439_ (.A(_13432_), .B(_07781_), .Y(_07782_));
NAND_g _29440_ (.A(cpuregs_7[26]), .B(_00012_[2]), .Y(_07783_));
NAND_g _29441_ (.A(cpuregs_3[26]), .B(_11214_), .Y(_07784_));
NAND_g _29442_ (.A(_07783_), .B(_07784_), .Y(_07785_));
AND_g _29443_ (.A(_00012_[0]), .B(_07785_), .Y(_07786_));
NAND_g _29444_ (.A(cpuregs_6[26]), .B(_00012_[2]), .Y(_07787_));
NAND_g _29445_ (.A(cpuregs_2[26]), .B(_11214_), .Y(_07788_));
AND_g _29446_ (.A(_07787_), .B(_07788_), .Y(_07789_));
NOR_g _29447_ (.A(_00012_[0]), .B(_07789_), .Y(_07790_));
NOR_g _29448_ (.A(_07786_), .B(_07790_), .Y(_07791_));
NAND_g _29449_ (.A(cpuregs_5[26]), .B(_00012_[2]), .Y(_07792_));
NAND_g _29450_ (.A(cpuregs_1[26]), .B(_11214_), .Y(_07793_));
NAND_g _29451_ (.A(_07792_), .B(_07793_), .Y(_07794_));
NAND_g _29452_ (.A(_00012_[0]), .B(_07794_), .Y(_07795_));
NAND_g _29453_ (.A(cpuregs_4[26]), .B(_00012_[2]), .Y(_07796_));
NAND_g _29454_ (.A(cpuregs_0[26]), .B(_11214_), .Y(_07797_));
AND_g _29455_ (.A(_07796_), .B(_07797_), .Y(_07798_));
NOR_g _29456_ (.A(_00012_[0]), .B(_07798_), .Y(_07799_));
NAND_g _29457_ (.A(_00012_[1]), .B(_07791_), .Y(_07800_));
NOR_g _29458_ (.A(_00012_[1]), .B(_07799_), .Y(_07801_));
NAND_g _29459_ (.A(_07795_), .B(_07801_), .Y(_07802_));
AND_g _29460_ (.A(_07800_), .B(_07802_), .Y(_07803_));
NAND_g _29461_ (.A(_11215_), .B(_07803_), .Y(_07804_));
NAND_g _29462_ (.A(cpuregs_13[26]), .B(_00012_[0]), .Y(_07805_));
NAND_g _29463_ (.A(cpuregs_12[26]), .B(_11212_), .Y(_07806_));
AND_g _29464_ (.A(_00012_[2]), .B(_07806_), .Y(_07807_));
NAND_g _29465_ (.A(_07805_), .B(_07807_), .Y(_07808_));
NAND_g _29466_ (.A(cpuregs_9[26]), .B(_00012_[0]), .Y(_07809_));
NAND_g _29467_ (.A(cpuregs_8[26]), .B(_11212_), .Y(_07810_));
AND_g _29468_ (.A(_11214_), .B(_07810_), .Y(_07811_));
NAND_g _29469_ (.A(_07809_), .B(_07811_), .Y(_07812_));
AND_g _29470_ (.A(_11213_), .B(_07812_), .Y(_07813_));
NAND_g _29471_ (.A(_07808_), .B(_07813_), .Y(_07814_));
NAND_g _29472_ (.A(cpuregs_15[26]), .B(_00012_[0]), .Y(_07815_));
NAND_g _29473_ (.A(cpuregs_14[26]), .B(_11212_), .Y(_07816_));
AND_g _29474_ (.A(_00012_[2]), .B(_07816_), .Y(_07817_));
NAND_g _29475_ (.A(_07815_), .B(_07817_), .Y(_07818_));
NAND_g _29476_ (.A(cpuregs_11[26]), .B(_00012_[0]), .Y(_07819_));
NAND_g _29477_ (.A(cpuregs_10[26]), .B(_11212_), .Y(_07820_));
AND_g _29478_ (.A(_11214_), .B(_07820_), .Y(_07821_));
NAND_g _29479_ (.A(_07819_), .B(_07821_), .Y(_07822_));
AND_g _29480_ (.A(_00012_[1]), .B(_07822_), .Y(_07823_));
NAND_g _29481_ (.A(_07818_), .B(_07823_), .Y(_07824_));
NAND_g _29482_ (.A(_07814_), .B(_07824_), .Y(_07825_));
NAND_g _29483_ (.A(_00012_[3]), .B(_07825_), .Y(_07826_));
AND_g _29484_ (.A(_07804_), .B(_07826_), .Y(_07827_));
NAND_g _29485_ (.A(_11216_), .B(_07827_), .Y(_07828_));
NAND_g _29486_ (.A(_11020_), .B(_00012_[2]), .Y(_07829_));
NOR_g _29487_ (.A(cpuregs_18[26]), .B(_00012_[2]), .Y(_07830_));
NOR_g _29488_ (.A(_00012_[0]), .B(_07830_), .Y(_07831_));
NAND_g _29489_ (.A(_07829_), .B(_07831_), .Y(_07832_));
NAND_g _29490_ (.A(_11189_), .B(_00012_[2]), .Y(_07833_));
NOR_g _29491_ (.A(cpuregs_19[26]), .B(_00012_[2]), .Y(_07834_));
NOR_g _29492_ (.A(_11212_), .B(_07834_), .Y(_07835_));
NAND_g _29493_ (.A(_07833_), .B(_07835_), .Y(_07836_));
AND_g _29494_ (.A(_07832_), .B(_07836_), .Y(_07837_));
NAND_g _29495_ (.A(_11201_), .B(_00012_[2]), .Y(_07838_));
NOR_g _29496_ (.A(cpuregs_16[26]), .B(_00012_[2]), .Y(_07839_));
NOR_g _29497_ (.A(_00012_[0]), .B(_07839_), .Y(_07840_));
NAND_g _29498_ (.A(_07838_), .B(_07840_), .Y(_07841_));
NAND_g _29499_ (.A(_11036_), .B(_00012_[2]), .Y(_07842_));
NOR_g _29500_ (.A(cpuregs_17[26]), .B(_00012_[2]), .Y(_07843_));
NOR_g _29501_ (.A(_11212_), .B(_07843_), .Y(_07844_));
NAND_g _29502_ (.A(_07842_), .B(_07844_), .Y(_07845_));
AND_g _29503_ (.A(_07841_), .B(_07845_), .Y(_07846_));
NAND_g _29504_ (.A(_00012_[1]), .B(_07837_), .Y(_07847_));
NAND_g _29505_ (.A(_11213_), .B(_07846_), .Y(_07848_));
AND_g _29506_ (.A(_07847_), .B(_07848_), .Y(_07849_));
NAND_g _29507_ (.A(_11215_), .B(_07849_), .Y(_07850_));
NAND_g _29508_ (.A(cpuregs_29[26]), .B(_11213_), .Y(_07851_));
NAND_g _29509_ (.A(cpuregs_31[26]), .B(_00012_[1]), .Y(_07852_));
AND_g _29510_ (.A(_00012_[2]), .B(_07852_), .Y(_07853_));
NAND_g _29511_ (.A(_07851_), .B(_07853_), .Y(_07854_));
NAND_g _29512_ (.A(cpuregs_25[26]), .B(_11213_), .Y(_07855_));
NAND_g _29513_ (.A(cpuregs_27[26]), .B(_00012_[1]), .Y(_07856_));
AND_g _29514_ (.A(_11214_), .B(_07856_), .Y(_07857_));
NAND_g _29515_ (.A(_07855_), .B(_07857_), .Y(_07858_));
AND_g _29516_ (.A(_00012_[0]), .B(_07858_), .Y(_07859_));
NAND_g _29517_ (.A(_07854_), .B(_07859_), .Y(_07860_));
NAND_g _29518_ (.A(cpuregs_28[26]), .B(_11213_), .Y(_07861_));
NAND_g _29519_ (.A(cpuregs_30[26]), .B(_00012_[1]), .Y(_07862_));
AND_g _29520_ (.A(_00012_[2]), .B(_07862_), .Y(_07863_));
NAND_g _29521_ (.A(_07861_), .B(_07863_), .Y(_07864_));
NAND_g _29522_ (.A(cpuregs_24[26]), .B(_11213_), .Y(_07865_));
NAND_g _29523_ (.A(cpuregs_26[26]), .B(_00012_[1]), .Y(_07866_));
AND_g _29524_ (.A(_11214_), .B(_07866_), .Y(_07867_));
NAND_g _29525_ (.A(_07865_), .B(_07867_), .Y(_07868_));
AND_g _29526_ (.A(_11212_), .B(_07868_), .Y(_07869_));
NAND_g _29527_ (.A(_07864_), .B(_07869_), .Y(_07870_));
NAND_g _29528_ (.A(_07860_), .B(_07870_), .Y(_07871_));
NAND_g _29529_ (.A(_00012_[3]), .B(_07871_), .Y(_07872_));
AND_g _29530_ (.A(_07850_), .B(_07872_), .Y(_07873_));
NAND_g _29531_ (.A(_00012_[4]), .B(_07873_), .Y(_07874_));
AND_g _29532_ (.A(_13409_), .B(_07874_), .Y(_07875_));
AND_g _29533_ (.A(_07828_), .B(_07875_), .Y(_07876_));
AND_g _29534_ (.A(_13613_), .B(_07876_), .Y(_07877_));
NAND_g _29535_ (.A(reg_pc[26]), .B(_13714_), .Y(_07878_));
NAND_g _29536_ (.A(pcpi_rs1[30]), .B(_13419_), .Y(_07879_));
AND_g _29537_ (.A(_13383_), .B(_07879_), .Y(_07880_));
NAND_g _29538_ (.A(_07544_), .B(_07880_), .Y(_07881_));
NAND_g _29539_ (.A(pcpi_rs1[25]), .B(_13420_), .Y(_07882_));
AND_g _29540_ (.A(_13382_), .B(_07882_), .Y(_07883_));
NAND_g _29541_ (.A(_07541_), .B(_07883_), .Y(_07884_));
AND_g _29542_ (.A(_07881_), .B(_07884_), .Y(_07885_));
NAND_g _29543_ (.A(_13389_), .B(_07885_), .Y(_07886_));
AND_g _29544_ (.A(_07878_), .B(_07886_), .Y(_07887_));
NAND_g _29545_ (.A(_13425_), .B(_07887_), .Y(_07888_));
NOR_g _29546_ (.A(_07877_), .B(_07888_), .Y(_07889_));
AND_g _29547_ (.A(_07782_), .B(_07889_), .Y(_07890_));
NOR_g _29548_ (.A(_07780_), .B(_07890_), .Y(_01233_));
NOR_g _29549_ (.A(pcpi_rs1[27]), .B(_13425_), .Y(_07891_));
XOR_g _29550_ (.A(decoded_imm[27]), .B(pcpi_rs1[27]), .Y(_07892_));
XNOR_g _29551_ (.A(_13545_), .B(_07892_), .Y(_07893_));
NAND_g _29552_ (.A(_13432_), .B(_07893_), .Y(_07894_));
NAND_g _29553_ (.A(reg_pc[27]), .B(_13714_), .Y(_07895_));
NAND_g _29554_ (.A(pcpi_rs1[31]), .B(_13419_), .Y(_07896_));
AND_g _29555_ (.A(_13383_), .B(_07656_), .Y(_07897_));
NAND_g _29556_ (.A(_07896_), .B(_07897_), .Y(_07898_));
NAND_g _29557_ (.A(pcpi_rs1[26]), .B(_13420_), .Y(_07899_));
AND_g _29558_ (.A(_13382_), .B(_07899_), .Y(_07900_));
NAND_g _29559_ (.A(_07653_), .B(_07900_), .Y(_07901_));
AND_g _29560_ (.A(_07898_), .B(_07901_), .Y(_07902_));
NAND_g _29561_ (.A(_13389_), .B(_07902_), .Y(_07903_));
AND_g _29562_ (.A(_07895_), .B(_07903_), .Y(_07904_));
AND_g _29563_ (.A(_13425_), .B(_07904_), .Y(_07905_));
NAND_g _29564_ (.A(cpuregs_23[27]), .B(_00012_[0]), .Y(_07906_));
NAND_g _29565_ (.A(cpuregs_22[27]), .B(_11212_), .Y(_07907_));
AND_g _29566_ (.A(_00012_[2]), .B(_07907_), .Y(_07908_));
NAND_g _29567_ (.A(_07906_), .B(_07908_), .Y(_07909_));
NAND_g _29568_ (.A(cpuregs_19[27]), .B(_00012_[0]), .Y(_07910_));
NAND_g _29569_ (.A(cpuregs_18[27]), .B(_11212_), .Y(_07911_));
AND_g _29570_ (.A(_11214_), .B(_07911_), .Y(_07912_));
NAND_g _29571_ (.A(_07910_), .B(_07912_), .Y(_07913_));
AND_g _29572_ (.A(_11215_), .B(_07913_), .Y(_07914_));
NAND_g _29573_ (.A(_07909_), .B(_07914_), .Y(_07915_));
NAND_g _29574_ (.A(cpuregs_31[27]), .B(_00012_[0]), .Y(_07916_));
NAND_g _29575_ (.A(cpuregs_30[27]), .B(_11212_), .Y(_07917_));
AND_g _29576_ (.A(_00012_[2]), .B(_07917_), .Y(_07918_));
NAND_g _29577_ (.A(_07916_), .B(_07918_), .Y(_07919_));
NAND_g _29578_ (.A(cpuregs_27[27]), .B(_00012_[0]), .Y(_07920_));
NAND_g _29579_ (.A(cpuregs_26[27]), .B(_11212_), .Y(_07921_));
AND_g _29580_ (.A(_11214_), .B(_07921_), .Y(_07922_));
NAND_g _29581_ (.A(_07920_), .B(_07922_), .Y(_07923_));
AND_g _29582_ (.A(_00012_[3]), .B(_07923_), .Y(_07924_));
NAND_g _29583_ (.A(_07919_), .B(_07924_), .Y(_07925_));
NAND_g _29584_ (.A(_07915_), .B(_07925_), .Y(_07926_));
AND_g _29585_ (.A(_00012_[4]), .B(_07926_), .Y(_07927_));
NAND_g _29586_ (.A(cpuregs_6[27]), .B(_00012_[2]), .Y(_07928_));
NAND_g _29587_ (.A(cpuregs_2[27]), .B(_11214_), .Y(_07929_));
AND_g _29588_ (.A(_07928_), .B(_07929_), .Y(_07930_));
NAND_g _29589_ (.A(_11212_), .B(_07930_), .Y(_07931_));
NAND_g _29590_ (.A(cpuregs_7[27]), .B(_00012_[2]), .Y(_07932_));
NAND_g _29591_ (.A(cpuregs_3[27]), .B(_11214_), .Y(_07933_));
AND_g _29592_ (.A(_00012_[0]), .B(_07933_), .Y(_07934_));
NAND_g _29593_ (.A(_07932_), .B(_07934_), .Y(_07935_));
AND_g _29594_ (.A(_07931_), .B(_07935_), .Y(_07936_));
NAND_g _29595_ (.A(_11215_), .B(_07936_), .Y(_07937_));
NOR_g _29596_ (.A(cpuregs_10[27]), .B(_00012_[2]), .Y(_07938_));
AND_g _29597_ (.A(_11106_), .B(_00012_[2]), .Y(_07939_));
NOR_g _29598_ (.A(_07938_), .B(_07939_), .Y(_07940_));
NOR_g _29599_ (.A(cpuregs_11[27]), .B(_00012_[2]), .Y(_07941_));
NOT_g _29600_ (.A(_07941_), .Y(_07942_));
NAND_g _29601_ (.A(_11170_), .B(_00012_[2]), .Y(_07943_));
AND_g _29602_ (.A(_00012_[0]), .B(_07943_), .Y(_07944_));
NAND_g _29603_ (.A(_07942_), .B(_07944_), .Y(_07945_));
NAND_g _29604_ (.A(_11212_), .B(_07940_), .Y(_07946_));
NAND_g _29605_ (.A(_07945_), .B(_07946_), .Y(_07947_));
NAND_g _29606_ (.A(_00012_[3]), .B(_07947_), .Y(_07948_));
NAND_g _29607_ (.A(_07937_), .B(_07948_), .Y(_07949_));
AND_g _29608_ (.A(_11216_), .B(_07949_), .Y(_07950_));
NOR_g _29609_ (.A(_07927_), .B(_07950_), .Y(_07951_));
NOR_g _29610_ (.A(_11213_), .B(_07951_), .Y(_07952_));
NAND_g _29611_ (.A(cpuregs_4[27]), .B(_00012_[2]), .Y(_07953_));
NAND_g _29612_ (.A(cpuregs_0[27]), .B(_11214_), .Y(_07954_));
AND_g _29613_ (.A(_11212_), .B(_07954_), .Y(_07955_));
NAND_g _29614_ (.A(_07953_), .B(_07955_), .Y(_07956_));
NAND_g _29615_ (.A(cpuregs_1[27]), .B(_11214_), .Y(_07957_));
NAND_g _29616_ (.A(cpuregs_5[27]), .B(_00012_[2]), .Y(_07958_));
AND_g _29617_ (.A(_00012_[0]), .B(_07958_), .Y(_07959_));
NAND_g _29618_ (.A(_07957_), .B(_07959_), .Y(_07960_));
NOR_g _29619_ (.A(cpuregs_9[27]), .B(_00012_[2]), .Y(_07961_));
NAND_g _29620_ (.A(_11154_), .B(_00012_[2]), .Y(_07962_));
NOR_g _29621_ (.A(cpuregs_8[27]), .B(_00012_[2]), .Y(_07963_));
AND_g _29622_ (.A(_11122_), .B(_00012_[2]), .Y(_07964_));
NOR_g _29623_ (.A(_07963_), .B(_07964_), .Y(_07965_));
NAND_g _29624_ (.A(_07956_), .B(_07960_), .Y(_07966_));
NAND_g _29625_ (.A(_11215_), .B(_07966_), .Y(_07967_));
NAND_g _29626_ (.A(_11212_), .B(_07965_), .Y(_07968_));
NOR_g _29627_ (.A(_11212_), .B(_07961_), .Y(_07969_));
NAND_g _29628_ (.A(_07962_), .B(_07969_), .Y(_07970_));
AND_g _29629_ (.A(_00012_[3]), .B(_07970_), .Y(_07971_));
NAND_g _29630_ (.A(_07968_), .B(_07971_), .Y(_07972_));
AND_g _29631_ (.A(_07967_), .B(_07972_), .Y(_07973_));
NAND_g _29632_ (.A(_11216_), .B(_07973_), .Y(_07974_));
NAND_g _29633_ (.A(cpuregs_25[27]), .B(_00012_[3]), .Y(_07975_));
NAND_g _29634_ (.A(cpuregs_17[27]), .B(_11215_), .Y(_07976_));
NAND_g _29635_ (.A(_07975_), .B(_07976_), .Y(_07977_));
NAND_g _29636_ (.A(_11214_), .B(_07977_), .Y(_07978_));
NAND_g _29637_ (.A(cpuregs_29[27]), .B(_00012_[3]), .Y(_07979_));
NAND_g _29638_ (.A(cpuregs_21[27]), .B(_11215_), .Y(_07980_));
NAND_g _29639_ (.A(_07979_), .B(_07980_), .Y(_07981_));
NAND_g _29640_ (.A(_00012_[2]), .B(_07981_), .Y(_07982_));
AND_g _29641_ (.A(_00012_[0]), .B(_07982_), .Y(_07983_));
NAND_g _29642_ (.A(_07978_), .B(_07983_), .Y(_07984_));
NAND_g _29643_ (.A(cpuregs_24[27]), .B(_00012_[3]), .Y(_07985_));
NAND_g _29644_ (.A(cpuregs_16[27]), .B(_11215_), .Y(_07986_));
NAND_g _29645_ (.A(_07985_), .B(_07986_), .Y(_07987_));
NAND_g _29646_ (.A(_11214_), .B(_07987_), .Y(_07988_));
NAND_g _29647_ (.A(cpuregs_28[27]), .B(_00012_[3]), .Y(_07989_));
NAND_g _29648_ (.A(cpuregs_20[27]), .B(_11215_), .Y(_07990_));
NAND_g _29649_ (.A(_07989_), .B(_07990_), .Y(_07991_));
NAND_g _29650_ (.A(_00012_[2]), .B(_07991_), .Y(_07992_));
AND_g _29651_ (.A(_11212_), .B(_07992_), .Y(_07993_));
NAND_g _29652_ (.A(_07988_), .B(_07993_), .Y(_07994_));
AND_g _29653_ (.A(_00012_[4]), .B(_07994_), .Y(_07995_));
NAND_g _29654_ (.A(_07984_), .B(_07995_), .Y(_07996_));
NAND_g _29655_ (.A(_07974_), .B(_07996_), .Y(_07997_));
AND_g _29656_ (.A(_11213_), .B(_07997_), .Y(_07998_));
NOR_g _29657_ (.A(_07952_), .B(_07998_), .Y(_07999_));
NOR_g _29658_ (.A(_13560_), .B(_07999_), .Y(_08000_));
NAND_g _29659_ (.A(_05765_), .B(_08000_), .Y(_08001_));
AND_g _29660_ (.A(_07905_), .B(_08001_), .Y(_08002_));
AND_g _29661_ (.A(_07894_), .B(_08002_), .Y(_08003_));
NOR_g _29662_ (.A(_07891_), .B(_08003_), .Y(_01234_));
NOR_g _29663_ (.A(pcpi_rs1[28]), .B(_13425_), .Y(_08004_));
NAND_g _29664_ (.A(cpuregs_7[28]), .B(_00012_[2]), .Y(_08005_));
NAND_g _29665_ (.A(cpuregs_3[28]), .B(_11214_), .Y(_08006_));
NAND_g _29666_ (.A(_08005_), .B(_08006_), .Y(_08007_));
AND_g _29667_ (.A(_00012_[0]), .B(_08007_), .Y(_08008_));
NAND_g _29668_ (.A(cpuregs_6[28]), .B(_00012_[2]), .Y(_08009_));
NAND_g _29669_ (.A(cpuregs_2[28]), .B(_11214_), .Y(_08010_));
AND_g _29670_ (.A(_08009_), .B(_08010_), .Y(_08011_));
NOR_g _29671_ (.A(_00012_[0]), .B(_08011_), .Y(_08012_));
NOR_g _29672_ (.A(_08008_), .B(_08012_), .Y(_08013_));
NAND_g _29673_ (.A(cpuregs_5[28]), .B(_00012_[2]), .Y(_08014_));
NAND_g _29674_ (.A(cpuregs_1[28]), .B(_11214_), .Y(_08015_));
NAND_g _29675_ (.A(_08014_), .B(_08015_), .Y(_08016_));
NAND_g _29676_ (.A(_00012_[0]), .B(_08016_), .Y(_08017_));
NAND_g _29677_ (.A(cpuregs_4[28]), .B(_00012_[2]), .Y(_08018_));
NAND_g _29678_ (.A(cpuregs_0[28]), .B(_11214_), .Y(_08019_));
AND_g _29679_ (.A(_08018_), .B(_08019_), .Y(_08020_));
NOR_g _29680_ (.A(_00012_[0]), .B(_08020_), .Y(_08021_));
NAND_g _29681_ (.A(_00012_[1]), .B(_08013_), .Y(_08022_));
NOR_g _29682_ (.A(_00012_[1]), .B(_08021_), .Y(_08023_));
NAND_g _29683_ (.A(_08017_), .B(_08023_), .Y(_08024_));
AND_g _29684_ (.A(_11215_), .B(_08024_), .Y(_08025_));
NAND_g _29685_ (.A(_08022_), .B(_08025_), .Y(_08026_));
NAND_g _29686_ (.A(cpuregs_13[28]), .B(_00012_[0]), .Y(_08027_));
NAND_g _29687_ (.A(cpuregs_12[28]), .B(_11212_), .Y(_08028_));
AND_g _29688_ (.A(_00012_[2]), .B(_08028_), .Y(_08029_));
NAND_g _29689_ (.A(_08027_), .B(_08029_), .Y(_08030_));
NAND_g _29690_ (.A(cpuregs_9[28]), .B(_00012_[0]), .Y(_08031_));
NAND_g _29691_ (.A(cpuregs_8[28]), .B(_11212_), .Y(_08032_));
AND_g _29692_ (.A(_11214_), .B(_08032_), .Y(_08033_));
NAND_g _29693_ (.A(_08031_), .B(_08033_), .Y(_08034_));
AND_g _29694_ (.A(_11213_), .B(_08034_), .Y(_08035_));
NAND_g _29695_ (.A(_08030_), .B(_08035_), .Y(_08036_));
NAND_g _29696_ (.A(cpuregs_15[28]), .B(_00012_[0]), .Y(_08037_));
NAND_g _29697_ (.A(cpuregs_14[28]), .B(_11212_), .Y(_08038_));
AND_g _29698_ (.A(_00012_[2]), .B(_08038_), .Y(_08039_));
NAND_g _29699_ (.A(_08037_), .B(_08039_), .Y(_08040_));
NAND_g _29700_ (.A(cpuregs_11[28]), .B(_00012_[0]), .Y(_08041_));
NAND_g _29701_ (.A(cpuregs_10[28]), .B(_11212_), .Y(_08042_));
AND_g _29702_ (.A(_11214_), .B(_08042_), .Y(_08043_));
NAND_g _29703_ (.A(_08041_), .B(_08043_), .Y(_08044_));
AND_g _29704_ (.A(_00012_[1]), .B(_08044_), .Y(_08045_));
NAND_g _29705_ (.A(_08040_), .B(_08045_), .Y(_08046_));
NAND_g _29706_ (.A(_08036_), .B(_08046_), .Y(_08047_));
NAND_g _29707_ (.A(_00012_[3]), .B(_08047_), .Y(_08048_));
AND_g _29708_ (.A(_08026_), .B(_08048_), .Y(_08049_));
NAND_g _29709_ (.A(_11216_), .B(_08049_), .Y(_08050_));
NAND_g _29710_ (.A(cpuregs_20[28]), .B(_11213_), .Y(_08051_));
NAND_g _29711_ (.A(cpuregs_22[28]), .B(_00012_[1]), .Y(_08052_));
AND_g _29712_ (.A(_00012_[2]), .B(_08052_), .Y(_08053_));
NAND_g _29713_ (.A(_08051_), .B(_08053_), .Y(_08054_));
NAND_g _29714_ (.A(cpuregs_16[28]), .B(_11213_), .Y(_08055_));
NAND_g _29715_ (.A(cpuregs_18[28]), .B(_00012_[1]), .Y(_08056_));
AND_g _29716_ (.A(_11214_), .B(_08056_), .Y(_08057_));
NAND_g _29717_ (.A(_08055_), .B(_08057_), .Y(_08058_));
AND_g _29718_ (.A(_11212_), .B(_08058_), .Y(_08059_));
NAND_g _29719_ (.A(_08054_), .B(_08059_), .Y(_08060_));
NAND_g _29720_ (.A(cpuregs_21[28]), .B(_11213_), .Y(_08061_));
NAND_g _29721_ (.A(cpuregs_23[28]), .B(_00012_[1]), .Y(_08062_));
AND_g _29722_ (.A(_00012_[2]), .B(_08062_), .Y(_08063_));
NAND_g _29723_ (.A(_08061_), .B(_08063_), .Y(_08064_));
NAND_g _29724_ (.A(cpuregs_17[28]), .B(_11213_), .Y(_08065_));
NAND_g _29725_ (.A(cpuregs_19[28]), .B(_00012_[1]), .Y(_08066_));
AND_g _29726_ (.A(_11214_), .B(_08066_), .Y(_08067_));
NAND_g _29727_ (.A(_08065_), .B(_08067_), .Y(_08068_));
AND_g _29728_ (.A(_00012_[0]), .B(_08068_), .Y(_08069_));
NAND_g _29729_ (.A(_08064_), .B(_08069_), .Y(_08070_));
NAND_g _29730_ (.A(_08060_), .B(_08070_), .Y(_08071_));
NAND_g _29731_ (.A(_11215_), .B(_08071_), .Y(_08072_));
NAND_g _29732_ (.A(cpuregs_26[28]), .B(_11214_), .Y(_08073_));
NAND_g _29733_ (.A(cpuregs_30[28]), .B(_00012_[2]), .Y(_08074_));
AND_g _29734_ (.A(_00012_[1]), .B(_08074_), .Y(_08075_));
NAND_g _29735_ (.A(_08073_), .B(_08075_), .Y(_08076_));
NAND_g _29736_ (.A(cpuregs_24[28]), .B(_11214_), .Y(_08077_));
NAND_g _29737_ (.A(cpuregs_28[28]), .B(_00012_[2]), .Y(_08078_));
AND_g _29738_ (.A(_11213_), .B(_08078_), .Y(_08079_));
NAND_g _29739_ (.A(_08077_), .B(_08079_), .Y(_08080_));
AND_g _29740_ (.A(_11212_), .B(_08080_), .Y(_08081_));
NAND_g _29741_ (.A(_08076_), .B(_08081_), .Y(_08082_));
NAND_g _29742_ (.A(cpuregs_27[28]), .B(_11214_), .Y(_08083_));
NAND_g _29743_ (.A(cpuregs_31[28]), .B(_00012_[2]), .Y(_08084_));
AND_g _29744_ (.A(_00012_[1]), .B(_08084_), .Y(_08085_));
NAND_g _29745_ (.A(_08083_), .B(_08085_), .Y(_08086_));
NAND_g _29746_ (.A(cpuregs_29[28]), .B(_00012_[2]), .Y(_08087_));
NAND_g _29747_ (.A(cpuregs_25[28]), .B(_11214_), .Y(_08088_));
AND_g _29748_ (.A(_11213_), .B(_08088_), .Y(_08089_));
NAND_g _29749_ (.A(_08087_), .B(_08089_), .Y(_08090_));
AND_g _29750_ (.A(_00012_[0]), .B(_08090_), .Y(_08091_));
NAND_g _29751_ (.A(_08086_), .B(_08091_), .Y(_08092_));
NAND_g _29752_ (.A(_08082_), .B(_08092_), .Y(_08093_));
NAND_g _29753_ (.A(_00012_[3]), .B(_08093_), .Y(_08094_));
AND_g _29754_ (.A(_00012_[4]), .B(_08072_), .Y(_08095_));
NAND_g _29755_ (.A(_08094_), .B(_08095_), .Y(_08096_));
AND_g _29756_ (.A(_13409_), .B(_08096_), .Y(_08097_));
AND_g _29757_ (.A(_08050_), .B(_08097_), .Y(_08098_));
AND_g _29758_ (.A(_13613_), .B(_08098_), .Y(_08099_));
NAND_g _29759_ (.A(reg_pc[28]), .B(_13714_), .Y(_08100_));
NAND_g _29760_ (.A(pcpi_rs1[31]), .B(_13380_), .Y(_08101_));
AND_g _29761_ (.A(_13383_), .B(_08101_), .Y(_08102_));
NAND_g _29762_ (.A(_07769_), .B(_08102_), .Y(_08103_));
AND_g _29763_ (.A(_13382_), .B(_13707_), .Y(_08104_));
NAND_g _29764_ (.A(_07766_), .B(_08104_), .Y(_08105_));
AND_g _29765_ (.A(_08103_), .B(_08105_), .Y(_08106_));
NAND_g _29766_ (.A(_13389_), .B(_08106_), .Y(_08107_));
AND_g _29767_ (.A(_08100_), .B(_08107_), .Y(_08108_));
NAND_g _29768_ (.A(_13425_), .B(_08108_), .Y(_08109_));
NOR_g _29769_ (.A(_08099_), .B(_08109_), .Y(_08110_));
XOR_g _29770_ (.A(_13438_), .B(_13547_), .Y(_08111_));
NAND_g _29771_ (.A(_13432_), .B(_08111_), .Y(_08112_));
AND_g _29772_ (.A(_08110_), .B(_08112_), .Y(_08113_));
NOR_g _29773_ (.A(_08004_), .B(_08113_), .Y(_01235_));
NOR_g _29774_ (.A(pcpi_rs1[29]), .B(_13425_), .Y(_08114_));
XOR_g _29775_ (.A(decoded_imm[29]), .B(pcpi_rs1[29]), .Y(_08115_));
XNOR_g _29776_ (.A(_13549_), .B(_08115_), .Y(_08116_));
NAND_g _29777_ (.A(_13432_), .B(_08116_), .Y(_08117_));
NAND_g _29778_ (.A(cpuregs_7[29]), .B(_00012_[2]), .Y(_08118_));
NAND_g _29779_ (.A(cpuregs_3[29]), .B(_11214_), .Y(_08119_));
NAND_g _29780_ (.A(_08118_), .B(_08119_), .Y(_08120_));
AND_g _29781_ (.A(_00012_[0]), .B(_08120_), .Y(_08121_));
NAND_g _29782_ (.A(cpuregs_6[29]), .B(_00012_[2]), .Y(_08122_));
NAND_g _29783_ (.A(cpuregs_2[29]), .B(_11214_), .Y(_08123_));
AND_g _29784_ (.A(_08122_), .B(_08123_), .Y(_08124_));
NOR_g _29785_ (.A(_00012_[0]), .B(_08124_), .Y(_08125_));
NOR_g _29786_ (.A(_08121_), .B(_08125_), .Y(_08126_));
NAND_g _29787_ (.A(cpuregs_5[29]), .B(_00012_[2]), .Y(_08127_));
NAND_g _29788_ (.A(cpuregs_1[29]), .B(_11214_), .Y(_08128_));
NAND_g _29789_ (.A(_08127_), .B(_08128_), .Y(_08129_));
NAND_g _29790_ (.A(_00012_[0]), .B(_08129_), .Y(_08130_));
NAND_g _29791_ (.A(cpuregs_4[29]), .B(_00012_[2]), .Y(_08131_));
NAND_g _29792_ (.A(cpuregs_0[29]), .B(_11214_), .Y(_08132_));
AND_g _29793_ (.A(_08131_), .B(_08132_), .Y(_08133_));
NOR_g _29794_ (.A(_00012_[0]), .B(_08133_), .Y(_08134_));
NAND_g _29795_ (.A(_00012_[1]), .B(_08126_), .Y(_08135_));
NOR_g _29796_ (.A(_00012_[1]), .B(_08134_), .Y(_08136_));
NAND_g _29797_ (.A(_08130_), .B(_08136_), .Y(_08137_));
AND_g _29798_ (.A(_11215_), .B(_08137_), .Y(_08138_));
NAND_g _29799_ (.A(_08135_), .B(_08138_), .Y(_08139_));
NAND_g _29800_ (.A(cpuregs_13[29]), .B(_00012_[0]), .Y(_08140_));
NAND_g _29801_ (.A(cpuregs_12[29]), .B(_11212_), .Y(_08141_));
AND_g _29802_ (.A(_00012_[2]), .B(_08141_), .Y(_08142_));
NAND_g _29803_ (.A(_08140_), .B(_08142_), .Y(_08143_));
NAND_g _29804_ (.A(cpuregs_9[29]), .B(_00012_[0]), .Y(_08144_));
NAND_g _29805_ (.A(cpuregs_8[29]), .B(_11212_), .Y(_08145_));
AND_g _29806_ (.A(_11214_), .B(_08145_), .Y(_08146_));
NAND_g _29807_ (.A(_08144_), .B(_08146_), .Y(_08147_));
AND_g _29808_ (.A(_11213_), .B(_08147_), .Y(_08148_));
NAND_g _29809_ (.A(_08143_), .B(_08148_), .Y(_08149_));
NAND_g _29810_ (.A(cpuregs_15[29]), .B(_00012_[0]), .Y(_08150_));
NAND_g _29811_ (.A(cpuregs_14[29]), .B(_11212_), .Y(_08151_));
AND_g _29812_ (.A(_00012_[2]), .B(_08151_), .Y(_08152_));
NAND_g _29813_ (.A(_08150_), .B(_08152_), .Y(_08153_));
NAND_g _29814_ (.A(cpuregs_11[29]), .B(_00012_[0]), .Y(_08154_));
NAND_g _29815_ (.A(cpuregs_10[29]), .B(_11212_), .Y(_08155_));
AND_g _29816_ (.A(_11214_), .B(_08155_), .Y(_08156_));
NAND_g _29817_ (.A(_08154_), .B(_08156_), .Y(_08157_));
AND_g _29818_ (.A(_00012_[1]), .B(_08157_), .Y(_08158_));
NAND_g _29819_ (.A(_08153_), .B(_08158_), .Y(_08159_));
NAND_g _29820_ (.A(_08149_), .B(_08159_), .Y(_08160_));
NAND_g _29821_ (.A(_00012_[3]), .B(_08160_), .Y(_08161_));
AND_g _29822_ (.A(_08139_), .B(_08161_), .Y(_08162_));
NAND_g _29823_ (.A(_11216_), .B(_08162_), .Y(_08163_));
NAND_g _29824_ (.A(_11021_), .B(_00012_[2]), .Y(_08164_));
NOR_g _29825_ (.A(cpuregs_18[29]), .B(_00012_[2]), .Y(_08165_));
NOR_g _29826_ (.A(_00012_[0]), .B(_08165_), .Y(_08166_));
NAND_g _29827_ (.A(_08164_), .B(_08166_), .Y(_08167_));
NAND_g _29828_ (.A(_11190_), .B(_00012_[2]), .Y(_08168_));
NOR_g _29829_ (.A(cpuregs_19[29]), .B(_00012_[2]), .Y(_08169_));
NOR_g _29830_ (.A(_11212_), .B(_08169_), .Y(_08170_));
NAND_g _29831_ (.A(_08168_), .B(_08170_), .Y(_08171_));
AND_g _29832_ (.A(_08167_), .B(_08171_), .Y(_08172_));
NAND_g _29833_ (.A(_11202_), .B(_00012_[2]), .Y(_08173_));
NOR_g _29834_ (.A(cpuregs_16[29]), .B(_00012_[2]), .Y(_08174_));
NOR_g _29835_ (.A(_00012_[0]), .B(_08174_), .Y(_08175_));
NAND_g _29836_ (.A(_08173_), .B(_08175_), .Y(_08176_));
NAND_g _29837_ (.A(_11037_), .B(_00012_[2]), .Y(_08177_));
NOR_g _29838_ (.A(cpuregs_17[29]), .B(_00012_[2]), .Y(_08178_));
NOR_g _29839_ (.A(_11212_), .B(_08178_), .Y(_08179_));
NAND_g _29840_ (.A(_08177_), .B(_08179_), .Y(_08180_));
AND_g _29841_ (.A(_08176_), .B(_08180_), .Y(_08181_));
NAND_g _29842_ (.A(_00012_[1]), .B(_08172_), .Y(_08182_));
NAND_g _29843_ (.A(_11213_), .B(_08181_), .Y(_08183_));
AND_g _29844_ (.A(_08182_), .B(_08183_), .Y(_08184_));
NAND_g _29845_ (.A(_11215_), .B(_08184_), .Y(_08185_));
NAND_g _29846_ (.A(cpuregs_29[29]), .B(_11213_), .Y(_08186_));
NAND_g _29847_ (.A(cpuregs_31[29]), .B(_00012_[1]), .Y(_08187_));
AND_g _29848_ (.A(_00012_[2]), .B(_08187_), .Y(_08188_));
NAND_g _29849_ (.A(_08186_), .B(_08188_), .Y(_08189_));
NAND_g _29850_ (.A(cpuregs_25[29]), .B(_11213_), .Y(_08190_));
NAND_g _29851_ (.A(cpuregs_27[29]), .B(_00012_[1]), .Y(_08191_));
AND_g _29852_ (.A(_11214_), .B(_08191_), .Y(_08192_));
NAND_g _29853_ (.A(_08190_), .B(_08192_), .Y(_08193_));
AND_g _29854_ (.A(_00012_[0]), .B(_08193_), .Y(_08194_));
NAND_g _29855_ (.A(_08189_), .B(_08194_), .Y(_08195_));
NAND_g _29856_ (.A(cpuregs_28[29]), .B(_11213_), .Y(_08196_));
NAND_g _29857_ (.A(cpuregs_30[29]), .B(_00012_[1]), .Y(_08197_));
AND_g _29858_ (.A(_00012_[2]), .B(_08197_), .Y(_08198_));
NAND_g _29859_ (.A(_08196_), .B(_08198_), .Y(_08199_));
NAND_g _29860_ (.A(cpuregs_24[29]), .B(_11213_), .Y(_08200_));
NAND_g _29861_ (.A(cpuregs_26[29]), .B(_00012_[1]), .Y(_08201_));
AND_g _29862_ (.A(_11214_), .B(_08201_), .Y(_08202_));
NAND_g _29863_ (.A(_08200_), .B(_08202_), .Y(_08203_));
AND_g _29864_ (.A(_11212_), .B(_08203_), .Y(_08204_));
NAND_g _29865_ (.A(_08199_), .B(_08204_), .Y(_08205_));
NAND_g _29866_ (.A(_08195_), .B(_08205_), .Y(_08206_));
NAND_g _29867_ (.A(_00012_[3]), .B(_08206_), .Y(_08207_));
AND_g _29868_ (.A(_08185_), .B(_08207_), .Y(_08208_));
NAND_g _29869_ (.A(_00012_[4]), .B(_08208_), .Y(_08209_));
AND_g _29870_ (.A(_13409_), .B(_08209_), .Y(_08210_));
AND_g _29871_ (.A(_08163_), .B(_08210_), .Y(_08211_));
AND_g _29872_ (.A(_13613_), .B(_08211_), .Y(_08212_));
NAND_g _29873_ (.A(reg_pc[29]), .B(_13714_), .Y(_08213_));
NAND_g _29874_ (.A(pcpi_rs1[28]), .B(_13420_), .Y(_08214_));
AND_g _29875_ (.A(_13382_), .B(_08214_), .Y(_08215_));
NAND_g _29876_ (.A(_07879_), .B(_08215_), .Y(_08216_));
NAND_g _29877_ (.A(_07882_), .B(_08102_), .Y(_08217_));
AND_g _29878_ (.A(_08216_), .B(_08217_), .Y(_08218_));
NAND_g _29879_ (.A(_13389_), .B(_08218_), .Y(_08219_));
AND_g _29880_ (.A(_08213_), .B(_08219_), .Y(_08220_));
NAND_g _29881_ (.A(_13425_), .B(_08220_), .Y(_08221_));
NOR_g _29882_ (.A(_08212_), .B(_08221_), .Y(_08222_));
AND_g _29883_ (.A(_08117_), .B(_08222_), .Y(_08223_));
NOR_g _29884_ (.A(_08114_), .B(_08223_), .Y(_01236_));
NOR_g _29885_ (.A(pcpi_rs1[30]), .B(_13425_), .Y(_08224_));
NAND_g _29886_ (.A(cpuregs_8[30]), .B(_11212_), .Y(_08225_));
NAND_g _29887_ (.A(cpuregs_9[30]), .B(_00012_[0]), .Y(_08226_));
NAND_g _29888_ (.A(_08225_), .B(_08226_), .Y(_08227_));
NAND_g _29889_ (.A(_11214_), .B(_08227_), .Y(_08228_));
NAND_g _29890_ (.A(cpuregs_12[30]), .B(_11212_), .Y(_08229_));
NAND_g _29891_ (.A(cpuregs_13[30]), .B(_00012_[0]), .Y(_08230_));
NAND_g _29892_ (.A(_08229_), .B(_08230_), .Y(_08231_));
NAND_g _29893_ (.A(_00012_[2]), .B(_08231_), .Y(_08232_));
AND_g _29894_ (.A(_11213_), .B(_08232_), .Y(_08233_));
NAND_g _29895_ (.A(_08228_), .B(_08233_), .Y(_08234_));
NAND_g _29896_ (.A(cpuregs_10[30]), .B(_11212_), .Y(_08235_));
NAND_g _29897_ (.A(cpuregs_11[30]), .B(_00012_[0]), .Y(_08236_));
NAND_g _29898_ (.A(_08235_), .B(_08236_), .Y(_08237_));
NAND_g _29899_ (.A(_11214_), .B(_08237_), .Y(_08238_));
NAND_g _29900_ (.A(cpuregs_14[30]), .B(_11212_), .Y(_08239_));
NAND_g _29901_ (.A(cpuregs_15[30]), .B(_00012_[0]), .Y(_08240_));
NAND_g _29902_ (.A(_08239_), .B(_08240_), .Y(_08241_));
NAND_g _29903_ (.A(_00012_[2]), .B(_08241_), .Y(_08242_));
AND_g _29904_ (.A(_00012_[1]), .B(_08242_), .Y(_08243_));
NAND_g _29905_ (.A(_08238_), .B(_08243_), .Y(_08244_));
AND_g _29906_ (.A(_08234_), .B(_08244_), .Y(_08245_));
NAND_g _29907_ (.A(cpuregs_1[30]), .B(_11213_), .Y(_08246_));
NAND_g _29908_ (.A(cpuregs_3[30]), .B(_00012_[1]), .Y(_08247_));
AND_g _29909_ (.A(_11214_), .B(_08247_), .Y(_08248_));
NAND_g _29910_ (.A(_08246_), .B(_08248_), .Y(_08249_));
NAND_g _29911_ (.A(cpuregs_5[30]), .B(_11213_), .Y(_08250_));
NAND_g _29912_ (.A(cpuregs_7[30]), .B(_00012_[1]), .Y(_08251_));
AND_g _29913_ (.A(_00012_[2]), .B(_08251_), .Y(_08252_));
NAND_g _29914_ (.A(_08250_), .B(_08252_), .Y(_08253_));
NAND_g _29915_ (.A(_08249_), .B(_08253_), .Y(_08254_));
NAND_g _29916_ (.A(_00012_[0]), .B(_08254_), .Y(_08255_));
NAND_g _29917_ (.A(cpuregs_0[30]), .B(_11213_), .Y(_08256_));
NAND_g _29918_ (.A(cpuregs_2[30]), .B(_00012_[1]), .Y(_08257_));
AND_g _29919_ (.A(_11214_), .B(_08257_), .Y(_08258_));
NAND_g _29920_ (.A(_08256_), .B(_08258_), .Y(_08259_));
NAND_g _29921_ (.A(cpuregs_4[30]), .B(_11213_), .Y(_08260_));
NAND_g _29922_ (.A(cpuregs_6[30]), .B(_00012_[1]), .Y(_08261_));
AND_g _29923_ (.A(_00012_[2]), .B(_08261_), .Y(_08262_));
NAND_g _29924_ (.A(_08260_), .B(_08262_), .Y(_08263_));
NAND_g _29925_ (.A(_08259_), .B(_08263_), .Y(_08264_));
NAND_g _29926_ (.A(_11212_), .B(_08264_), .Y(_08265_));
AND_g _29927_ (.A(_08255_), .B(_08265_), .Y(_08266_));
NAND_g _29928_ (.A(_00012_[3]), .B(_08245_), .Y(_08267_));
NAND_g _29929_ (.A(_11215_), .B(_08266_), .Y(_08268_));
AND_g _29930_ (.A(_11216_), .B(_08268_), .Y(_08269_));
NAND_g _29931_ (.A(_08267_), .B(_08269_), .Y(_08270_));
NAND_g _29932_ (.A(cpuregs_16[30]), .B(_11214_), .Y(_08271_));
NAND_g _29933_ (.A(cpuregs_20[30]), .B(_00012_[2]), .Y(_08272_));
AND_g _29934_ (.A(_08271_), .B(_08272_), .Y(_08273_));
NOR_g _29935_ (.A(_00012_[0]), .B(_08273_), .Y(_08274_));
NAND_g _29936_ (.A(_11038_), .B(_00012_[2]), .Y(_08275_));
NOR_g _29937_ (.A(cpuregs_17[30]), .B(_00012_[2]), .Y(_08276_));
NOR_g _29938_ (.A(_11212_), .B(_08276_), .Y(_08277_));
AND_g _29939_ (.A(_08275_), .B(_08277_), .Y(_08278_));
NOR_g _29940_ (.A(_08274_), .B(_08278_), .Y(_08279_));
NAND_g _29941_ (.A(_11213_), .B(_08279_), .Y(_08280_));
NAND_g _29942_ (.A(cpuregs_22[30]), .B(_00012_[2]), .Y(_08281_));
NAND_g _29943_ (.A(cpuregs_18[30]), .B(_11214_), .Y(_08282_));
NAND_g _29944_ (.A(_08281_), .B(_08282_), .Y(_08283_));
NAND_g _29945_ (.A(_11212_), .B(_08283_), .Y(_08284_));
NOR_g _29946_ (.A(cpuregs_19[30]), .B(_00012_[2]), .Y(_08285_));
NAND_g _29947_ (.A(_11191_), .B(_00012_[2]), .Y(_08286_));
NOR_g _29948_ (.A(_11212_), .B(_08285_), .Y(_08287_));
NAND_g _29949_ (.A(_08286_), .B(_08287_), .Y(_08288_));
AND_g _29950_ (.A(_00012_[1]), .B(_08288_), .Y(_08289_));
NAND_g _29951_ (.A(_08284_), .B(_08289_), .Y(_08290_));
AND_g _29952_ (.A(_08280_), .B(_08290_), .Y(_08291_));
NAND_g _29953_ (.A(cpuregs_27[30]), .B(_00012_[0]), .Y(_08292_));
NAND_g _29954_ (.A(cpuregs_26[30]), .B(_11212_), .Y(_08293_));
AND_g _29955_ (.A(_11214_), .B(_08293_), .Y(_08294_));
NAND_g _29956_ (.A(_08292_), .B(_08294_), .Y(_08295_));
NAND_g _29957_ (.A(cpuregs_31[30]), .B(_00012_[0]), .Y(_08296_));
NAND_g _29958_ (.A(cpuregs_30[30]), .B(_11212_), .Y(_08297_));
AND_g _29959_ (.A(_00012_[2]), .B(_08297_), .Y(_08298_));
NAND_g _29960_ (.A(_08296_), .B(_08298_), .Y(_08299_));
NAND_g _29961_ (.A(_08295_), .B(_08299_), .Y(_08300_));
NAND_g _29962_ (.A(_00012_[1]), .B(_08300_), .Y(_08301_));
NAND_g _29963_ (.A(cpuregs_25[30]), .B(_00012_[0]), .Y(_08302_));
NAND_g _29964_ (.A(cpuregs_24[30]), .B(_11212_), .Y(_08303_));
AND_g _29965_ (.A(_11214_), .B(_08303_), .Y(_08304_));
NAND_g _29966_ (.A(_08302_), .B(_08304_), .Y(_08305_));
NAND_g _29967_ (.A(cpuregs_29[30]), .B(_00012_[0]), .Y(_08306_));
NAND_g _29968_ (.A(cpuregs_28[30]), .B(_11212_), .Y(_08307_));
AND_g _29969_ (.A(_00012_[2]), .B(_08307_), .Y(_08308_));
NAND_g _29970_ (.A(_08306_), .B(_08308_), .Y(_08309_));
NAND_g _29971_ (.A(_08305_), .B(_08309_), .Y(_08310_));
NAND_g _29972_ (.A(_11213_), .B(_08310_), .Y(_08311_));
AND_g _29973_ (.A(_08301_), .B(_08311_), .Y(_08312_));
NAND_g _29974_ (.A(_00012_[3]), .B(_08312_), .Y(_08313_));
NAND_g _29975_ (.A(_11215_), .B(_08291_), .Y(_08314_));
AND_g _29976_ (.A(_00012_[4]), .B(_08314_), .Y(_08315_));
NAND_g _29977_ (.A(_08313_), .B(_08315_), .Y(_08316_));
AND_g _29978_ (.A(_08270_), .B(_08316_), .Y(_08317_));
AND_g _29979_ (.A(_13613_), .B(_08317_), .Y(_08318_));
NAND_g _29980_ (.A(_13409_), .B(_08318_), .Y(_08319_));
NAND_g _29981_ (.A(reg_pc[30]), .B(_13714_), .Y(_08320_));
NAND_g _29982_ (.A(_07899_), .B(_08102_), .Y(_08321_));
NAND_g _29983_ (.A(pcpi_rs1[29]), .B(_13420_), .Y(_08322_));
AND_g _29984_ (.A(_07896_), .B(_08322_), .Y(_08323_));
NAND_g _29985_ (.A(_13382_), .B(_08323_), .Y(_08324_));
AND_g _29986_ (.A(_08321_), .B(_08324_), .Y(_08325_));
NAND_g _29987_ (.A(_13389_), .B(_08325_), .Y(_08326_));
AND_g _29988_ (.A(_08320_), .B(_08326_), .Y(_08327_));
AND_g _29989_ (.A(_13425_), .B(_08327_), .Y(_08328_));
AND_g _29990_ (.A(_08319_), .B(_08328_), .Y(_08329_));
XOR_g _29991_ (.A(_13434_), .B(_13551_), .Y(_08330_));
NAND_g _29992_ (.A(_13432_), .B(_08330_), .Y(_08331_));
AND_g _29993_ (.A(_08329_), .B(_08331_), .Y(_08332_));
NOR_g _29994_ (.A(_08224_), .B(_08332_), .Y(_01237_));
NAND_g _29995_ (.A(_11918_), .B(_00798_), .Y(_08333_));
NAND_g _29996_ (.A(decoded_imm_j[6]), .B(_11919_), .Y(_08334_));
NAND_g _29997_ (.A(_08333_), .B(_08334_), .Y(_01270_));
NAND_g _29998_ (.A(_11918_), .B(_00799_), .Y(_08335_));
NAND_g _29999_ (.A(decoded_imm_j[7]), .B(_11919_), .Y(_08336_));
NAND_g _30000_ (.A(_08335_), .B(_08336_), .Y(_01271_));
NAND_g _30001_ (.A(_11918_), .B(_00802_), .Y(_08337_));
NAND_g _30002_ (.A(decoded_imm_j[10]), .B(_11919_), .Y(_08338_));
NAND_g _30003_ (.A(_08337_), .B(_08338_), .Y(_01272_));
NAND_g _30004_ (.A(_11918_), .B(_00796_), .Y(_08339_));
NAND_g _30005_ (.A(decoded_imm_j[4]), .B(_11919_), .Y(_08340_));
NAND_g _30006_ (.A(_08339_), .B(_08340_), .Y(_01273_));
NAND_g _30007_ (.A(_11918_), .B(_00803_), .Y(_08341_));
NAND_g _30008_ (.A(decoded_imm_j[31]), .B(_11919_), .Y(_08342_));
NAND_g _30009_ (.A(_08341_), .B(_08342_), .Y(_01274_));
AND_g _30010_ (.A(_11289_), .B(_04426_), .Y(_08343_));
NAND_g _30011_ (.A(_11289_), .B(_04426_), .Y(_08344_));
NAND_g _30012_ (.A(cpuregs_13[0]), .B(_08344_), .Y(_08345_));
NAND_g _30013_ (.A(_11301_), .B(_08343_), .Y(_08346_));
NAND_g _30014_ (.A(_08345_), .B(_08346_), .Y(_01275_));
NAND_g _30015_ (.A(cpuregs_13[1]), .B(_08344_), .Y(_08347_));
NAND_g _30016_ (.A(_11310_), .B(_08343_), .Y(_08348_));
NAND_g _30017_ (.A(_08347_), .B(_08348_), .Y(_01276_));
NAND_g _30018_ (.A(cpuregs_13[2]), .B(_08344_), .Y(_08349_));
NAND_g _30019_ (.A(_11319_), .B(_08343_), .Y(_08350_));
NAND_g _30020_ (.A(_08349_), .B(_08350_), .Y(_01277_));
NAND_g _30021_ (.A(cpuregs_13[3]), .B(_08344_), .Y(_08351_));
NAND_g _30022_ (.A(_11332_), .B(_08343_), .Y(_08352_));
NAND_g _30023_ (.A(_08351_), .B(_08352_), .Y(_01278_));
NAND_g _30024_ (.A(cpuregs_13[4]), .B(_08344_), .Y(_08353_));
NAND_g _30025_ (.A(_11345_), .B(_08343_), .Y(_08354_));
NAND_g _30026_ (.A(_08353_), .B(_08354_), .Y(_01279_));
NAND_g _30027_ (.A(cpuregs_13[5]), .B(_08344_), .Y(_08355_));
NAND_g _30028_ (.A(_11358_), .B(_08343_), .Y(_08356_));
NAND_g _30029_ (.A(_08355_), .B(_08356_), .Y(_01280_));
NAND_g _30030_ (.A(cpuregs_13[6]), .B(_08344_), .Y(_08357_));
NAND_g _30031_ (.A(_11371_), .B(_08343_), .Y(_08358_));
NAND_g _30032_ (.A(_08357_), .B(_08358_), .Y(_01281_));
NAND_g _30033_ (.A(cpuregs_13[7]), .B(_08344_), .Y(_08359_));
NAND_g _30034_ (.A(_11384_), .B(_08343_), .Y(_08360_));
NAND_g _30035_ (.A(_08359_), .B(_08360_), .Y(_01282_));
NAND_g _30036_ (.A(cpuregs_13[8]), .B(_08344_), .Y(_08361_));
NAND_g _30037_ (.A(_11397_), .B(_08343_), .Y(_08362_));
NAND_g _30038_ (.A(_08361_), .B(_08362_), .Y(_01283_));
NAND_g _30039_ (.A(cpuregs_13[9]), .B(_08344_), .Y(_08363_));
NAND_g _30040_ (.A(_11410_), .B(_08343_), .Y(_08364_));
NAND_g _30041_ (.A(_08363_), .B(_08364_), .Y(_01284_));
NAND_g _30042_ (.A(cpuregs_13[10]), .B(_08344_), .Y(_08365_));
NAND_g _30043_ (.A(_11423_), .B(_08343_), .Y(_08366_));
NAND_g _30044_ (.A(_08365_), .B(_08366_), .Y(_01285_));
NAND_g _30045_ (.A(cpuregs_13[11]), .B(_08344_), .Y(_08367_));
NAND_g _30046_ (.A(_11436_), .B(_08343_), .Y(_08368_));
NAND_g _30047_ (.A(_08367_), .B(_08368_), .Y(_01286_));
NAND_g _30048_ (.A(cpuregs_13[12]), .B(_08344_), .Y(_08369_));
NAND_g _30049_ (.A(_11449_), .B(_08343_), .Y(_08370_));
NAND_g _30050_ (.A(_08369_), .B(_08370_), .Y(_01287_));
NAND_g _30051_ (.A(cpuregs_13[13]), .B(_08344_), .Y(_08371_));
NAND_g _30052_ (.A(_11462_), .B(_08343_), .Y(_08372_));
NAND_g _30053_ (.A(_08371_), .B(_08372_), .Y(_01288_));
NAND_g _30054_ (.A(cpuregs_13[14]), .B(_08344_), .Y(_08373_));
NAND_g _30055_ (.A(_11475_), .B(_08343_), .Y(_08374_));
NAND_g _30056_ (.A(_08373_), .B(_08374_), .Y(_01289_));
NAND_g _30057_ (.A(cpuregs_13[15]), .B(_08344_), .Y(_08375_));
NAND_g _30058_ (.A(_11488_), .B(_08343_), .Y(_08376_));
NAND_g _30059_ (.A(_08375_), .B(_08376_), .Y(_01290_));
NAND_g _30060_ (.A(cpuregs_13[16]), .B(_08344_), .Y(_08377_));
NAND_g _30061_ (.A(_11501_), .B(_08343_), .Y(_08378_));
NAND_g _30062_ (.A(_08377_), .B(_08378_), .Y(_01291_));
NAND_g _30063_ (.A(cpuregs_13[17]), .B(_08344_), .Y(_08379_));
NAND_g _30064_ (.A(_11514_), .B(_08343_), .Y(_08380_));
NAND_g _30065_ (.A(_08379_), .B(_08380_), .Y(_01292_));
NAND_g _30066_ (.A(cpuregs_13[18]), .B(_08344_), .Y(_08381_));
NAND_g _30067_ (.A(_11527_), .B(_08343_), .Y(_08382_));
NAND_g _30068_ (.A(_08381_), .B(_08382_), .Y(_01293_));
NAND_g _30069_ (.A(cpuregs_13[19]), .B(_08344_), .Y(_08383_));
NAND_g _30070_ (.A(_11540_), .B(_08343_), .Y(_08384_));
NAND_g _30071_ (.A(_08383_), .B(_08384_), .Y(_01294_));
NAND_g _30072_ (.A(cpuregs_13[20]), .B(_08344_), .Y(_08385_));
NAND_g _30073_ (.A(_11553_), .B(_08343_), .Y(_08386_));
NAND_g _30074_ (.A(_08385_), .B(_08386_), .Y(_01295_));
NAND_g _30075_ (.A(cpuregs_13[21]), .B(_08344_), .Y(_08387_));
NAND_g _30076_ (.A(_11566_), .B(_08343_), .Y(_08388_));
NAND_g _30077_ (.A(_08387_), .B(_08388_), .Y(_01296_));
NAND_g _30078_ (.A(cpuregs_13[22]), .B(_08344_), .Y(_08389_));
NAND_g _30079_ (.A(_11579_), .B(_08343_), .Y(_08390_));
NAND_g _30080_ (.A(_08389_), .B(_08390_), .Y(_01297_));
NAND_g _30081_ (.A(cpuregs_13[23]), .B(_08344_), .Y(_08391_));
NAND_g _30082_ (.A(_11592_), .B(_08343_), .Y(_08392_));
NAND_g _30083_ (.A(_08391_), .B(_08392_), .Y(_01298_));
NAND_g _30084_ (.A(cpuregs_13[24]), .B(_08344_), .Y(_08393_));
NAND_g _30085_ (.A(_11605_), .B(_08343_), .Y(_08394_));
NAND_g _30086_ (.A(_08393_), .B(_08394_), .Y(_01299_));
NAND_g _30087_ (.A(cpuregs_13[25]), .B(_08344_), .Y(_08395_));
NAND_g _30088_ (.A(_11618_), .B(_08343_), .Y(_08396_));
NAND_g _30089_ (.A(_08395_), .B(_08396_), .Y(_01300_));
NAND_g _30090_ (.A(cpuregs_13[26]), .B(_08344_), .Y(_08397_));
NAND_g _30091_ (.A(_11631_), .B(_08343_), .Y(_08398_));
NAND_g _30092_ (.A(_08397_), .B(_08398_), .Y(_01301_));
NAND_g _30093_ (.A(cpuregs_13[27]), .B(_08344_), .Y(_08399_));
NAND_g _30094_ (.A(_11644_), .B(_08343_), .Y(_08400_));
NAND_g _30095_ (.A(_08399_), .B(_08400_), .Y(_01302_));
NAND_g _30096_ (.A(cpuregs_13[28]), .B(_08344_), .Y(_08401_));
NAND_g _30097_ (.A(_11657_), .B(_08343_), .Y(_08402_));
NAND_g _30098_ (.A(_08401_), .B(_08402_), .Y(_01303_));
NAND_g _30099_ (.A(cpuregs_13[29]), .B(_08344_), .Y(_08403_));
NAND_g _30100_ (.A(_11670_), .B(_08343_), .Y(_08404_));
NAND_g _30101_ (.A(_08403_), .B(_08404_), .Y(_01304_));
NAND_g _30102_ (.A(cpuregs_13[30]), .B(_08344_), .Y(_08405_));
NAND_g _30103_ (.A(_11683_), .B(_08343_), .Y(_08406_));
NAND_g _30104_ (.A(_08405_), .B(_08406_), .Y(_01305_));
NAND_g _30105_ (.A(cpuregs_13[31]), .B(_08344_), .Y(_08407_));
NAND_g _30106_ (.A(_11695_), .B(_08343_), .Y(_08408_));
NAND_g _30107_ (.A(_08407_), .B(_08408_), .Y(_01306_));
NAND_g _30108_ (.A(decoded_imm_j[12]), .B(_11919_), .Y(_08409_));
NAND_g _30109_ (.A(_11918_), .B(_00784_), .Y(_08410_));
NAND_g _30110_ (.A(_08409_), .B(_08410_), .Y(_01307_));
NAND_g _30111_ (.A(_11918_), .B(_00785_), .Y(_08411_));
NAND_g _30112_ (.A(decoded_imm_j[13]), .B(_11919_), .Y(_08412_));
NAND_g _30113_ (.A(_08411_), .B(_08412_), .Y(_01308_));
NOR_g _30114_ (.A(decoded_imm_j[14]), .B(_11918_), .Y(_08413_));
NOR_g _30115_ (.A(_12273_), .B(_08413_), .Y(_01309_));
NAND_g _30116_ (.A(_11918_), .B(_00790_), .Y(_08414_));
NAND_g _30117_ (.A(decoded_imm_j[18]), .B(_11919_), .Y(_08415_));
NAND_g _30118_ (.A(_08414_), .B(_08415_), .Y(_01310_));
NAND_g _30119_ (.A(_11918_), .B(_00791_), .Y(_08416_));
NAND_g _30120_ (.A(decoded_imm_j[19]), .B(_11919_), .Y(_08417_));
NAND_g _30121_ (.A(_08416_), .B(_08417_), .Y(_01311_));
NAND_g _30122_ (.A(_11918_), .B(_00787_), .Y(_08418_));
NAND_g _30123_ (.A(decoded_imm_j[15]), .B(_11919_), .Y(_08419_));
NAND_g _30124_ (.A(_08418_), .B(_08419_), .Y(_01312_));
NAND_g _30125_ (.A(_11918_), .B(_00788_), .Y(_08420_));
NAND_g _30126_ (.A(decoded_imm_j[16]), .B(_11919_), .Y(_08421_));
NAND_g _30127_ (.A(_08420_), .B(_08421_), .Y(_01313_));
NAND_g _30128_ (.A(_11918_), .B(_00789_), .Y(_08422_));
NAND_g _30129_ (.A(decoded_imm_j[17]), .B(_11919_), .Y(_08423_));
NAND_g _30130_ (.A(_08422_), .B(_08423_), .Y(_01314_));
AND_g _30131_ (.A(_11932_), .B(_04426_), .Y(_08424_));
NAND_g _30132_ (.A(_11932_), .B(_04426_), .Y(_08425_));
NAND_g _30133_ (.A(cpuregs_15[0]), .B(_08425_), .Y(_08426_));
NAND_g _30134_ (.A(_11301_), .B(_08424_), .Y(_08427_));
NAND_g _30135_ (.A(_08426_), .B(_08427_), .Y(_01315_));
NAND_g _30136_ (.A(cpuregs_15[1]), .B(_08425_), .Y(_08428_));
NAND_g _30137_ (.A(_11310_), .B(_08424_), .Y(_08429_));
NAND_g _30138_ (.A(_08428_), .B(_08429_), .Y(_01316_));
NAND_g _30139_ (.A(cpuregs_15[2]), .B(_08425_), .Y(_08430_));
NAND_g _30140_ (.A(_11319_), .B(_08424_), .Y(_08431_));
NAND_g _30141_ (.A(_08430_), .B(_08431_), .Y(_01317_));
NAND_g _30142_ (.A(cpuregs_15[3]), .B(_08425_), .Y(_08432_));
NAND_g _30143_ (.A(_11332_), .B(_08424_), .Y(_08433_));
NAND_g _30144_ (.A(_08432_), .B(_08433_), .Y(_01318_));
NAND_g _30145_ (.A(cpuregs_15[4]), .B(_08425_), .Y(_08434_));
NAND_g _30146_ (.A(_11345_), .B(_08424_), .Y(_08435_));
NAND_g _30147_ (.A(_08434_), .B(_08435_), .Y(_01319_));
NAND_g _30148_ (.A(cpuregs_15[5]), .B(_08425_), .Y(_08436_));
NAND_g _30149_ (.A(_11358_), .B(_08424_), .Y(_08437_));
NAND_g _30150_ (.A(_08436_), .B(_08437_), .Y(_01320_));
NAND_g _30151_ (.A(cpuregs_15[6]), .B(_08425_), .Y(_08438_));
NAND_g _30152_ (.A(_11371_), .B(_08424_), .Y(_08439_));
NAND_g _30153_ (.A(_08438_), .B(_08439_), .Y(_01321_));
NAND_g _30154_ (.A(cpuregs_15[7]), .B(_08425_), .Y(_08440_));
NAND_g _30155_ (.A(_11384_), .B(_08424_), .Y(_08441_));
NAND_g _30156_ (.A(_08440_), .B(_08441_), .Y(_01322_));
NAND_g _30157_ (.A(cpuregs_15[8]), .B(_08425_), .Y(_08442_));
NAND_g _30158_ (.A(_11397_), .B(_08424_), .Y(_08443_));
NAND_g _30159_ (.A(_08442_), .B(_08443_), .Y(_01323_));
NAND_g _30160_ (.A(cpuregs_15[9]), .B(_08425_), .Y(_08444_));
NAND_g _30161_ (.A(_11410_), .B(_08424_), .Y(_08445_));
NAND_g _30162_ (.A(_08444_), .B(_08445_), .Y(_01324_));
NAND_g _30163_ (.A(cpuregs_15[10]), .B(_08425_), .Y(_08446_));
NAND_g _30164_ (.A(_11423_), .B(_08424_), .Y(_08447_));
NAND_g _30165_ (.A(_08446_), .B(_08447_), .Y(_01325_));
NAND_g _30166_ (.A(cpuregs_15[11]), .B(_08425_), .Y(_08448_));
NAND_g _30167_ (.A(_11436_), .B(_08424_), .Y(_08449_));
NAND_g _30168_ (.A(_08448_), .B(_08449_), .Y(_01326_));
NAND_g _30169_ (.A(cpuregs_15[12]), .B(_08425_), .Y(_08450_));
NAND_g _30170_ (.A(_11449_), .B(_08424_), .Y(_08451_));
NAND_g _30171_ (.A(_08450_), .B(_08451_), .Y(_01327_));
NAND_g _30172_ (.A(cpuregs_15[13]), .B(_08425_), .Y(_08452_));
NAND_g _30173_ (.A(_11462_), .B(_08424_), .Y(_08453_));
NAND_g _30174_ (.A(_08452_), .B(_08453_), .Y(_01328_));
NAND_g _30175_ (.A(cpuregs_15[14]), .B(_08425_), .Y(_08454_));
NAND_g _30176_ (.A(_11475_), .B(_08424_), .Y(_08455_));
NAND_g _30177_ (.A(_08454_), .B(_08455_), .Y(_01329_));
NAND_g _30178_ (.A(cpuregs_15[15]), .B(_08425_), .Y(_08456_));
NAND_g _30179_ (.A(_11488_), .B(_08424_), .Y(_08457_));
NAND_g _30180_ (.A(_08456_), .B(_08457_), .Y(_01330_));
NAND_g _30181_ (.A(cpuregs_15[16]), .B(_08425_), .Y(_08458_));
NAND_g _30182_ (.A(_11501_), .B(_08424_), .Y(_08459_));
NAND_g _30183_ (.A(_08458_), .B(_08459_), .Y(_01331_));
NAND_g _30184_ (.A(_11514_), .B(_08424_), .Y(_08460_));
NAND_g _30185_ (.A(cpuregs_15[17]), .B(_08425_), .Y(_08461_));
NAND_g _30186_ (.A(_08460_), .B(_08461_), .Y(_01332_));
NAND_g _30187_ (.A(_11527_), .B(_08424_), .Y(_08462_));
NAND_g _30188_ (.A(cpuregs_15[18]), .B(_08425_), .Y(_08463_));
NAND_g _30189_ (.A(_08462_), .B(_08463_), .Y(_01333_));
NAND_g _30190_ (.A(_11540_), .B(_08424_), .Y(_08464_));
NAND_g _30191_ (.A(cpuregs_15[19]), .B(_08425_), .Y(_08465_));
NAND_g _30192_ (.A(_08464_), .B(_08465_), .Y(_01334_));
NAND_g _30193_ (.A(_11553_), .B(_08424_), .Y(_08466_));
NAND_g _30194_ (.A(cpuregs_15[20]), .B(_08425_), .Y(_08467_));
NAND_g _30195_ (.A(_08466_), .B(_08467_), .Y(_01335_));
NAND_g _30196_ (.A(_11566_), .B(_08424_), .Y(_08468_));
NAND_g _30197_ (.A(cpuregs_15[21]), .B(_08425_), .Y(_08469_));
NAND_g _30198_ (.A(_08468_), .B(_08469_), .Y(_01336_));
NAND_g _30199_ (.A(_11579_), .B(_08424_), .Y(_08470_));
NAND_g _30200_ (.A(cpuregs_15[22]), .B(_08425_), .Y(_08471_));
NAND_g _30201_ (.A(_08470_), .B(_08471_), .Y(_01337_));
NAND_g _30202_ (.A(_11592_), .B(_08424_), .Y(_08472_));
NAND_g _30203_ (.A(cpuregs_15[23]), .B(_08425_), .Y(_08473_));
NAND_g _30204_ (.A(_08472_), .B(_08473_), .Y(_01338_));
NAND_g _30205_ (.A(_11605_), .B(_08424_), .Y(_08474_));
NAND_g _30206_ (.A(cpuregs_15[24]), .B(_08425_), .Y(_08475_));
NAND_g _30207_ (.A(_08474_), .B(_08475_), .Y(_01339_));
NAND_g _30208_ (.A(_11618_), .B(_08424_), .Y(_08476_));
NAND_g _30209_ (.A(cpuregs_15[25]), .B(_08425_), .Y(_08477_));
NAND_g _30210_ (.A(_08476_), .B(_08477_), .Y(_01340_));
NAND_g _30211_ (.A(_11631_), .B(_08424_), .Y(_08478_));
NAND_g _30212_ (.A(cpuregs_15[26]), .B(_08425_), .Y(_08479_));
NAND_g _30213_ (.A(_08478_), .B(_08479_), .Y(_01341_));
NAND_g _30214_ (.A(_11644_), .B(_08424_), .Y(_08480_));
NAND_g _30215_ (.A(cpuregs_15[27]), .B(_08425_), .Y(_08481_));
NAND_g _30216_ (.A(_08480_), .B(_08481_), .Y(_01342_));
NAND_g _30217_ (.A(_11657_), .B(_08424_), .Y(_08482_));
NAND_g _30218_ (.A(cpuregs_15[28]), .B(_08425_), .Y(_08483_));
NAND_g _30219_ (.A(_08482_), .B(_08483_), .Y(_01343_));
NAND_g _30220_ (.A(_11670_), .B(_08424_), .Y(_08484_));
NAND_g _30221_ (.A(cpuregs_15[29]), .B(_08425_), .Y(_08485_));
NAND_g _30222_ (.A(_08484_), .B(_08485_), .Y(_01344_));
NAND_g _30223_ (.A(_11683_), .B(_08424_), .Y(_08486_));
NAND_g _30224_ (.A(cpuregs_15[30]), .B(_08425_), .Y(_08487_));
NAND_g _30225_ (.A(_08486_), .B(_08487_), .Y(_01345_));
NAND_g _30226_ (.A(_11695_), .B(_08424_), .Y(_08488_));
NAND_g _30227_ (.A(cpuregs_15[31]), .B(_08425_), .Y(_08489_));
NAND_g _30228_ (.A(_08488_), .B(_08489_), .Y(_01346_));
NAND_g _30229_ (.A(count_instr[0]), .B(launch_next_insn), .Y(_08490_));
NOR_g _30230_ (.A(count_instr[0]), .B(launch_next_insn), .Y(_08491_));
NOR_g _30231_ (.A(_10963_), .B(_08491_), .Y(_08492_));
AND_g _30232_ (.A(_08490_), .B(_08492_), .Y(_01347_));
NAND_g _30233_ (.A(_10892_), .B(_08490_), .Y(_08493_));
NAND_g _30234_ (.A(resetn), .B(_08493_), .Y(_08494_));
NOR_g _30235_ (.A(_10892_), .B(_08490_), .Y(_08495_));
AND_g _30236_ (.A(count_instr[1]), .B(count_instr[0]), .Y(_08496_));
NOR_g _30237_ (.A(_08494_), .B(_08495_), .Y(_01348_));
NOR_g _30238_ (.A(count_instr[2]), .B(_08495_), .Y(_08497_));
NOR_g _30239_ (.A(_10963_), .B(_08497_), .Y(_08498_));
NAND_g _30240_ (.A(count_instr[2]), .B(_08495_), .Y(_08499_));
AND_g _30241_ (.A(_08498_), .B(_08499_), .Y(_01349_));
NAND_g _30242_ (.A(_10891_), .B(_08499_), .Y(_08500_));
AND_g _30243_ (.A(count_instr[3]), .B(count_instr[2]), .Y(_08501_));
AND_g _30244_ (.A(_08495_), .B(_08501_), .Y(_08502_));
NAND_g _30245_ (.A(resetn), .B(_08500_), .Y(_08503_));
AND_g _30246_ (.A(count_instr[3]), .B(_08496_), .Y(_08504_));
AND_g _30247_ (.A(count_instr[2]), .B(_08504_), .Y(_08505_));
AND_g _30248_ (.A(launch_next_insn), .B(_08505_), .Y(_08506_));
NOR_g _30249_ (.A(_08503_), .B(_08506_), .Y(_01350_));
NOR_g _30250_ (.A(count_instr[4]), .B(_08506_), .Y(_08507_));
NOR_g _30251_ (.A(_10963_), .B(_08507_), .Y(_08508_));
NAND_g _30252_ (.A(count_instr[4]), .B(_08506_), .Y(_08509_));
AND_g _30253_ (.A(_08508_), .B(_08509_), .Y(_01351_));
NAND_g _30254_ (.A(_10890_), .B(_08509_), .Y(_08510_));
AND_g _30255_ (.A(count_instr[5]), .B(count_instr[4]), .Y(_08511_));
AND_g _30256_ (.A(_08502_), .B(_08511_), .Y(_08512_));
NAND_g _30257_ (.A(_08502_), .B(_08511_), .Y(_08513_));
NAND_g _30258_ (.A(resetn), .B(_08510_), .Y(_08514_));
NOR_g _30259_ (.A(_10890_), .B(_08509_), .Y(_08515_));
NOR_g _30260_ (.A(_08514_), .B(_08515_), .Y(_01352_));
NAND_g _30261_ (.A(_10889_), .B(_08513_), .Y(_08516_));
AND_g _30262_ (.A(resetn), .B(_08516_), .Y(_08517_));
NAND_g _30263_ (.A(count_instr[6]), .B(_08515_), .Y(_08518_));
AND_g _30264_ (.A(_08517_), .B(_08518_), .Y(_01353_));
NAND_g _30265_ (.A(_10888_), .B(_08518_), .Y(_08519_));
AND_g _30266_ (.A(count_instr[7]), .B(count_instr[6]), .Y(_08520_));
AND_g _30267_ (.A(_08512_), .B(_08520_), .Y(_08521_));
NAND_g _30268_ (.A(resetn), .B(_08519_), .Y(_08522_));
NOR_g _30269_ (.A(_10888_), .B(_08518_), .Y(_08523_));
NOR_g _30270_ (.A(_08522_), .B(_08523_), .Y(_01354_));
NOR_g _30271_ (.A(count_instr[8]), .B(_08521_), .Y(_08524_));
NOR_g _30272_ (.A(_10963_), .B(_08524_), .Y(_08525_));
NAND_g _30273_ (.A(count_instr[8]), .B(_08523_), .Y(_08526_));
AND_g _30274_ (.A(_08525_), .B(_08526_), .Y(_01355_));
NAND_g _30275_ (.A(_10887_), .B(_08526_), .Y(_08527_));
AND_g _30276_ (.A(count_instr[9]), .B(count_instr[8]), .Y(_08528_));
AND_g _30277_ (.A(_08521_), .B(_08528_), .Y(_08529_));
NOR_g _30278_ (.A(_10963_), .B(_08529_), .Y(_08530_));
AND_g _30279_ (.A(_08527_), .B(_08530_), .Y(_01356_));
NOR_g _30280_ (.A(count_instr[10]), .B(_08529_), .Y(_08531_));
NOR_g _30281_ (.A(_10963_), .B(_08531_), .Y(_08532_));
NAND_g _30282_ (.A(count_instr[10]), .B(_08529_), .Y(_08533_));
NOT_g _30283_ (.A(_08533_), .Y(_08534_));
AND_g _30284_ (.A(_08532_), .B(_08533_), .Y(_01357_));
NAND_g _30285_ (.A(_10886_), .B(_08533_), .Y(_08535_));
AND_g _30286_ (.A(resetn), .B(_08535_), .Y(_08536_));
NAND_g _30287_ (.A(count_instr[11]), .B(_08534_), .Y(_08537_));
NOT_g _30288_ (.A(_08537_), .Y(_08538_));
AND_g _30289_ (.A(count_instr[11]), .B(_08528_), .Y(_08539_));
AND_g _30290_ (.A(count_instr[10]), .B(_08539_), .Y(_08540_));
AND_g _30291_ (.A(_08536_), .B(_08537_), .Y(_01358_));
NAND_g _30292_ (.A(_10885_), .B(_08537_), .Y(_08541_));
AND_g _30293_ (.A(resetn), .B(_08541_), .Y(_08542_));
NAND_g _30294_ (.A(count_instr[12]), .B(_08538_), .Y(_08543_));
AND_g _30295_ (.A(_08542_), .B(_08543_), .Y(_01359_));
XNOR_g _30296_ (.A(count_instr[13]), .B(_08543_), .Y(_08544_));
AND_g _30297_ (.A(resetn), .B(_08544_), .Y(_01360_));
AND_g _30298_ (.A(count_instr[13]), .B(count_instr[12]), .Y(_08545_));
AND_g _30299_ (.A(count_instr[11]), .B(count_instr[10]), .Y(_08546_));
AND_g _30300_ (.A(_08545_), .B(_08546_), .Y(_08547_));
AND_g _30301_ (.A(_08528_), .B(_08547_), .Y(_08548_));
AND_g _30302_ (.A(_08521_), .B(_08548_), .Y(_08549_));
AND_g _30303_ (.A(count_instr[12]), .B(count_instr[5]), .Y(_08550_));
AND_g _30304_ (.A(count_instr[13]), .B(count_instr[4]), .Y(_08551_));
AND_g _30305_ (.A(_08520_), .B(_08551_), .Y(_08552_));
AND_g _30306_ (.A(_08550_), .B(_08552_), .Y(_08553_));
AND_g _30307_ (.A(_08540_), .B(_08553_), .Y(_08554_));
AND_g _30308_ (.A(_08506_), .B(_08554_), .Y(_08555_));
AND_g _30309_ (.A(_08520_), .B(_08545_), .Y(_08556_));
AND_g _30310_ (.A(_08511_), .B(_08556_), .Y(_08557_));
AND_g _30311_ (.A(_08540_), .B(_08557_), .Y(_08558_));
AND_g _30312_ (.A(_08505_), .B(_08558_), .Y(_08559_));
AND_g _30313_ (.A(launch_next_insn), .B(_08559_), .Y(_08560_));
NOR_g _30314_ (.A(count_instr[14]), .B(_08560_), .Y(_08561_));
NOR_g _30315_ (.A(_10963_), .B(_08561_), .Y(_08562_));
AND_g _30316_ (.A(count_instr[14]), .B(_08555_), .Y(_08563_));
NAND_g _30317_ (.A(count_instr[14]), .B(_08560_), .Y(_08564_));
AND_g _30318_ (.A(_08562_), .B(_08564_), .Y(_01361_));
NAND_g _30319_ (.A(_10884_), .B(_08564_), .Y(_08565_));
AND_g _30320_ (.A(count_instr[15]), .B(count_instr[14]), .Y(_08566_));
AND_g _30321_ (.A(resetn), .B(_08565_), .Y(_08567_));
NAND_g _30322_ (.A(count_instr[15]), .B(_08563_), .Y(_08568_));
AND_g _30323_ (.A(_08567_), .B(_08568_), .Y(_01362_));
NAND_g _30324_ (.A(_10883_), .B(_08568_), .Y(_08569_));
NAND_g _30325_ (.A(resetn), .B(_08569_), .Y(_08570_));
NOR_g _30326_ (.A(_10883_), .B(_08568_), .Y(_08571_));
AND_g _30327_ (.A(count_instr[16]), .B(_08566_), .Y(_08572_));
AND_g _30328_ (.A(_08560_), .B(_08572_), .Y(_08573_));
NOR_g _30329_ (.A(_08570_), .B(_08573_), .Y(_01363_));
NOR_g _30330_ (.A(count_instr[17]), .B(_08573_), .Y(_08574_));
AND_g _30331_ (.A(count_instr[17]), .B(count_instr[16]), .Y(_08575_));
AND_g _30332_ (.A(_08566_), .B(_08575_), .Y(_08576_));
AND_g _30333_ (.A(_08549_), .B(_08576_), .Y(_08577_));
NAND_g _30334_ (.A(_08549_), .B(_08576_), .Y(_08578_));
NAND_g _30335_ (.A(resetn), .B(_08578_), .Y(_08579_));
NAND_g _30336_ (.A(count_instr[17]), .B(_08571_), .Y(_08580_));
NOR_g _30337_ (.A(_08574_), .B(_08579_), .Y(_01364_));
NAND_g _30338_ (.A(_10882_), .B(_08580_), .Y(_08581_));
NAND_g _30339_ (.A(resetn), .B(_08581_), .Y(_08582_));
NOR_g _30340_ (.A(_10882_), .B(_08580_), .Y(_08583_));
NOR_g _30341_ (.A(_08582_), .B(_08583_), .Y(_01365_));
NOR_g _30342_ (.A(count_instr[19]), .B(_08583_), .Y(_08584_));
AND_g _30343_ (.A(count_instr[19]), .B(count_instr[18]), .Y(_08585_));
NOR_g _30344_ (.A(_10963_), .B(_08584_), .Y(_08586_));
NAND_g _30345_ (.A(count_instr[19]), .B(_08583_), .Y(_08587_));
AND_g _30346_ (.A(count_instr[18]), .B(count_instr[17]), .Y(_08588_));
AND_g _30347_ (.A(count_instr[19]), .B(_08588_), .Y(_08589_));
AND_g _30348_ (.A(_08573_), .B(_08589_), .Y(_08590_));
AND_g _30349_ (.A(_08586_), .B(_08587_), .Y(_01366_));
NAND_g _30350_ (.A(_10881_), .B(_08587_), .Y(_08591_));
AND_g _30351_ (.A(resetn), .B(_08591_), .Y(_08592_));
NAND_g _30352_ (.A(count_instr[20]), .B(_08590_), .Y(_08593_));
AND_g _30353_ (.A(_08592_), .B(_08593_), .Y(_01367_));
NAND_g _30354_ (.A(_10880_), .B(_08593_), .Y(_08594_));
AND_g _30355_ (.A(count_instr[21]), .B(count_instr[20]), .Y(_08595_));
AND_g _30356_ (.A(_08585_), .B(_08595_), .Y(_08596_));
NAND_g _30357_ (.A(_08577_), .B(_08596_), .Y(_08597_));
NAND_g _30358_ (.A(resetn), .B(_08594_), .Y(_08598_));
NOR_g _30359_ (.A(_10880_), .B(_08593_), .Y(_08599_));
NOR_g _30360_ (.A(_08598_), .B(_08599_), .Y(_01368_));
NAND_g _30361_ (.A(_10879_), .B(_08597_), .Y(_08600_));
AND_g _30362_ (.A(resetn), .B(_08600_), .Y(_08601_));
NAND_g _30363_ (.A(count_instr[22]), .B(_08599_), .Y(_08602_));
AND_g _30364_ (.A(_08601_), .B(_08602_), .Y(_01369_));
NAND_g _30365_ (.A(_10878_), .B(_08602_), .Y(_08603_));
AND_g _30366_ (.A(count_instr[23]), .B(count_instr[22]), .Y(_08604_));
AND_g _30367_ (.A(_08596_), .B(_08604_), .Y(_08605_));
AND_g _30368_ (.A(_08577_), .B(_08605_), .Y(_08606_));
NOR_g _30369_ (.A(_10963_), .B(_08606_), .Y(_08607_));
AND_g _30370_ (.A(_08603_), .B(_08607_), .Y(_01370_));
AND_g _30371_ (.A(count_instr[16]), .B(count_instr[14]), .Y(_08608_));
AND_g _30372_ (.A(_08595_), .B(_08608_), .Y(_08609_));
AND_g _30373_ (.A(count_instr[15]), .B(_08604_), .Y(_08610_));
AND_g _30374_ (.A(_08589_), .B(_08610_), .Y(_08611_));
AND_g _30375_ (.A(_08609_), .B(_08611_), .Y(_08612_));
AND_g _30376_ (.A(_08555_), .B(_08612_), .Y(_08613_));
AND_g _30377_ (.A(count_instr[22]), .B(_08589_), .Y(_08614_));
AND_g _30378_ (.A(count_instr[23]), .B(count_instr[21]), .Y(_08615_));
AND_g _30379_ (.A(count_instr[20]), .B(_08615_), .Y(_08616_));
AND_g _30380_ (.A(_08572_), .B(_08616_), .Y(_08617_));
AND_g _30381_ (.A(_08614_), .B(_08617_), .Y(_08618_));
NAND_g _30382_ (.A(_08560_), .B(_08618_), .Y(_08619_));
NAND_g _30383_ (.A(_10877_), .B(_08619_), .Y(_08620_));
NAND_g _30384_ (.A(resetn), .B(_08620_), .Y(_08621_));
AND_g _30385_ (.A(count_instr[24]), .B(_08606_), .Y(_08622_));
NOR_g _30386_ (.A(_08621_), .B(_08622_), .Y(_01371_));
NOR_g _30387_ (.A(count_instr[25]), .B(_08622_), .Y(_08623_));
NOR_g _30388_ (.A(_10963_), .B(_08623_), .Y(_08624_));
NAND_g _30389_ (.A(count_instr[25]), .B(_08622_), .Y(_08625_));
AND_g _30390_ (.A(count_instr[25]), .B(count_instr[24]), .Y(_08626_));
AND_g _30391_ (.A(_08613_), .B(_08626_), .Y(_08627_));
AND_g _30392_ (.A(_08624_), .B(_08625_), .Y(_01372_));
NAND_g _30393_ (.A(_10876_), .B(_08625_), .Y(_08628_));
AND_g _30394_ (.A(resetn), .B(_08628_), .Y(_08629_));
AND_g _30395_ (.A(count_instr[26]), .B(_08627_), .Y(_08630_));
NAND_g _30396_ (.A(count_instr[26]), .B(_08627_), .Y(_08631_));
AND_g _30397_ (.A(_08629_), .B(_08631_), .Y(_01373_));
NAND_g _30398_ (.A(_10875_), .B(_08631_), .Y(_08632_));
AND_g _30399_ (.A(count_instr[27]), .B(count_instr[26]), .Y(_08633_));
NAND_g _30400_ (.A(resetn), .B(_08632_), .Y(_08634_));
AND_g _30401_ (.A(count_instr[27]), .B(_08630_), .Y(_08635_));
NOR_g _30402_ (.A(_08634_), .B(_08635_), .Y(_01374_));
NOR_g _30403_ (.A(count_instr[28]), .B(_08635_), .Y(_08636_));
NOR_g _30404_ (.A(_10963_), .B(_08636_), .Y(_08637_));
NAND_g _30405_ (.A(count_instr[28]), .B(_08635_), .Y(_08638_));
NOT_g _30406_ (.A(_08638_), .Y(_08639_));
AND_g _30407_ (.A(_08637_), .B(_08638_), .Y(_01375_));
NAND_g _30408_ (.A(_10874_), .B(_08638_), .Y(_08640_));
AND_g _30409_ (.A(count_instr[29]), .B(count_instr[28]), .Y(_08641_));
AND_g _30410_ (.A(_08633_), .B(_08641_), .Y(_08642_));
AND_g _30411_ (.A(resetn), .B(_08640_), .Y(_08643_));
NAND_g _30412_ (.A(count_instr[29]), .B(_08639_), .Y(_08644_));
NOT_g _30413_ (.A(_08644_), .Y(_08645_));
AND_g _30414_ (.A(_08643_), .B(_08644_), .Y(_01376_));
NAND_g _30415_ (.A(_10873_), .B(_08644_), .Y(_08646_));
AND_g _30416_ (.A(resetn), .B(_08646_), .Y(_08647_));
NAND_g _30417_ (.A(count_instr[30]), .B(_08645_), .Y(_08648_));
AND_g _30418_ (.A(_08647_), .B(_08648_), .Y(_01377_));
NAND_g _30419_ (.A(_10872_), .B(_08648_), .Y(_08649_));
AND_g _30420_ (.A(count_instr[31]), .B(count_instr[30]), .Y(_08650_));
AND_g _30421_ (.A(count_instr[25]), .B(_08650_), .Y(_08651_));
AND_g _30422_ (.A(_08642_), .B(_08651_), .Y(_08652_));
AND_g _30423_ (.A(_08622_), .B(_08652_), .Y(_08653_));
NAND_g _30424_ (.A(resetn), .B(_08649_), .Y(_08654_));
AND_g _30425_ (.A(count_instr[31]), .B(_08641_), .Y(_08655_));
AND_g _30426_ (.A(count_instr[30]), .B(_08655_), .Y(_08656_));
AND_g _30427_ (.A(_08633_), .B(_08656_), .Y(_08657_));
AND_g _30428_ (.A(_08626_), .B(_08657_), .Y(_08658_));
AND_g _30429_ (.A(_08613_), .B(_08658_), .Y(_08659_));
AND_g _30430_ (.A(_08618_), .B(_08658_), .Y(_08660_));
AND_g _30431_ (.A(_08560_), .B(_08660_), .Y(_08661_));
NOR_g _30432_ (.A(_08654_), .B(_08659_), .Y(_01378_));
NOR_g _30433_ (.A(count_instr[32]), .B(_08661_), .Y(_08662_));
NOR_g _30434_ (.A(_10963_), .B(_08662_), .Y(_08663_));
AND_g _30435_ (.A(count_instr[32]), .B(_08659_), .Y(_08664_));
NAND_g _30436_ (.A(count_instr[32]), .B(_08661_), .Y(_08665_));
NOT_g _30437_ (.A(_08665_), .Y(_08666_));
AND_g _30438_ (.A(_08663_), .B(_08665_), .Y(_01379_));
NAND_g _30439_ (.A(_10871_), .B(_08665_), .Y(_08667_));
AND_g _30440_ (.A(count_instr[33]), .B(count_instr[32]), .Y(_08668_));
AND_g _30441_ (.A(resetn), .B(_08667_), .Y(_08669_));
NAND_g _30442_ (.A(count_instr[33]), .B(_08664_), .Y(_08670_));
NOT_g _30443_ (.A(_08670_), .Y(_08671_));
NAND_g _30444_ (.A(count_instr[33]), .B(_08666_), .Y(_08672_));
AND_g _30445_ (.A(_08669_), .B(_08672_), .Y(_01380_));
NAND_g _30446_ (.A(_10870_), .B(_08672_), .Y(_08673_));
AND_g _30447_ (.A(resetn), .B(_08673_), .Y(_08674_));
NAND_g _30448_ (.A(count_instr[34]), .B(_08671_), .Y(_08675_));
AND_g _30449_ (.A(count_instr[34]), .B(count_instr[33]), .Y(_08676_));
AND_g _30450_ (.A(_08674_), .B(_08675_), .Y(_01381_));
NAND_g _30451_ (.A(_10869_), .B(_08675_), .Y(_08677_));
AND_g _30452_ (.A(count_instr[35]), .B(count_instr[34]), .Y(_08678_));
AND_g _30453_ (.A(_08668_), .B(_08678_), .Y(_08679_));
AND_g _30454_ (.A(_08653_), .B(_08679_), .Y(_08680_));
NAND_g _30455_ (.A(resetn), .B(_08677_), .Y(_08681_));
AND_g _30456_ (.A(count_instr[35]), .B(_08676_), .Y(_08682_));
AND_g _30457_ (.A(_08666_), .B(_08682_), .Y(_08683_));
NOR_g _30458_ (.A(_08681_), .B(_08683_), .Y(_01382_));
NOR_g _30459_ (.A(count_instr[36]), .B(_08683_), .Y(_08684_));
NOR_g _30460_ (.A(_10963_), .B(_08684_), .Y(_08685_));
AND_g _30461_ (.A(count_instr[36]), .B(_08680_), .Y(_08686_));
NAND_g _30462_ (.A(count_instr[36]), .B(_08683_), .Y(_08687_));
NOT_g _30463_ (.A(_08687_), .Y(_08688_));
AND_g _30464_ (.A(_08685_), .B(_08687_), .Y(_01383_));
NAND_g _30465_ (.A(_10868_), .B(_08687_), .Y(_08689_));
AND_g _30466_ (.A(resetn), .B(_08689_), .Y(_08690_));
AND_g _30467_ (.A(count_instr[37]), .B(_08686_), .Y(_08691_));
NAND_g _30468_ (.A(count_instr[37]), .B(_08688_), .Y(_08692_));
AND_g _30469_ (.A(_08690_), .B(_08692_), .Y(_01384_));
NAND_g _30470_ (.A(_10867_), .B(_08692_), .Y(_08693_));
AND_g _30471_ (.A(resetn), .B(_08693_), .Y(_08694_));
NAND_g _30472_ (.A(count_instr[38]), .B(_08691_), .Y(_08695_));
AND_g _30473_ (.A(_08694_), .B(_08695_), .Y(_01385_));
XNOR_g _30474_ (.A(count_instr[39]), .B(_08695_), .Y(_08696_));
AND_g _30475_ (.A(resetn), .B(_08696_), .Y(_01386_));
AND_g _30476_ (.A(count_instr[39]), .B(count_instr[38]), .Y(_08697_));
AND_g _30477_ (.A(count_instr[37]), .B(_08697_), .Y(_08698_));
AND_g _30478_ (.A(_08686_), .B(_08698_), .Y(_08699_));
AND_g _30479_ (.A(count_instr[38]), .B(_08660_), .Y(_08700_));
AND_g _30480_ (.A(count_instr[39]), .B(count_instr[32]), .Y(_08701_));
AND_g _30481_ (.A(_08682_), .B(_08701_), .Y(_08702_));
AND_g _30482_ (.A(count_instr[37]), .B(_08702_), .Y(_08703_));
AND_g _30483_ (.A(count_instr[36]), .B(_08703_), .Y(_08704_));
AND_g _30484_ (.A(_08559_), .B(_08704_), .Y(_08705_));
AND_g _30485_ (.A(_08700_), .B(_08705_), .Y(_08706_));
AND_g _30486_ (.A(launch_next_insn), .B(_08706_), .Y(_08707_));
NOR_g _30487_ (.A(count_instr[40]), .B(_08707_), .Y(_08708_));
NOR_g _30488_ (.A(_10963_), .B(_08708_), .Y(_08709_));
NAND_g _30489_ (.A(count_instr[40]), .B(_08699_), .Y(_08710_));
AND_g _30490_ (.A(_08709_), .B(_08710_), .Y(_01387_));
NAND_g _30491_ (.A(_10866_), .B(_08710_), .Y(_08711_));
AND_g _30492_ (.A(count_instr[41]), .B(count_instr[40]), .Y(_08712_));
AND_g _30493_ (.A(_08699_), .B(_08712_), .Y(_08713_));
NOR_g _30494_ (.A(_10963_), .B(_08713_), .Y(_08714_));
AND_g _30495_ (.A(_08707_), .B(_08712_), .Y(_08715_));
AND_g _30496_ (.A(_08711_), .B(_08714_), .Y(_01388_));
NOR_g _30497_ (.A(count_instr[42]), .B(_08715_), .Y(_08716_));
NOR_g _30498_ (.A(_10963_), .B(_08716_), .Y(_08717_));
NAND_g _30499_ (.A(count_instr[42]), .B(_08713_), .Y(_08718_));
NOT_g _30500_ (.A(_08718_), .Y(_08719_));
AND_g _30501_ (.A(count_instr[42]), .B(_08715_), .Y(_08720_));
AND_g _30502_ (.A(_08717_), .B(_08718_), .Y(_01389_));
NAND_g _30503_ (.A(_10865_), .B(_08718_), .Y(_08721_));
AND_g _30504_ (.A(resetn), .B(_08721_), .Y(_08722_));
NAND_g _30505_ (.A(count_instr[43]), .B(_08719_), .Y(_08723_));
AND_g _30506_ (.A(count_instr[43]), .B(_08720_), .Y(_08724_));
AND_g _30507_ (.A(_08722_), .B(_08723_), .Y(_01390_));
NAND_g _30508_ (.A(_10864_), .B(_08723_), .Y(_08725_));
AND_g _30509_ (.A(resetn), .B(_08725_), .Y(_08726_));
AND_g _30510_ (.A(count_instr[44]), .B(_08724_), .Y(_08727_));
NAND_g _30511_ (.A(count_instr[44]), .B(_08724_), .Y(_08728_));
AND_g _30512_ (.A(_08726_), .B(_08728_), .Y(_01391_));
NAND_g _30513_ (.A(_10863_), .B(_08728_), .Y(_08729_));
AND_g _30514_ (.A(resetn), .B(_08729_), .Y(_08730_));
NAND_g _30515_ (.A(count_instr[45]), .B(_08727_), .Y(_08731_));
AND_g _30516_ (.A(_08730_), .B(_08731_), .Y(_01392_));
NAND_g _30517_ (.A(_10862_), .B(_08731_), .Y(_08732_));
NAND_g _30518_ (.A(resetn), .B(_08732_), .Y(_08733_));
NOR_g _30519_ (.A(_10862_), .B(_08731_), .Y(_08734_));
NOR_g _30520_ (.A(_08733_), .B(_08734_), .Y(_01393_));
AND_g _30521_ (.A(count_instr[47]), .B(_08734_), .Y(_08735_));
NOR_g _30522_ (.A(count_instr[47]), .B(_08734_), .Y(_08736_));
NOT_g _30523_ (.A(_08736_), .Y(_08737_));
NAND_g _30524_ (.A(resetn), .B(_08737_), .Y(_08738_));
NOR_g _30525_ (.A(_08735_), .B(_08738_), .Y(_01394_));
AND_g _30526_ (.A(count_instr[48]), .B(_08735_), .Y(_08739_));
NAND_g _30527_ (.A(count_instr[48]), .B(_08735_), .Y(_08740_));
NOR_g _30528_ (.A(count_instr[48]), .B(_08735_), .Y(_08741_));
NOR_g _30529_ (.A(_10963_), .B(_08741_), .Y(_08742_));
AND_g _30530_ (.A(_08740_), .B(_08742_), .Y(_01395_));
NOR_g _30531_ (.A(count_instr[49]), .B(_08739_), .Y(_08743_));
NOR_g _30532_ (.A(_10963_), .B(_08743_), .Y(_08744_));
NAND_g _30533_ (.A(count_instr[49]), .B(_08739_), .Y(_08745_));
NOT_g _30534_ (.A(_08745_), .Y(_08746_));
AND_g _30535_ (.A(count_instr[49]), .B(count_instr[48]), .Y(_08747_));
AND_g _30536_ (.A(_08744_), .B(_08745_), .Y(_01396_));
NAND_g _30537_ (.A(_10861_), .B(_08745_), .Y(_08748_));
AND_g _30538_ (.A(resetn), .B(_08748_), .Y(_08749_));
NAND_g _30539_ (.A(count_instr[50]), .B(_08746_), .Y(_08750_));
AND_g _30540_ (.A(_08749_), .B(_08750_), .Y(_01397_));
NAND_g _30541_ (.A(_10860_), .B(_08750_), .Y(_08751_));
NAND_g _30542_ (.A(count_instr[51]), .B(count_instr[50]), .Y(_08752_));
NOR_g _30543_ (.A(_08745_), .B(_08752_), .Y(_08753_));
NOR_g _30544_ (.A(_10963_), .B(_08753_), .Y(_08754_));
AND_g _30545_ (.A(_08751_), .B(_08754_), .Y(_01398_));
AND_g _30546_ (.A(count_instr[51]), .B(_08747_), .Y(_08755_));
AND_g _30547_ (.A(count_instr[50]), .B(_08755_), .Y(_08756_));
AND_g _30548_ (.A(_08735_), .B(_08756_), .Y(_08757_));
NOR_g _30549_ (.A(count_instr[52]), .B(_08757_), .Y(_08758_));
NOR_g _30550_ (.A(_10963_), .B(_08758_), .Y(_08759_));
NAND_g _30551_ (.A(count_instr[52]), .B(_08757_), .Y(_08760_));
AND_g _30552_ (.A(_08759_), .B(_08760_), .Y(_01399_));
NAND_g _30553_ (.A(_10859_), .B(_08760_), .Y(_08761_));
AND_g _30554_ (.A(count_instr[53]), .B(count_instr[52]), .Y(_08762_));
AND_g _30555_ (.A(_08756_), .B(_08762_), .Y(_08763_));
NAND_g _30556_ (.A(_08735_), .B(_08763_), .Y(_08764_));
AND_g _30557_ (.A(resetn), .B(_08764_), .Y(_08765_));
AND_g _30558_ (.A(_08761_), .B(_08765_), .Y(_01400_));
NOR_g _30559_ (.A(_10858_), .B(_08764_), .Y(_08766_));
NAND_g _30560_ (.A(_10858_), .B(_08764_), .Y(_08767_));
NAND_g _30561_ (.A(resetn), .B(_08767_), .Y(_08768_));
NOR_g _30562_ (.A(_08766_), .B(_08768_), .Y(_01401_));
NAND_g _30563_ (.A(count_instr[55]), .B(_08766_), .Y(_08769_));
NOR_g _30564_ (.A(count_instr[55]), .B(_08766_), .Y(_08770_));
NOR_g _30565_ (.A(_10963_), .B(_08770_), .Y(_08771_));
AND_g _30566_ (.A(_08769_), .B(_08771_), .Y(_01402_));
NAND_g _30567_ (.A(_10857_), .B(_08769_), .Y(_08772_));
NAND_g _30568_ (.A(resetn), .B(_08772_), .Y(_08773_));
NOR_g _30569_ (.A(_10857_), .B(_08769_), .Y(_08774_));
NOR_g _30570_ (.A(_08773_), .B(_08774_), .Y(_01403_));
NOR_g _30571_ (.A(count_instr[57]), .B(_08774_), .Y(_08775_));
NOR_g _30572_ (.A(_10963_), .B(_08775_), .Y(_08776_));
NAND_g _30573_ (.A(count_instr[57]), .B(_08774_), .Y(_08777_));
AND_g _30574_ (.A(_08776_), .B(_08777_), .Y(_01404_));
NAND_g _30575_ (.A(_10856_), .B(_08777_), .Y(_08778_));
NAND_g _30576_ (.A(resetn), .B(_08778_), .Y(_08779_));
NOR_g _30577_ (.A(_10856_), .B(_08777_), .Y(_08780_));
NOR_g _30578_ (.A(_08779_), .B(_08780_), .Y(_01405_));
NOR_g _30579_ (.A(count_instr[59]), .B(_08780_), .Y(_08781_));
NOR_g _30580_ (.A(_10963_), .B(_08781_), .Y(_08782_));
NAND_g _30581_ (.A(count_instr[59]), .B(_08780_), .Y(_08783_));
AND_g _30582_ (.A(_08782_), .B(_08783_), .Y(_01406_));
NAND_g _30583_ (.A(_10855_), .B(_08783_), .Y(_08784_));
NAND_g _30584_ (.A(resetn), .B(_08784_), .Y(_08785_));
NOR_g _30585_ (.A(_10855_), .B(_08783_), .Y(_08786_));
NOR_g _30586_ (.A(_08785_), .B(_08786_), .Y(_01407_));
NOR_g _30587_ (.A(count_instr[61]), .B(_08786_), .Y(_08787_));
NOR_g _30588_ (.A(_10963_), .B(_08787_), .Y(_08788_));
NAND_g _30589_ (.A(count_instr[61]), .B(_08786_), .Y(_08789_));
NOT_g _30590_ (.A(_08789_), .Y(_08790_));
AND_g _30591_ (.A(_08788_), .B(_08789_), .Y(_01408_));
NAND_g _30592_ (.A(_10854_), .B(_08789_), .Y(_08791_));
AND_g _30593_ (.A(resetn), .B(_08791_), .Y(_08792_));
NAND_g _30594_ (.A(count_instr[62]), .B(_08790_), .Y(_08793_));
AND_g _30595_ (.A(_08792_), .B(_08793_), .Y(_01409_));
XNOR_g _30596_ (.A(count_instr[63]), .B(_08793_), .Y(_08794_));
AND_g _30597_ (.A(resetn), .B(_08794_), .Y(_01410_));
AND_g _30598_ (.A(_11287_), .B(_11765_), .Y(_08795_));
NAND_g _30599_ (.A(_11287_), .B(_11765_), .Y(_08796_));
NAND_g _30600_ (.A(_11301_), .B(_08795_), .Y(_08797_));
NAND_g _30601_ (.A(cpuregs_30[0]), .B(_08796_), .Y(_08798_));
NAND_g _30602_ (.A(_08797_), .B(_08798_), .Y(_01411_));
NAND_g _30603_ (.A(_11310_), .B(_08795_), .Y(_08799_));
NAND_g _30604_ (.A(cpuregs_30[1]), .B(_08796_), .Y(_08800_));
NAND_g _30605_ (.A(_08799_), .B(_08800_), .Y(_01412_));
NAND_g _30606_ (.A(_11319_), .B(_08795_), .Y(_08801_));
NAND_g _30607_ (.A(cpuregs_30[2]), .B(_08796_), .Y(_08802_));
NAND_g _30608_ (.A(_08801_), .B(_08802_), .Y(_01413_));
NAND_g _30609_ (.A(_11332_), .B(_08795_), .Y(_08803_));
NAND_g _30610_ (.A(cpuregs_30[3]), .B(_08796_), .Y(_08804_));
NAND_g _30611_ (.A(_08803_), .B(_08804_), .Y(_01414_));
NAND_g _30612_ (.A(_11345_), .B(_08795_), .Y(_08805_));
NAND_g _30613_ (.A(cpuregs_30[4]), .B(_08796_), .Y(_08806_));
NAND_g _30614_ (.A(_08805_), .B(_08806_), .Y(_01415_));
NAND_g _30615_ (.A(_11358_), .B(_08795_), .Y(_08807_));
NAND_g _30616_ (.A(cpuregs_30[5]), .B(_08796_), .Y(_08808_));
NAND_g _30617_ (.A(_08807_), .B(_08808_), .Y(_01416_));
NAND_g _30618_ (.A(_11371_), .B(_08795_), .Y(_08809_));
NAND_g _30619_ (.A(cpuregs_30[6]), .B(_08796_), .Y(_08810_));
NAND_g _30620_ (.A(_08809_), .B(_08810_), .Y(_01417_));
NAND_g _30621_ (.A(_11384_), .B(_08795_), .Y(_08811_));
NAND_g _30622_ (.A(cpuregs_30[7]), .B(_08796_), .Y(_08812_));
NAND_g _30623_ (.A(_08811_), .B(_08812_), .Y(_01418_));
NAND_g _30624_ (.A(_11397_), .B(_08795_), .Y(_08813_));
NAND_g _30625_ (.A(cpuregs_30[8]), .B(_08796_), .Y(_08814_));
NAND_g _30626_ (.A(_08813_), .B(_08814_), .Y(_01419_));
NAND_g _30627_ (.A(_11410_), .B(_08795_), .Y(_08815_));
NAND_g _30628_ (.A(cpuregs_30[9]), .B(_08796_), .Y(_08816_));
NAND_g _30629_ (.A(_08815_), .B(_08816_), .Y(_01420_));
NAND_g _30630_ (.A(_11423_), .B(_08795_), .Y(_08817_));
NAND_g _30631_ (.A(cpuregs_30[10]), .B(_08796_), .Y(_08818_));
NAND_g _30632_ (.A(_08817_), .B(_08818_), .Y(_01421_));
NAND_g _30633_ (.A(_11436_), .B(_08795_), .Y(_08819_));
NAND_g _30634_ (.A(cpuregs_30[11]), .B(_08796_), .Y(_08820_));
NAND_g _30635_ (.A(_08819_), .B(_08820_), .Y(_01422_));
NAND_g _30636_ (.A(_11449_), .B(_08795_), .Y(_08821_));
NAND_g _30637_ (.A(cpuregs_30[12]), .B(_08796_), .Y(_08822_));
NAND_g _30638_ (.A(_08821_), .B(_08822_), .Y(_01423_));
NAND_g _30639_ (.A(_11462_), .B(_08795_), .Y(_08823_));
NAND_g _30640_ (.A(cpuregs_30[13]), .B(_08796_), .Y(_08824_));
NAND_g _30641_ (.A(_08823_), .B(_08824_), .Y(_01424_));
NAND_g _30642_ (.A(_11475_), .B(_08795_), .Y(_08825_));
NAND_g _30643_ (.A(cpuregs_30[14]), .B(_08796_), .Y(_08826_));
NAND_g _30644_ (.A(_08825_), .B(_08826_), .Y(_01425_));
NAND_g _30645_ (.A(_11488_), .B(_08795_), .Y(_08827_));
NAND_g _30646_ (.A(cpuregs_30[15]), .B(_08796_), .Y(_08828_));
NAND_g _30647_ (.A(_08827_), .B(_08828_), .Y(_01426_));
NAND_g _30648_ (.A(_11501_), .B(_08795_), .Y(_08829_));
NAND_g _30649_ (.A(cpuregs_30[16]), .B(_08796_), .Y(_08830_));
NAND_g _30650_ (.A(_08829_), .B(_08830_), .Y(_01427_));
NAND_g _30651_ (.A(_11514_), .B(_08795_), .Y(_08831_));
NAND_g _30652_ (.A(cpuregs_30[17]), .B(_08796_), .Y(_08832_));
NAND_g _30653_ (.A(_08831_), .B(_08832_), .Y(_01428_));
NAND_g _30654_ (.A(_11527_), .B(_08795_), .Y(_08833_));
NAND_g _30655_ (.A(cpuregs_30[18]), .B(_08796_), .Y(_08834_));
NAND_g _30656_ (.A(_08833_), .B(_08834_), .Y(_01429_));
NAND_g _30657_ (.A(_11540_), .B(_08795_), .Y(_08835_));
NAND_g _30658_ (.A(cpuregs_30[19]), .B(_08796_), .Y(_08836_));
NAND_g _30659_ (.A(_08835_), .B(_08836_), .Y(_01430_));
NAND_g _30660_ (.A(_11553_), .B(_08795_), .Y(_08837_));
NAND_g _30661_ (.A(cpuregs_30[20]), .B(_08796_), .Y(_08838_));
NAND_g _30662_ (.A(_08837_), .B(_08838_), .Y(_01431_));
NAND_g _30663_ (.A(_11566_), .B(_08795_), .Y(_08839_));
NAND_g _30664_ (.A(cpuregs_30[21]), .B(_08796_), .Y(_08840_));
NAND_g _30665_ (.A(_08839_), .B(_08840_), .Y(_01432_));
NAND_g _30666_ (.A(_11579_), .B(_08795_), .Y(_08841_));
NAND_g _30667_ (.A(cpuregs_30[22]), .B(_08796_), .Y(_08842_));
NAND_g _30668_ (.A(_08841_), .B(_08842_), .Y(_01433_));
NAND_g _30669_ (.A(_11592_), .B(_08795_), .Y(_08843_));
NAND_g _30670_ (.A(cpuregs_30[23]), .B(_08796_), .Y(_08844_));
NAND_g _30671_ (.A(_08843_), .B(_08844_), .Y(_01434_));
NAND_g _30672_ (.A(_11605_), .B(_08795_), .Y(_08845_));
NAND_g _30673_ (.A(cpuregs_30[24]), .B(_08796_), .Y(_08846_));
NAND_g _30674_ (.A(_08845_), .B(_08846_), .Y(_01435_));
NAND_g _30675_ (.A(_11618_), .B(_08795_), .Y(_08847_));
NAND_g _30676_ (.A(cpuregs_30[25]), .B(_08796_), .Y(_08848_));
NAND_g _30677_ (.A(_08847_), .B(_08848_), .Y(_01436_));
NAND_g _30678_ (.A(_11631_), .B(_08795_), .Y(_08849_));
NAND_g _30679_ (.A(cpuregs_30[26]), .B(_08796_), .Y(_08850_));
NAND_g _30680_ (.A(_08849_), .B(_08850_), .Y(_01437_));
NAND_g _30681_ (.A(_11644_), .B(_08795_), .Y(_08851_));
NAND_g _30682_ (.A(cpuregs_30[27]), .B(_08796_), .Y(_08852_));
NAND_g _30683_ (.A(_08851_), .B(_08852_), .Y(_01438_));
NAND_g _30684_ (.A(_11657_), .B(_08795_), .Y(_08853_));
NAND_g _30685_ (.A(cpuregs_30[28]), .B(_08796_), .Y(_08854_));
NAND_g _30686_ (.A(_08853_), .B(_08854_), .Y(_01439_));
NAND_g _30687_ (.A(_11670_), .B(_08795_), .Y(_08855_));
NAND_g _30688_ (.A(cpuregs_30[29]), .B(_08796_), .Y(_08856_));
NAND_g _30689_ (.A(_08855_), .B(_08856_), .Y(_01440_));
NAND_g _30690_ (.A(_11683_), .B(_08795_), .Y(_08857_));
NAND_g _30691_ (.A(cpuregs_30[30]), .B(_08796_), .Y(_08858_));
NAND_g _30692_ (.A(_08857_), .B(_08858_), .Y(_01441_));
NAND_g _30693_ (.A(_11695_), .B(_08795_), .Y(_08859_));
NAND_g _30694_ (.A(cpuregs_30[31]), .B(_08796_), .Y(_08860_));
NAND_g _30695_ (.A(_08859_), .B(_08860_), .Y(_01442_));
AND_g _30696_ (.A(_12002_), .B(_04359_), .Y(_08861_));
NAND_g _30697_ (.A(_12002_), .B(_04359_), .Y(_08862_));
NAND_g _30698_ (.A(cpuregs_24[0]), .B(_08862_), .Y(_08863_));
NAND_g _30699_ (.A(_11301_), .B(_08861_), .Y(_08864_));
AND_g _30700_ (.A(_12000_), .B(_12075_), .Y(_08865_));
NAND_g _30701_ (.A(_12000_), .B(_12075_), .Y(_08866_));
NAND_g _30702_ (.A(_08863_), .B(_08864_), .Y(_01443_));
NAND_g _30703_ (.A(cpuregs_24[1]), .B(_08862_), .Y(_08867_));
NAND_g _30704_ (.A(_11310_), .B(_08861_), .Y(_08868_));
NAND_g _30705_ (.A(_08867_), .B(_08868_), .Y(_01444_));
NAND_g _30706_ (.A(cpuregs_24[2]), .B(_08862_), .Y(_08869_));
NAND_g _30707_ (.A(_11319_), .B(_08861_), .Y(_08870_));
NAND_g _30708_ (.A(_08869_), .B(_08870_), .Y(_01445_));
NAND_g _30709_ (.A(cpuregs_24[3]), .B(_08862_), .Y(_08871_));
NAND_g _30710_ (.A(_11332_), .B(_08861_), .Y(_08872_));
NAND_g _30711_ (.A(_08871_), .B(_08872_), .Y(_01446_));
NAND_g _30712_ (.A(cpuregs_24[4]), .B(_08862_), .Y(_08873_));
NAND_g _30713_ (.A(_11345_), .B(_08861_), .Y(_08874_));
NAND_g _30714_ (.A(_08873_), .B(_08874_), .Y(_01447_));
NAND_g _30715_ (.A(cpuregs_24[5]), .B(_08862_), .Y(_08875_));
NAND_g _30716_ (.A(_11358_), .B(_08861_), .Y(_08876_));
NAND_g _30717_ (.A(_08875_), .B(_08876_), .Y(_01448_));
NAND_g _30718_ (.A(cpuregs_24[6]), .B(_08862_), .Y(_08877_));
NAND_g _30719_ (.A(_11371_), .B(_08861_), .Y(_08878_));
NAND_g _30720_ (.A(_08877_), .B(_08878_), .Y(_01449_));
NAND_g _30721_ (.A(cpuregs_24[7]), .B(_08862_), .Y(_08879_));
NAND_g _30722_ (.A(_11384_), .B(_08861_), .Y(_08880_));
NAND_g _30723_ (.A(_08879_), .B(_08880_), .Y(_01450_));
NAND_g _30724_ (.A(cpuregs_24[8]), .B(_08862_), .Y(_08881_));
NAND_g _30725_ (.A(_11397_), .B(_08861_), .Y(_08882_));
NAND_g _30726_ (.A(_08881_), .B(_08882_), .Y(_01451_));
NAND_g _30727_ (.A(cpuregs_24[9]), .B(_08862_), .Y(_08883_));
NAND_g _30728_ (.A(_11410_), .B(_08861_), .Y(_08884_));
NAND_g _30729_ (.A(_08883_), .B(_08884_), .Y(_01452_));
NAND_g _30730_ (.A(cpuregs_24[10]), .B(_08862_), .Y(_08885_));
NAND_g _30731_ (.A(_11423_), .B(_08861_), .Y(_08886_));
NAND_g _30732_ (.A(_08885_), .B(_08886_), .Y(_01453_));
NAND_g _30733_ (.A(cpuregs_24[11]), .B(_08862_), .Y(_08887_));
NAND_g _30734_ (.A(_11436_), .B(_08861_), .Y(_08888_));
NAND_g _30735_ (.A(_08887_), .B(_08888_), .Y(_01454_));
NAND_g _30736_ (.A(cpuregs_24[12]), .B(_08862_), .Y(_08889_));
NAND_g _30737_ (.A(_11449_), .B(_08861_), .Y(_08890_));
NAND_g _30738_ (.A(_08889_), .B(_08890_), .Y(_01455_));
NAND_g _30739_ (.A(cpuregs_24[13]), .B(_08862_), .Y(_08891_));
NAND_g _30740_ (.A(_11462_), .B(_08861_), .Y(_08892_));
NAND_g _30741_ (.A(_08891_), .B(_08892_), .Y(_01456_));
NAND_g _30742_ (.A(cpuregs_24[14]), .B(_08862_), .Y(_08893_));
NAND_g _30743_ (.A(_11475_), .B(_08861_), .Y(_08894_));
NAND_g _30744_ (.A(_08893_), .B(_08894_), .Y(_01457_));
NAND_g _30745_ (.A(cpuregs_24[15]), .B(_08862_), .Y(_08895_));
NAND_g _30746_ (.A(_11488_), .B(_08861_), .Y(_08896_));
NAND_g _30747_ (.A(_08895_), .B(_08896_), .Y(_01458_));
NAND_g _30748_ (.A(cpuregs_24[16]), .B(_08862_), .Y(_08897_));
NAND_g _30749_ (.A(_11501_), .B(_08861_), .Y(_08898_));
NAND_g _30750_ (.A(_08897_), .B(_08898_), .Y(_01459_));
NAND_g _30751_ (.A(cpuregs_24[17]), .B(_08866_), .Y(_08899_));
NAND_g _30752_ (.A(_11514_), .B(_08865_), .Y(_08900_));
NAND_g _30753_ (.A(_08899_), .B(_08900_), .Y(_01460_));
NAND_g _30754_ (.A(cpuregs_24[18]), .B(_08866_), .Y(_08901_));
NAND_g _30755_ (.A(_11527_), .B(_08865_), .Y(_08902_));
NAND_g _30756_ (.A(_08901_), .B(_08902_), .Y(_01461_));
NAND_g _30757_ (.A(cpuregs_24[19]), .B(_08866_), .Y(_08903_));
NAND_g _30758_ (.A(_11540_), .B(_08865_), .Y(_08904_));
NAND_g _30759_ (.A(_08903_), .B(_08904_), .Y(_01462_));
NAND_g _30760_ (.A(cpuregs_24[20]), .B(_08866_), .Y(_08905_));
NAND_g _30761_ (.A(_11553_), .B(_08865_), .Y(_08906_));
NAND_g _30762_ (.A(_08905_), .B(_08906_), .Y(_01463_));
NAND_g _30763_ (.A(cpuregs_24[21]), .B(_08866_), .Y(_08907_));
NAND_g _30764_ (.A(_11566_), .B(_08865_), .Y(_08908_));
NAND_g _30765_ (.A(_08907_), .B(_08908_), .Y(_01464_));
NAND_g _30766_ (.A(cpuregs_24[22]), .B(_08866_), .Y(_08909_));
NAND_g _30767_ (.A(_11579_), .B(_08865_), .Y(_08910_));
NAND_g _30768_ (.A(_08909_), .B(_08910_), .Y(_01465_));
NAND_g _30769_ (.A(cpuregs_24[23]), .B(_08866_), .Y(_08911_));
NAND_g _30770_ (.A(_11592_), .B(_08865_), .Y(_08912_));
NAND_g _30771_ (.A(_08911_), .B(_08912_), .Y(_01466_));
NAND_g _30772_ (.A(cpuregs_24[24]), .B(_08866_), .Y(_08913_));
NAND_g _30773_ (.A(_11605_), .B(_08865_), .Y(_08914_));
NAND_g _30774_ (.A(_08913_), .B(_08914_), .Y(_01467_));
NAND_g _30775_ (.A(cpuregs_24[25]), .B(_08866_), .Y(_08915_));
NAND_g _30776_ (.A(_11618_), .B(_08865_), .Y(_08916_));
NAND_g _30777_ (.A(_08915_), .B(_08916_), .Y(_01468_));
NAND_g _30778_ (.A(cpuregs_24[26]), .B(_08866_), .Y(_08917_));
NAND_g _30779_ (.A(_11631_), .B(_08865_), .Y(_08918_));
NAND_g _30780_ (.A(_08917_), .B(_08918_), .Y(_01469_));
NAND_g _30781_ (.A(cpuregs_24[27]), .B(_08866_), .Y(_08919_));
NAND_g _30782_ (.A(_11644_), .B(_08865_), .Y(_08920_));
NAND_g _30783_ (.A(_08919_), .B(_08920_), .Y(_01470_));
NAND_g _30784_ (.A(cpuregs_24[28]), .B(_08866_), .Y(_08921_));
NAND_g _30785_ (.A(_11657_), .B(_08865_), .Y(_08922_));
NAND_g _30786_ (.A(_08921_), .B(_08922_), .Y(_01471_));
NAND_g _30787_ (.A(cpuregs_24[29]), .B(_08866_), .Y(_08923_));
NAND_g _30788_ (.A(_11670_), .B(_08865_), .Y(_08924_));
NAND_g _30789_ (.A(_08923_), .B(_08924_), .Y(_01472_));
NAND_g _30790_ (.A(cpuregs_24[30]), .B(_08866_), .Y(_08925_));
NAND_g _30791_ (.A(_11683_), .B(_08865_), .Y(_08926_));
NAND_g _30792_ (.A(_08925_), .B(_08926_), .Y(_01473_));
NAND_g _30793_ (.A(cpuregs_24[31]), .B(_08866_), .Y(_08927_));
NAND_g _30794_ (.A(_11695_), .B(_08865_), .Y(_08928_));
NAND_g _30795_ (.A(_08927_), .B(_08928_), .Y(_01474_));
AND_g _30796_ (.A(_11765_), .B(_04292_), .Y(_08929_));
NAND_g _30797_ (.A(_11765_), .B(_04292_), .Y(_08930_));
NAND_g _30798_ (.A(_11301_), .B(_08929_), .Y(_08931_));
NAND_g _30799_ (.A(cpuregs_2[0]), .B(_08930_), .Y(_08932_));
NAND_g _30800_ (.A(_08931_), .B(_08932_), .Y(_01475_));
NAND_g _30801_ (.A(_11310_), .B(_08929_), .Y(_08933_));
NAND_g _30802_ (.A(cpuregs_2[1]), .B(_08930_), .Y(_08934_));
NAND_g _30803_ (.A(_08933_), .B(_08934_), .Y(_01476_));
NAND_g _30804_ (.A(_11319_), .B(_08929_), .Y(_08935_));
NAND_g _30805_ (.A(cpuregs_2[2]), .B(_08930_), .Y(_08936_));
NAND_g _30806_ (.A(_08935_), .B(_08936_), .Y(_01477_));
NAND_g _30807_ (.A(_11332_), .B(_08929_), .Y(_08937_));
NAND_g _30808_ (.A(cpuregs_2[3]), .B(_08930_), .Y(_08938_));
NAND_g _30809_ (.A(_08937_), .B(_08938_), .Y(_01478_));
NAND_g _30810_ (.A(_11345_), .B(_08929_), .Y(_08939_));
NAND_g _30811_ (.A(cpuregs_2[4]), .B(_08930_), .Y(_08940_));
NAND_g _30812_ (.A(_08939_), .B(_08940_), .Y(_01479_));
NAND_g _30813_ (.A(_11358_), .B(_08929_), .Y(_08941_));
NAND_g _30814_ (.A(cpuregs_2[5]), .B(_08930_), .Y(_08942_));
NAND_g _30815_ (.A(_08941_), .B(_08942_), .Y(_01480_));
NAND_g _30816_ (.A(_11371_), .B(_08929_), .Y(_08943_));
NAND_g _30817_ (.A(cpuregs_2[6]), .B(_08930_), .Y(_08944_));
NAND_g _30818_ (.A(_08943_), .B(_08944_), .Y(_01481_));
NAND_g _30819_ (.A(_11384_), .B(_08929_), .Y(_08945_));
NAND_g _30820_ (.A(cpuregs_2[7]), .B(_08930_), .Y(_08946_));
NAND_g _30821_ (.A(_08945_), .B(_08946_), .Y(_01482_));
NAND_g _30822_ (.A(_11397_), .B(_08929_), .Y(_08947_));
NAND_g _30823_ (.A(cpuregs_2[8]), .B(_08930_), .Y(_08948_));
NAND_g _30824_ (.A(_08947_), .B(_08948_), .Y(_01483_));
NAND_g _30825_ (.A(_11410_), .B(_08929_), .Y(_08949_));
NAND_g _30826_ (.A(cpuregs_2[9]), .B(_08930_), .Y(_08950_));
NAND_g _30827_ (.A(_08949_), .B(_08950_), .Y(_01484_));
NAND_g _30828_ (.A(_11423_), .B(_08929_), .Y(_08951_));
NAND_g _30829_ (.A(cpuregs_2[10]), .B(_08930_), .Y(_08952_));
NAND_g _30830_ (.A(_08951_), .B(_08952_), .Y(_01485_));
NAND_g _30831_ (.A(_11436_), .B(_08929_), .Y(_08953_));
NAND_g _30832_ (.A(cpuregs_2[11]), .B(_08930_), .Y(_08954_));
NAND_g _30833_ (.A(_08953_), .B(_08954_), .Y(_01486_));
NAND_g _30834_ (.A(_11449_), .B(_08929_), .Y(_08955_));
NAND_g _30835_ (.A(cpuregs_2[12]), .B(_08930_), .Y(_08956_));
NAND_g _30836_ (.A(_08955_), .B(_08956_), .Y(_01487_));
NAND_g _30837_ (.A(_11462_), .B(_08929_), .Y(_08957_));
NAND_g _30838_ (.A(cpuregs_2[13]), .B(_08930_), .Y(_08958_));
NAND_g _30839_ (.A(_08957_), .B(_08958_), .Y(_01488_));
NAND_g _30840_ (.A(_11475_), .B(_08929_), .Y(_08959_));
NAND_g _30841_ (.A(cpuregs_2[14]), .B(_08930_), .Y(_08960_));
NAND_g _30842_ (.A(_08959_), .B(_08960_), .Y(_01489_));
NAND_g _30843_ (.A(_11488_), .B(_08929_), .Y(_08961_));
NAND_g _30844_ (.A(cpuregs_2[15]), .B(_08930_), .Y(_08962_));
NAND_g _30845_ (.A(_08961_), .B(_08962_), .Y(_01490_));
NAND_g _30846_ (.A(_11501_), .B(_08929_), .Y(_08963_));
NAND_g _30847_ (.A(cpuregs_2[16]), .B(_08930_), .Y(_08964_));
NAND_g _30848_ (.A(_08963_), .B(_08964_), .Y(_01491_));
NOR_g _30849_ (.A(cpuregs_2[17]), .B(_08929_), .Y(_08965_));
NOR_g _30850_ (.A(_11514_), .B(_08930_), .Y(_08966_));
NOR_g _30851_ (.A(_08965_), .B(_08966_), .Y(_01492_));
NAND_g _30852_ (.A(_11527_), .B(_08929_), .Y(_08967_));
NAND_g _30853_ (.A(cpuregs_2[18]), .B(_08930_), .Y(_08968_));
NAND_g _30854_ (.A(_08967_), .B(_08968_), .Y(_01493_));
NAND_g _30855_ (.A(_11540_), .B(_08929_), .Y(_08969_));
NAND_g _30856_ (.A(cpuregs_2[19]), .B(_08930_), .Y(_08970_));
NAND_g _30857_ (.A(_08969_), .B(_08970_), .Y(_01494_));
NAND_g _30858_ (.A(_11553_), .B(_08929_), .Y(_08971_));
NAND_g _30859_ (.A(cpuregs_2[20]), .B(_08930_), .Y(_08972_));
NAND_g _30860_ (.A(_08971_), .B(_08972_), .Y(_01495_));
NAND_g _30861_ (.A(_11566_), .B(_08929_), .Y(_08973_));
NAND_g _30862_ (.A(cpuregs_2[21]), .B(_08930_), .Y(_08974_));
NAND_g _30863_ (.A(_08973_), .B(_08974_), .Y(_01496_));
NAND_g _30864_ (.A(_11579_), .B(_08929_), .Y(_08975_));
NAND_g _30865_ (.A(cpuregs_2[22]), .B(_08930_), .Y(_08976_));
NAND_g _30866_ (.A(_08975_), .B(_08976_), .Y(_01497_));
NAND_g _30867_ (.A(_11592_), .B(_08929_), .Y(_08977_));
NAND_g _30868_ (.A(cpuregs_2[23]), .B(_08930_), .Y(_08978_));
NAND_g _30869_ (.A(_08977_), .B(_08978_), .Y(_01498_));
NAND_g _30870_ (.A(_11605_), .B(_08929_), .Y(_08979_));
NAND_g _30871_ (.A(cpuregs_2[24]), .B(_08930_), .Y(_08980_));
NAND_g _30872_ (.A(_08979_), .B(_08980_), .Y(_01499_));
NAND_g _30873_ (.A(_11618_), .B(_08929_), .Y(_08981_));
NAND_g _30874_ (.A(cpuregs_2[25]), .B(_08930_), .Y(_08982_));
NAND_g _30875_ (.A(_08981_), .B(_08982_), .Y(_01500_));
NAND_g _30876_ (.A(_11631_), .B(_08929_), .Y(_08983_));
NAND_g _30877_ (.A(cpuregs_2[26]), .B(_08930_), .Y(_08984_));
NAND_g _30878_ (.A(_08983_), .B(_08984_), .Y(_01501_));
NAND_g _30879_ (.A(_11644_), .B(_08929_), .Y(_08985_));
NAND_g _30880_ (.A(cpuregs_2[27]), .B(_08930_), .Y(_08986_));
NAND_g _30881_ (.A(_08985_), .B(_08986_), .Y(_01502_));
NAND_g _30882_ (.A(_11657_), .B(_08929_), .Y(_08987_));
NAND_g _30883_ (.A(cpuregs_2[28]), .B(_08930_), .Y(_08988_));
NAND_g _30884_ (.A(_08987_), .B(_08988_), .Y(_01503_));
NAND_g _30885_ (.A(_11670_), .B(_08929_), .Y(_08989_));
NAND_g _30886_ (.A(cpuregs_2[29]), .B(_08930_), .Y(_08990_));
NAND_g _30887_ (.A(_08989_), .B(_08990_), .Y(_01504_));
NAND_g _30888_ (.A(_11683_), .B(_08929_), .Y(_08991_));
NAND_g _30889_ (.A(cpuregs_2[30]), .B(_08930_), .Y(_08992_));
NAND_g _30890_ (.A(_08991_), .B(_08992_), .Y(_01505_));
NAND_g _30891_ (.A(_11695_), .B(_08929_), .Y(_08993_));
NAND_g _30892_ (.A(cpuregs_2[31]), .B(_08930_), .Y(_08994_));
NAND_g _30893_ (.A(_08993_), .B(_08994_), .Y(_01506_));
AND_g _30894_ (.A(_11932_), .B(_02634_), .Y(_08995_));
NAND_g _30895_ (.A(_11932_), .B(_02634_), .Y(_08996_));
NAND_g _30896_ (.A(cpuregs_23[0]), .B(_08996_), .Y(_08997_));
NAND_g _30897_ (.A(_11301_), .B(_08995_), .Y(_08998_));
NAND_g _30898_ (.A(_08997_), .B(_08998_), .Y(_01507_));
NAND_g _30899_ (.A(cpuregs_23[1]), .B(_08996_), .Y(_08999_));
NAND_g _30900_ (.A(_11310_), .B(_08995_), .Y(_09000_));
NAND_g _30901_ (.A(_08999_), .B(_09000_), .Y(_01508_));
NAND_g _30902_ (.A(cpuregs_23[2]), .B(_08996_), .Y(_09001_));
NAND_g _30903_ (.A(_11319_), .B(_08995_), .Y(_09002_));
NAND_g _30904_ (.A(_09001_), .B(_09002_), .Y(_01509_));
NAND_g _30905_ (.A(cpuregs_23[3]), .B(_08996_), .Y(_09003_));
NAND_g _30906_ (.A(_11332_), .B(_08995_), .Y(_09004_));
NAND_g _30907_ (.A(_09003_), .B(_09004_), .Y(_01510_));
NAND_g _30908_ (.A(_11345_), .B(_08995_), .Y(_09005_));
NAND_g _30909_ (.A(cpuregs_23[4]), .B(_08996_), .Y(_09006_));
NAND_g _30910_ (.A(_09005_), .B(_09006_), .Y(_01511_));
NAND_g _30911_ (.A(cpuregs_23[5]), .B(_08996_), .Y(_09007_));
NAND_g _30912_ (.A(_11358_), .B(_08995_), .Y(_09008_));
NAND_g _30913_ (.A(_09007_), .B(_09008_), .Y(_01512_));
NAND_g _30914_ (.A(cpuregs_23[6]), .B(_08996_), .Y(_09009_));
NAND_g _30915_ (.A(_11371_), .B(_08995_), .Y(_09010_));
NAND_g _30916_ (.A(_09009_), .B(_09010_), .Y(_01513_));
NAND_g _30917_ (.A(cpuregs_23[7]), .B(_08996_), .Y(_09011_));
NAND_g _30918_ (.A(_11384_), .B(_08995_), .Y(_09012_));
NAND_g _30919_ (.A(_09011_), .B(_09012_), .Y(_01514_));
NAND_g _30920_ (.A(_11397_), .B(_08995_), .Y(_09013_));
NAND_g _30921_ (.A(cpuregs_23[8]), .B(_08996_), .Y(_09014_));
NAND_g _30922_ (.A(_09013_), .B(_09014_), .Y(_01515_));
NAND_g _30923_ (.A(cpuregs_23[9]), .B(_08996_), .Y(_09015_));
NAND_g _30924_ (.A(_11410_), .B(_08995_), .Y(_09016_));
NAND_g _30925_ (.A(_09015_), .B(_09016_), .Y(_01516_));
NAND_g _30926_ (.A(cpuregs_23[10]), .B(_08996_), .Y(_09017_));
NAND_g _30927_ (.A(_11423_), .B(_08995_), .Y(_09018_));
NAND_g _30928_ (.A(_09017_), .B(_09018_), .Y(_01517_));
NAND_g _30929_ (.A(cpuregs_23[11]), .B(_08996_), .Y(_09019_));
NAND_g _30930_ (.A(_11436_), .B(_08995_), .Y(_09020_));
NAND_g _30931_ (.A(_09019_), .B(_09020_), .Y(_01518_));
NAND_g _30932_ (.A(cpuregs_23[12]), .B(_08996_), .Y(_09021_));
NAND_g _30933_ (.A(_11449_), .B(_08995_), .Y(_09022_));
NAND_g _30934_ (.A(_09021_), .B(_09022_), .Y(_01519_));
NAND_g _30935_ (.A(_11462_), .B(_08995_), .Y(_09023_));
NAND_g _30936_ (.A(cpuregs_23[13]), .B(_08996_), .Y(_09024_));
NAND_g _30937_ (.A(_09023_), .B(_09024_), .Y(_01520_));
NAND_g _30938_ (.A(cpuregs_23[14]), .B(_08996_), .Y(_09025_));
NAND_g _30939_ (.A(_11475_), .B(_08995_), .Y(_09026_));
NAND_g _30940_ (.A(_09025_), .B(_09026_), .Y(_01521_));
NAND_g _30941_ (.A(cpuregs_23[15]), .B(_08996_), .Y(_09027_));
NAND_g _30942_ (.A(_11488_), .B(_08995_), .Y(_09028_));
NAND_g _30943_ (.A(_09027_), .B(_09028_), .Y(_01522_));
NAND_g _30944_ (.A(cpuregs_23[16]), .B(_08996_), .Y(_09029_));
NAND_g _30945_ (.A(_11501_), .B(_08995_), .Y(_09030_));
NAND_g _30946_ (.A(_09029_), .B(_09030_), .Y(_01523_));
AND_g _30947_ (.A(_11184_), .B(_08996_), .Y(_09031_));
NOR_g _30948_ (.A(_11514_), .B(_08996_), .Y(_09032_));
NOR_g _30949_ (.A(_09031_), .B(_09032_), .Y(_01524_));
NAND_g _30950_ (.A(_11527_), .B(_08995_), .Y(_09033_));
NAND_g _30951_ (.A(cpuregs_23[18]), .B(_08996_), .Y(_09034_));
NAND_g _30952_ (.A(_09033_), .B(_09034_), .Y(_01525_));
NAND_g _30953_ (.A(_11540_), .B(_08995_), .Y(_09035_));
NAND_g _30954_ (.A(cpuregs_23[19]), .B(_08996_), .Y(_09036_));
NAND_g _30955_ (.A(_09035_), .B(_09036_), .Y(_01526_));
NAND_g _30956_ (.A(_11553_), .B(_08995_), .Y(_09037_));
NAND_g _30957_ (.A(cpuregs_23[20]), .B(_08996_), .Y(_09038_));
NAND_g _30958_ (.A(_09037_), .B(_09038_), .Y(_01527_));
NAND_g _30959_ (.A(_11566_), .B(_08995_), .Y(_09039_));
NAND_g _30960_ (.A(cpuregs_23[21]), .B(_08996_), .Y(_09040_));
NAND_g _30961_ (.A(_09039_), .B(_09040_), .Y(_01528_));
NAND_g _30962_ (.A(_11579_), .B(_08995_), .Y(_09041_));
NAND_g _30963_ (.A(cpuregs_23[22]), .B(_08996_), .Y(_09042_));
NAND_g _30964_ (.A(_09041_), .B(_09042_), .Y(_01529_));
NAND_g _30965_ (.A(_11592_), .B(_08995_), .Y(_09043_));
NAND_g _30966_ (.A(cpuregs_23[23]), .B(_08996_), .Y(_09044_));
NAND_g _30967_ (.A(_09043_), .B(_09044_), .Y(_01530_));
NAND_g _30968_ (.A(_11605_), .B(_08995_), .Y(_09045_));
NAND_g _30969_ (.A(cpuregs_23[24]), .B(_08996_), .Y(_09046_));
NAND_g _30970_ (.A(_09045_), .B(_09046_), .Y(_01531_));
NAND_g _30971_ (.A(_11618_), .B(_08995_), .Y(_09047_));
NAND_g _30972_ (.A(cpuregs_23[25]), .B(_08996_), .Y(_09048_));
NAND_g _30973_ (.A(_09047_), .B(_09048_), .Y(_01532_));
NAND_g _30974_ (.A(_11631_), .B(_08995_), .Y(_09049_));
NAND_g _30975_ (.A(cpuregs_23[26]), .B(_08996_), .Y(_09050_));
NAND_g _30976_ (.A(_09049_), .B(_09050_), .Y(_01533_));
NAND_g _30977_ (.A(_11644_), .B(_08995_), .Y(_09051_));
NAND_g _30978_ (.A(cpuregs_23[27]), .B(_08996_), .Y(_09052_));
NAND_g _30979_ (.A(_09051_), .B(_09052_), .Y(_01534_));
NAND_g _30980_ (.A(_11657_), .B(_08995_), .Y(_09053_));
NAND_g _30981_ (.A(cpuregs_23[28]), .B(_08996_), .Y(_09054_));
NAND_g _30982_ (.A(_09053_), .B(_09054_), .Y(_01535_));
NAND_g _30983_ (.A(_11670_), .B(_08995_), .Y(_09055_));
NAND_g _30984_ (.A(cpuregs_23[29]), .B(_08996_), .Y(_09056_));
NAND_g _30985_ (.A(_09055_), .B(_09056_), .Y(_01536_));
NAND_g _30986_ (.A(_11683_), .B(_08995_), .Y(_09057_));
NAND_g _30987_ (.A(cpuregs_23[30]), .B(_08996_), .Y(_09058_));
NAND_g _30988_ (.A(_09057_), .B(_09058_), .Y(_01537_));
NAND_g _30989_ (.A(_11695_), .B(_08995_), .Y(_09059_));
NAND_g _30990_ (.A(cpuregs_23[31]), .B(_08996_), .Y(_09060_));
NAND_g _30991_ (.A(_09059_), .B(_09060_), .Y(_01538_));
AND_g _30992_ (.A(_02634_), .B(_04359_), .Y(_09061_));
NAND_g _30993_ (.A(_02634_), .B(_04359_), .Y(_09062_));
NAND_g _30994_ (.A(_11301_), .B(_09061_), .Y(_09063_));
NAND_g _30995_ (.A(cpuregs_20[0]), .B(_09062_), .Y(_09064_));
NAND_g _30996_ (.A(_09063_), .B(_09064_), .Y(_01539_));
NAND_g _30997_ (.A(cpuregs_20[1]), .B(_09062_), .Y(_09065_));
NAND_g _30998_ (.A(_11310_), .B(_09061_), .Y(_09066_));
NAND_g _30999_ (.A(_09065_), .B(_09066_), .Y(_01540_));
NAND_g _31000_ (.A(cpuregs_20[2]), .B(_09062_), .Y(_09067_));
NAND_g _31001_ (.A(_11319_), .B(_09061_), .Y(_09068_));
NAND_g _31002_ (.A(_09067_), .B(_09068_), .Y(_01541_));
NAND_g _31003_ (.A(_11332_), .B(_09061_), .Y(_09069_));
NAND_g _31004_ (.A(cpuregs_20[3]), .B(_09062_), .Y(_09070_));
NAND_g _31005_ (.A(_09069_), .B(_09070_), .Y(_01542_));
NAND_g _31006_ (.A(cpuregs_20[4]), .B(_09062_), .Y(_09071_));
NAND_g _31007_ (.A(_11345_), .B(_09061_), .Y(_09072_));
NAND_g _31008_ (.A(_09071_), .B(_09072_), .Y(_01543_));
NAND_g _31009_ (.A(cpuregs_20[5]), .B(_09062_), .Y(_09073_));
NAND_g _31010_ (.A(_11358_), .B(_09061_), .Y(_09074_));
NAND_g _31011_ (.A(_09073_), .B(_09074_), .Y(_01544_));
NAND_g _31012_ (.A(_11371_), .B(_09061_), .Y(_09075_));
NAND_g _31013_ (.A(cpuregs_20[6]), .B(_09062_), .Y(_09076_));
NAND_g _31014_ (.A(_09075_), .B(_09076_), .Y(_01545_));
NAND_g _31015_ (.A(cpuregs_20[7]), .B(_09062_), .Y(_09077_));
NAND_g _31016_ (.A(_11384_), .B(_09061_), .Y(_09078_));
NAND_g _31017_ (.A(_09077_), .B(_09078_), .Y(_01546_));
NAND_g _31018_ (.A(cpuregs_20[8]), .B(_09062_), .Y(_09079_));
NAND_g _31019_ (.A(_11397_), .B(_09061_), .Y(_09080_));
NAND_g _31020_ (.A(_09079_), .B(_09080_), .Y(_01547_));
NAND_g _31021_ (.A(cpuregs_20[9]), .B(_09062_), .Y(_09081_));
NAND_g _31022_ (.A(_11410_), .B(_09061_), .Y(_09082_));
NAND_g _31023_ (.A(_09081_), .B(_09082_), .Y(_01548_));
NAND_g _31024_ (.A(cpuregs_20[10]), .B(_09062_), .Y(_09083_));
NAND_g _31025_ (.A(_11423_), .B(_09061_), .Y(_09084_));
NAND_g _31026_ (.A(_09083_), .B(_09084_), .Y(_01549_));
NAND_g _31027_ (.A(cpuregs_20[11]), .B(_09062_), .Y(_09085_));
NAND_g _31028_ (.A(_11436_), .B(_09061_), .Y(_09086_));
NAND_g _31029_ (.A(_09085_), .B(_09086_), .Y(_01550_));
NAND_g _31030_ (.A(_11449_), .B(_09061_), .Y(_09087_));
NAND_g _31031_ (.A(cpuregs_20[12]), .B(_09062_), .Y(_09088_));
NAND_g _31032_ (.A(_09087_), .B(_09088_), .Y(_01551_));
NAND_g _31033_ (.A(cpuregs_20[13]), .B(_09062_), .Y(_09089_));
NAND_g _31034_ (.A(_11462_), .B(_09061_), .Y(_09090_));
NAND_g _31035_ (.A(_09089_), .B(_09090_), .Y(_01552_));
NAND_g _31036_ (.A(_11475_), .B(_09061_), .Y(_09091_));
NAND_g _31037_ (.A(cpuregs_20[14]), .B(_09062_), .Y(_09092_));
NAND_g _31038_ (.A(_09091_), .B(_09092_), .Y(_01553_));
NAND_g _31039_ (.A(cpuregs_20[15]), .B(_09062_), .Y(_09093_));
NAND_g _31040_ (.A(_11488_), .B(_09061_), .Y(_09094_));
NAND_g _31041_ (.A(_09093_), .B(_09094_), .Y(_01554_));
NAND_g _31042_ (.A(cpuregs_20[16]), .B(_09062_), .Y(_09095_));
NAND_g _31043_ (.A(_11501_), .B(_09061_), .Y(_09096_));
NAND_g _31044_ (.A(_09095_), .B(_09096_), .Y(_01555_));
AND_g _31045_ (.A(_11198_), .B(_09062_), .Y(_09097_));
NOR_g _31046_ (.A(_11514_), .B(_09062_), .Y(_09098_));
NOR_g _31047_ (.A(_09097_), .B(_09098_), .Y(_01556_));
NAND_g _31048_ (.A(_11527_), .B(_09061_), .Y(_09099_));
NAND_g _31049_ (.A(cpuregs_20[18]), .B(_09062_), .Y(_09100_));
NAND_g _31050_ (.A(_09099_), .B(_09100_), .Y(_01557_));
NAND_g _31051_ (.A(cpuregs_20[19]), .B(_09062_), .Y(_09101_));
NAND_g _31052_ (.A(_11540_), .B(_09061_), .Y(_09102_));
NAND_g _31053_ (.A(_09101_), .B(_09102_), .Y(_01558_));
NAND_g _31054_ (.A(_11553_), .B(_09061_), .Y(_09103_));
NAND_g _31055_ (.A(cpuregs_20[20]), .B(_09062_), .Y(_09104_));
NAND_g _31056_ (.A(_09103_), .B(_09104_), .Y(_01559_));
NAND_g _31057_ (.A(cpuregs_20[21]), .B(_09062_), .Y(_09105_));
NAND_g _31058_ (.A(_11566_), .B(_09061_), .Y(_09106_));
NAND_g _31059_ (.A(_09105_), .B(_09106_), .Y(_01560_));
NAND_g _31060_ (.A(cpuregs_20[22]), .B(_09062_), .Y(_09107_));
NAND_g _31061_ (.A(_11579_), .B(_09061_), .Y(_09108_));
NAND_g _31062_ (.A(_09107_), .B(_09108_), .Y(_01561_));
NAND_g _31063_ (.A(cpuregs_20[23]), .B(_09062_), .Y(_09109_));
NAND_g _31064_ (.A(_11592_), .B(_09061_), .Y(_09110_));
NAND_g _31065_ (.A(_09109_), .B(_09110_), .Y(_01562_));
NAND_g _31066_ (.A(cpuregs_20[24]), .B(_09062_), .Y(_09111_));
NAND_g _31067_ (.A(_11605_), .B(_09061_), .Y(_09112_));
NAND_g _31068_ (.A(_09111_), .B(_09112_), .Y(_01563_));
NAND_g _31069_ (.A(cpuregs_20[25]), .B(_09062_), .Y(_09113_));
NAND_g _31070_ (.A(_11618_), .B(_09061_), .Y(_09114_));
NAND_g _31071_ (.A(_09113_), .B(_09114_), .Y(_01564_));
NAND_g _31072_ (.A(cpuregs_20[26]), .B(_09062_), .Y(_09115_));
NAND_g _31073_ (.A(_11631_), .B(_09061_), .Y(_09116_));
NAND_g _31074_ (.A(_09115_), .B(_09116_), .Y(_01565_));
NAND_g _31075_ (.A(cpuregs_20[27]), .B(_09062_), .Y(_09117_));
NAND_g _31076_ (.A(_11644_), .B(_09061_), .Y(_09118_));
NAND_g _31077_ (.A(_09117_), .B(_09118_), .Y(_01566_));
NAND_g _31078_ (.A(cpuregs_20[28]), .B(_09062_), .Y(_09119_));
NAND_g _31079_ (.A(_11657_), .B(_09061_), .Y(_09120_));
NAND_g _31080_ (.A(_09119_), .B(_09120_), .Y(_01567_));
NAND_g _31081_ (.A(cpuregs_20[29]), .B(_09062_), .Y(_09121_));
NAND_g _31082_ (.A(_11670_), .B(_09061_), .Y(_09122_));
NAND_g _31083_ (.A(_09121_), .B(_09122_), .Y(_01568_));
NAND_g _31084_ (.A(cpuregs_20[30]), .B(_09062_), .Y(_09123_));
NAND_g _31085_ (.A(_11683_), .B(_09061_), .Y(_09124_));
NAND_g _31086_ (.A(_09123_), .B(_09124_), .Y(_01569_));
NAND_g _31087_ (.A(cpuregs_20[31]), .B(_09062_), .Y(_09125_));
NAND_g _31088_ (.A(_11695_), .B(_09061_), .Y(_09126_));
NAND_g _31089_ (.A(_09125_), .B(_09126_), .Y(_01570_));
AND_g _31090_ (.A(_11836_), .B(_11932_), .Y(_09127_));
NAND_g _31091_ (.A(_11836_), .B(_11932_), .Y(_09128_));
NAND_g _31092_ (.A(cpuregs_19[0]), .B(_09128_), .Y(_09129_));
NAND_g _31093_ (.A(_11301_), .B(_09127_), .Y(_09130_));
NAND_g _31094_ (.A(_09129_), .B(_09130_), .Y(_01571_));
NAND_g _31095_ (.A(cpuregs_19[1]), .B(_09128_), .Y(_09131_));
NAND_g _31096_ (.A(_11310_), .B(_09127_), .Y(_09132_));
NAND_g _31097_ (.A(_09131_), .B(_09132_), .Y(_01572_));
NAND_g _31098_ (.A(cpuregs_19[2]), .B(_09128_), .Y(_09133_));
NAND_g _31099_ (.A(_11319_), .B(_09127_), .Y(_09134_));
NAND_g _31100_ (.A(_09133_), .B(_09134_), .Y(_01573_));
NAND_g _31101_ (.A(cpuregs_19[3]), .B(_09128_), .Y(_09135_));
NAND_g _31102_ (.A(_11332_), .B(_09127_), .Y(_09136_));
NAND_g _31103_ (.A(_09135_), .B(_09136_), .Y(_01574_));
NAND_g _31104_ (.A(cpuregs_19[4]), .B(_09128_), .Y(_09137_));
NAND_g _31105_ (.A(_11345_), .B(_09127_), .Y(_09138_));
NAND_g _31106_ (.A(_09137_), .B(_09138_), .Y(_01575_));
NAND_g _31107_ (.A(cpuregs_19[5]), .B(_09128_), .Y(_09139_));
NAND_g _31108_ (.A(_11358_), .B(_09127_), .Y(_09140_));
NAND_g _31109_ (.A(_09139_), .B(_09140_), .Y(_01576_));
NAND_g _31110_ (.A(cpuregs_19[6]), .B(_09128_), .Y(_09141_));
NAND_g _31111_ (.A(_11371_), .B(_09127_), .Y(_09142_));
NAND_g _31112_ (.A(_09141_), .B(_09142_), .Y(_01577_));
NAND_g _31113_ (.A(cpuregs_19[7]), .B(_09128_), .Y(_09143_));
NAND_g _31114_ (.A(_11384_), .B(_09127_), .Y(_09144_));
NAND_g _31115_ (.A(_09143_), .B(_09144_), .Y(_01578_));
NAND_g _31116_ (.A(cpuregs_19[8]), .B(_09128_), .Y(_09145_));
NAND_g _31117_ (.A(_11397_), .B(_09127_), .Y(_09146_));
NAND_g _31118_ (.A(_09145_), .B(_09146_), .Y(_01579_));
NAND_g _31119_ (.A(cpuregs_19[9]), .B(_09128_), .Y(_09147_));
NAND_g _31120_ (.A(_11410_), .B(_09127_), .Y(_09148_));
NAND_g _31121_ (.A(_09147_), .B(_09148_), .Y(_01580_));
NAND_g _31122_ (.A(cpuregs_19[10]), .B(_09128_), .Y(_09149_));
NAND_g _31123_ (.A(_11423_), .B(_09127_), .Y(_09150_));
NAND_g _31124_ (.A(_09149_), .B(_09150_), .Y(_01581_));
NAND_g _31125_ (.A(cpuregs_19[11]), .B(_09128_), .Y(_09151_));
NAND_g _31126_ (.A(_11436_), .B(_09127_), .Y(_09152_));
NAND_g _31127_ (.A(_09151_), .B(_09152_), .Y(_01582_));
NAND_g _31128_ (.A(cpuregs_19[12]), .B(_09128_), .Y(_09153_));
NAND_g _31129_ (.A(_11449_), .B(_09127_), .Y(_09154_));
NAND_g _31130_ (.A(_09153_), .B(_09154_), .Y(_01583_));
NAND_g _31131_ (.A(cpuregs_19[13]), .B(_09128_), .Y(_09155_));
NAND_g _31132_ (.A(_11462_), .B(_09127_), .Y(_09156_));
NAND_g _31133_ (.A(_09155_), .B(_09156_), .Y(_01584_));
NAND_g _31134_ (.A(cpuregs_19[14]), .B(_09128_), .Y(_09157_));
NAND_g _31135_ (.A(_11475_), .B(_09127_), .Y(_09158_));
NAND_g _31136_ (.A(_09157_), .B(_09158_), .Y(_01585_));
NAND_g _31137_ (.A(cpuregs_19[15]), .B(_09128_), .Y(_09159_));
NAND_g _31138_ (.A(_11488_), .B(_09127_), .Y(_09160_));
NAND_g _31139_ (.A(_09159_), .B(_09160_), .Y(_01586_));
NAND_g _31140_ (.A(cpuregs_19[16]), .B(_09128_), .Y(_09161_));
NAND_g _31141_ (.A(_11501_), .B(_09127_), .Y(_09162_));
NAND_g _31142_ (.A(_09161_), .B(_09162_), .Y(_01587_));
NOR_g _31143_ (.A(cpuregs_19[17]), .B(_09127_), .Y(_09163_));
NOR_g _31144_ (.A(_11514_), .B(_09128_), .Y(_09164_));
NOR_g _31145_ (.A(_09163_), .B(_09164_), .Y(_01588_));
NAND_g _31146_ (.A(_11527_), .B(_09127_), .Y(_09165_));
NAND_g _31147_ (.A(cpuregs_19[18]), .B(_09128_), .Y(_09166_));
NAND_g _31148_ (.A(_09165_), .B(_09166_), .Y(_01589_));
NAND_g _31149_ (.A(_11540_), .B(_09127_), .Y(_09167_));
NAND_g _31150_ (.A(cpuregs_19[19]), .B(_09128_), .Y(_09168_));
NAND_g _31151_ (.A(_09167_), .B(_09168_), .Y(_01590_));
NAND_g _31152_ (.A(_11553_), .B(_09127_), .Y(_09169_));
NAND_g _31153_ (.A(cpuregs_19[20]), .B(_09128_), .Y(_09170_));
NAND_g _31154_ (.A(_09169_), .B(_09170_), .Y(_01591_));
NAND_g _31155_ (.A(_11566_), .B(_09127_), .Y(_09171_));
NAND_g _31156_ (.A(cpuregs_19[21]), .B(_09128_), .Y(_09172_));
NAND_g _31157_ (.A(_09171_), .B(_09172_), .Y(_01592_));
NAND_g _31158_ (.A(_11579_), .B(_09127_), .Y(_09173_));
NAND_g _31159_ (.A(cpuregs_19[22]), .B(_09128_), .Y(_09174_));
NAND_g _31160_ (.A(_09173_), .B(_09174_), .Y(_01593_));
NAND_g _31161_ (.A(_11592_), .B(_09127_), .Y(_09175_));
NAND_g _31162_ (.A(cpuregs_19[23]), .B(_09128_), .Y(_09176_));
NAND_g _31163_ (.A(_09175_), .B(_09176_), .Y(_01594_));
NAND_g _31164_ (.A(_11605_), .B(_09127_), .Y(_09177_));
NAND_g _31165_ (.A(cpuregs_19[24]), .B(_09128_), .Y(_09178_));
NAND_g _31166_ (.A(_09177_), .B(_09178_), .Y(_01595_));
NAND_g _31167_ (.A(_11618_), .B(_09127_), .Y(_09179_));
NAND_g _31168_ (.A(cpuregs_19[25]), .B(_09128_), .Y(_09180_));
NAND_g _31169_ (.A(_09179_), .B(_09180_), .Y(_01596_));
NAND_g _31170_ (.A(_11631_), .B(_09127_), .Y(_09181_));
NAND_g _31171_ (.A(cpuregs_19[26]), .B(_09128_), .Y(_09182_));
NAND_g _31172_ (.A(_09181_), .B(_09182_), .Y(_01597_));
NAND_g _31173_ (.A(_11644_), .B(_09127_), .Y(_09183_));
NAND_g _31174_ (.A(cpuregs_19[27]), .B(_09128_), .Y(_09184_));
NAND_g _31175_ (.A(_09183_), .B(_09184_), .Y(_01598_));
NAND_g _31176_ (.A(_11657_), .B(_09127_), .Y(_09185_));
NAND_g _31177_ (.A(cpuregs_19[28]), .B(_09128_), .Y(_09186_));
NAND_g _31178_ (.A(_09185_), .B(_09186_), .Y(_01599_));
NAND_g _31179_ (.A(_11670_), .B(_09127_), .Y(_09187_));
NAND_g _31180_ (.A(cpuregs_19[29]), .B(_09128_), .Y(_09188_));
NAND_g _31181_ (.A(_09187_), .B(_09188_), .Y(_01600_));
NAND_g _31182_ (.A(_11683_), .B(_09127_), .Y(_09189_));
NAND_g _31183_ (.A(cpuregs_19[30]), .B(_09128_), .Y(_09190_));
NAND_g _31184_ (.A(_09189_), .B(_09190_), .Y(_01601_));
NAND_g _31185_ (.A(_11695_), .B(_09127_), .Y(_09191_));
NAND_g _31186_ (.A(cpuregs_19[31]), .B(_09128_), .Y(_09192_));
NAND_g _31187_ (.A(_09191_), .B(_09192_), .Y(_01602_));
AND_g _31188_ (.A(_11836_), .B(_04359_), .Y(_09193_));
NAND_g _31189_ (.A(_11836_), .B(_04359_), .Y(_09194_));
NAND_g _31190_ (.A(cpuregs_16[0]), .B(_09194_), .Y(_09195_));
NAND_g _31191_ (.A(_11301_), .B(_09193_), .Y(_09196_));
NAND_g _31192_ (.A(_09195_), .B(_09196_), .Y(_01603_));
NAND_g _31193_ (.A(cpuregs_16[1]), .B(_09194_), .Y(_09197_));
NAND_g _31194_ (.A(_11310_), .B(_09193_), .Y(_09198_));
NAND_g _31195_ (.A(_09197_), .B(_09198_), .Y(_01604_));
NAND_g _31196_ (.A(cpuregs_16[2]), .B(_09194_), .Y(_09199_));
NAND_g _31197_ (.A(_11319_), .B(_09193_), .Y(_09200_));
NAND_g _31198_ (.A(_09199_), .B(_09200_), .Y(_01605_));
NAND_g _31199_ (.A(cpuregs_16[3]), .B(_09194_), .Y(_09201_));
NAND_g _31200_ (.A(_11332_), .B(_09193_), .Y(_09202_));
NAND_g _31201_ (.A(_09201_), .B(_09202_), .Y(_01606_));
NAND_g _31202_ (.A(cpuregs_16[4]), .B(_09194_), .Y(_09203_));
NAND_g _31203_ (.A(_11345_), .B(_09193_), .Y(_09204_));
NAND_g _31204_ (.A(_09203_), .B(_09204_), .Y(_01607_));
NAND_g _31205_ (.A(cpuregs_16[5]), .B(_09194_), .Y(_09205_));
NAND_g _31206_ (.A(_11358_), .B(_09193_), .Y(_09206_));
NAND_g _31207_ (.A(_09205_), .B(_09206_), .Y(_01608_));
NAND_g _31208_ (.A(cpuregs_16[6]), .B(_09194_), .Y(_09207_));
NAND_g _31209_ (.A(_11371_), .B(_09193_), .Y(_09208_));
NAND_g _31210_ (.A(_09207_), .B(_09208_), .Y(_01609_));
NAND_g _31211_ (.A(cpuregs_16[7]), .B(_09194_), .Y(_09209_));
NAND_g _31212_ (.A(_11384_), .B(_09193_), .Y(_09210_));
NAND_g _31213_ (.A(_09209_), .B(_09210_), .Y(_01610_));
NAND_g _31214_ (.A(cpuregs_16[8]), .B(_09194_), .Y(_09211_));
NAND_g _31215_ (.A(_11397_), .B(_09193_), .Y(_09212_));
NAND_g _31216_ (.A(_09211_), .B(_09212_), .Y(_01611_));
NAND_g _31217_ (.A(cpuregs_16[9]), .B(_09194_), .Y(_09213_));
NAND_g _31218_ (.A(_11410_), .B(_09193_), .Y(_09214_));
NAND_g _31219_ (.A(_09213_), .B(_09214_), .Y(_01612_));
NAND_g _31220_ (.A(cpuregs_16[10]), .B(_09194_), .Y(_09215_));
NAND_g _31221_ (.A(_11423_), .B(_09193_), .Y(_09216_));
NAND_g _31222_ (.A(_09215_), .B(_09216_), .Y(_01613_));
NAND_g _31223_ (.A(cpuregs_16[11]), .B(_09194_), .Y(_09217_));
NAND_g _31224_ (.A(_11436_), .B(_09193_), .Y(_09218_));
NAND_g _31225_ (.A(_09217_), .B(_09218_), .Y(_01614_));
NAND_g _31226_ (.A(cpuregs_16[12]), .B(_09194_), .Y(_09219_));
NAND_g _31227_ (.A(_11449_), .B(_09193_), .Y(_09220_));
NAND_g _31228_ (.A(_09219_), .B(_09220_), .Y(_01615_));
NAND_g _31229_ (.A(cpuregs_16[13]), .B(_09194_), .Y(_09221_));
NAND_g _31230_ (.A(_11462_), .B(_09193_), .Y(_09222_));
NAND_g _31231_ (.A(_09221_), .B(_09222_), .Y(_01616_));
NAND_g _31232_ (.A(cpuregs_16[14]), .B(_09194_), .Y(_09223_));
NAND_g _31233_ (.A(_11475_), .B(_09193_), .Y(_09224_));
NAND_g _31234_ (.A(_09223_), .B(_09224_), .Y(_01617_));
NAND_g _31235_ (.A(cpuregs_16[15]), .B(_09194_), .Y(_09225_));
NAND_g _31236_ (.A(_11488_), .B(_09193_), .Y(_09226_));
NAND_g _31237_ (.A(_09225_), .B(_09226_), .Y(_01618_));
NAND_g _31238_ (.A(cpuregs_16[16]), .B(_09194_), .Y(_09227_));
NAND_g _31239_ (.A(_11501_), .B(_09193_), .Y(_09228_));
NAND_g _31240_ (.A(_09227_), .B(_09228_), .Y(_01619_));
NOR_g _31241_ (.A(cpuregs_16[17]), .B(_09193_), .Y(_09229_));
NOR_g _31242_ (.A(_11514_), .B(_09194_), .Y(_09230_));
NOR_g _31243_ (.A(_09229_), .B(_09230_), .Y(_01620_));
NOR_g _31244_ (.A(cpuregs_16[18]), .B(_09193_), .Y(_09231_));
NOR_g _31245_ (.A(_11527_), .B(_09194_), .Y(_09232_));
NOR_g _31246_ (.A(_09231_), .B(_09232_), .Y(_01621_));
NOR_g _31247_ (.A(cpuregs_16[19]), .B(_09193_), .Y(_09233_));
NOR_g _31248_ (.A(_11540_), .B(_09194_), .Y(_09234_));
NOR_g _31249_ (.A(_09233_), .B(_09234_), .Y(_01622_));
NOR_g _31250_ (.A(cpuregs_16[20]), .B(_09193_), .Y(_09235_));
NOR_g _31251_ (.A(_11553_), .B(_09194_), .Y(_09236_));
NOR_g _31252_ (.A(_09235_), .B(_09236_), .Y(_01623_));
NOR_g _31253_ (.A(cpuregs_16[21]), .B(_09193_), .Y(_09237_));
NOR_g _31254_ (.A(_11566_), .B(_09194_), .Y(_09238_));
NOR_g _31255_ (.A(_09237_), .B(_09238_), .Y(_01624_));
NOR_g _31256_ (.A(cpuregs_16[22]), .B(_09193_), .Y(_09239_));
NOR_g _31257_ (.A(_11579_), .B(_09194_), .Y(_09240_));
NOR_g _31258_ (.A(_09239_), .B(_09240_), .Y(_01625_));
NOR_g _31259_ (.A(cpuregs_16[23]), .B(_09193_), .Y(_09241_));
NOR_g _31260_ (.A(_11592_), .B(_09194_), .Y(_09242_));
NOR_g _31261_ (.A(_09241_), .B(_09242_), .Y(_01626_));
NOR_g _31262_ (.A(cpuregs_16[24]), .B(_09193_), .Y(_09243_));
NOR_g _31263_ (.A(_11605_), .B(_09194_), .Y(_09244_));
NOR_g _31264_ (.A(_09243_), .B(_09244_), .Y(_01627_));
NOR_g _31265_ (.A(cpuregs_16[25]), .B(_09193_), .Y(_09245_));
NOR_g _31266_ (.A(_11618_), .B(_09194_), .Y(_09246_));
NOR_g _31267_ (.A(_09245_), .B(_09246_), .Y(_01628_));
NOR_g _31268_ (.A(cpuregs_16[26]), .B(_09193_), .Y(_09247_));
NOR_g _31269_ (.A(_11631_), .B(_09194_), .Y(_09248_));
NOR_g _31270_ (.A(_09247_), .B(_09248_), .Y(_01629_));
NOR_g _31271_ (.A(cpuregs_16[27]), .B(_09193_), .Y(_09249_));
NOR_g _31272_ (.A(_11644_), .B(_09194_), .Y(_09250_));
NOR_g _31273_ (.A(_09249_), .B(_09250_), .Y(_01630_));
NOR_g _31274_ (.A(cpuregs_16[28]), .B(_09193_), .Y(_09251_));
NOR_g _31275_ (.A(_11657_), .B(_09194_), .Y(_09252_));
NOR_g _31276_ (.A(_09251_), .B(_09252_), .Y(_01631_));
NOR_g _31277_ (.A(cpuregs_16[29]), .B(_09193_), .Y(_09253_));
NOR_g _31278_ (.A(_11670_), .B(_09194_), .Y(_09254_));
NOR_g _31279_ (.A(_09253_), .B(_09254_), .Y(_01632_));
NOR_g _31280_ (.A(cpuregs_16[30]), .B(_09193_), .Y(_09255_));
NOR_g _31281_ (.A(_11683_), .B(_09194_), .Y(_09256_));
NOR_g _31282_ (.A(_09255_), .B(_09256_), .Y(_01633_));
NOR_g _31283_ (.A(cpuregs_16[31]), .B(_09193_), .Y(_09257_));
NOR_g _31284_ (.A(_11695_), .B(_09194_), .Y(_09258_));
NOR_g _31285_ (.A(_09257_), .B(_09258_), .Y(_01634_));
AND_g _31286_ (.A(_11289_), .B(_04292_), .Y(_09259_));
NAND_g _31287_ (.A(_11289_), .B(_04292_), .Y(_09260_));
NAND_g _31288_ (.A(cpuregs_1[0]), .B(_09260_), .Y(_09261_));
NAND_g _31289_ (.A(_11301_), .B(_09259_), .Y(_09262_));
NAND_g _31290_ (.A(_09261_), .B(_09262_), .Y(_01635_));
NAND_g _31291_ (.A(cpuregs_1[1]), .B(_09260_), .Y(_09263_));
NAND_g _31292_ (.A(_11310_), .B(_09259_), .Y(_09264_));
NAND_g _31293_ (.A(_09263_), .B(_09264_), .Y(_01636_));
NAND_g _31294_ (.A(cpuregs_1[2]), .B(_09260_), .Y(_09265_));
NAND_g _31295_ (.A(_11319_), .B(_09259_), .Y(_09266_));
NAND_g _31296_ (.A(_09265_), .B(_09266_), .Y(_01637_));
NAND_g _31297_ (.A(cpuregs_1[3]), .B(_09260_), .Y(_09267_));
NAND_g _31298_ (.A(_11332_), .B(_09259_), .Y(_09268_));
NAND_g _31299_ (.A(_09267_), .B(_09268_), .Y(_01638_));
NAND_g _31300_ (.A(cpuregs_1[4]), .B(_09260_), .Y(_09269_));
NAND_g _31301_ (.A(_11345_), .B(_09259_), .Y(_09270_));
NAND_g _31302_ (.A(_09269_), .B(_09270_), .Y(_01639_));
NAND_g _31303_ (.A(cpuregs_1[5]), .B(_09260_), .Y(_09271_));
NAND_g _31304_ (.A(_11358_), .B(_09259_), .Y(_09272_));
NAND_g _31305_ (.A(_09271_), .B(_09272_), .Y(_01640_));
NAND_g _31306_ (.A(cpuregs_1[6]), .B(_09260_), .Y(_09273_));
NAND_g _31307_ (.A(_11371_), .B(_09259_), .Y(_09274_));
NAND_g _31308_ (.A(_09273_), .B(_09274_), .Y(_01641_));
NAND_g _31309_ (.A(cpuregs_1[7]), .B(_09260_), .Y(_09275_));
NAND_g _31310_ (.A(_11384_), .B(_09259_), .Y(_09276_));
NAND_g _31311_ (.A(_09275_), .B(_09276_), .Y(_01642_));
NAND_g _31312_ (.A(cpuregs_1[8]), .B(_09260_), .Y(_09277_));
NAND_g _31313_ (.A(_11397_), .B(_09259_), .Y(_09278_));
NAND_g _31314_ (.A(_09277_), .B(_09278_), .Y(_01643_));
NAND_g _31315_ (.A(cpuregs_1[9]), .B(_09260_), .Y(_09279_));
NAND_g _31316_ (.A(_11410_), .B(_09259_), .Y(_09280_));
NAND_g _31317_ (.A(_09279_), .B(_09280_), .Y(_01644_));
NAND_g _31318_ (.A(cpuregs_1[10]), .B(_09260_), .Y(_09281_));
NAND_g _31319_ (.A(_11423_), .B(_09259_), .Y(_09282_));
NAND_g _31320_ (.A(_09281_), .B(_09282_), .Y(_01645_));
NAND_g _31321_ (.A(cpuregs_1[11]), .B(_09260_), .Y(_09283_));
NAND_g _31322_ (.A(_11436_), .B(_09259_), .Y(_09284_));
NAND_g _31323_ (.A(_09283_), .B(_09284_), .Y(_01646_));
NAND_g _31324_ (.A(cpuregs_1[12]), .B(_09260_), .Y(_09285_));
NAND_g _31325_ (.A(_11449_), .B(_09259_), .Y(_09286_));
NAND_g _31326_ (.A(_09285_), .B(_09286_), .Y(_01647_));
NAND_g _31327_ (.A(cpuregs_1[13]), .B(_09260_), .Y(_09287_));
NAND_g _31328_ (.A(_11462_), .B(_09259_), .Y(_09288_));
NAND_g _31329_ (.A(_09287_), .B(_09288_), .Y(_01648_));
NAND_g _31330_ (.A(cpuregs_1[14]), .B(_09260_), .Y(_09289_));
NAND_g _31331_ (.A(_11475_), .B(_09259_), .Y(_09290_));
NAND_g _31332_ (.A(_09289_), .B(_09290_), .Y(_01649_));
NAND_g _31333_ (.A(cpuregs_1[15]), .B(_09260_), .Y(_09291_));
NAND_g _31334_ (.A(_11488_), .B(_09259_), .Y(_09292_));
NAND_g _31335_ (.A(_09291_), .B(_09292_), .Y(_01650_));
NAND_g _31336_ (.A(cpuregs_1[16]), .B(_09260_), .Y(_09293_));
NAND_g _31337_ (.A(_11501_), .B(_09259_), .Y(_09294_));
NAND_g _31338_ (.A(_09293_), .B(_09294_), .Y(_01651_));
NOR_g _31339_ (.A(cpuregs_1[17]), .B(_09259_), .Y(_09295_));
NOR_g _31340_ (.A(_11514_), .B(_09260_), .Y(_09296_));
NOR_g _31341_ (.A(_09295_), .B(_09296_), .Y(_01652_));
NAND_g _31342_ (.A(cpuregs_1[18]), .B(_09260_), .Y(_09297_));
NAND_g _31343_ (.A(_11527_), .B(_09259_), .Y(_09298_));
NAND_g _31344_ (.A(_09297_), .B(_09298_), .Y(_01653_));
NAND_g _31345_ (.A(cpuregs_1[19]), .B(_09260_), .Y(_09299_));
NAND_g _31346_ (.A(_11540_), .B(_09259_), .Y(_09300_));
NAND_g _31347_ (.A(_09299_), .B(_09300_), .Y(_01654_));
NAND_g _31348_ (.A(cpuregs_1[20]), .B(_09260_), .Y(_09301_));
NAND_g _31349_ (.A(_11553_), .B(_09259_), .Y(_09302_));
NAND_g _31350_ (.A(_09301_), .B(_09302_), .Y(_01655_));
NAND_g _31351_ (.A(cpuregs_1[21]), .B(_09260_), .Y(_09303_));
NAND_g _31352_ (.A(_11566_), .B(_09259_), .Y(_09304_));
NAND_g _31353_ (.A(_09303_), .B(_09304_), .Y(_01656_));
NAND_g _31354_ (.A(cpuregs_1[22]), .B(_09260_), .Y(_09305_));
NAND_g _31355_ (.A(_11579_), .B(_09259_), .Y(_09306_));
NAND_g _31356_ (.A(_09305_), .B(_09306_), .Y(_01657_));
NAND_g _31357_ (.A(cpuregs_1[23]), .B(_09260_), .Y(_09307_));
NAND_g _31358_ (.A(_11592_), .B(_09259_), .Y(_09308_));
NAND_g _31359_ (.A(_09307_), .B(_09308_), .Y(_01658_));
NAND_g _31360_ (.A(cpuregs_1[24]), .B(_09260_), .Y(_09309_));
NAND_g _31361_ (.A(_11605_), .B(_09259_), .Y(_09310_));
NAND_g _31362_ (.A(_09309_), .B(_09310_), .Y(_01659_));
NAND_g _31363_ (.A(cpuregs_1[25]), .B(_09260_), .Y(_09311_));
NAND_g _31364_ (.A(_11618_), .B(_09259_), .Y(_09312_));
NAND_g _31365_ (.A(_09311_), .B(_09312_), .Y(_01660_));
NAND_g _31366_ (.A(cpuregs_1[26]), .B(_09260_), .Y(_09313_));
NAND_g _31367_ (.A(_11631_), .B(_09259_), .Y(_09314_));
NAND_g _31368_ (.A(_09313_), .B(_09314_), .Y(_01661_));
NAND_g _31369_ (.A(cpuregs_1[27]), .B(_09260_), .Y(_09315_));
NAND_g _31370_ (.A(_11644_), .B(_09259_), .Y(_09316_));
NAND_g _31371_ (.A(_09315_), .B(_09316_), .Y(_01662_));
NAND_g _31372_ (.A(cpuregs_1[28]), .B(_09260_), .Y(_09317_));
NAND_g _31373_ (.A(_11657_), .B(_09259_), .Y(_09318_));
NAND_g _31374_ (.A(_09317_), .B(_09318_), .Y(_01663_));
NAND_g _31375_ (.A(cpuregs_1[29]), .B(_09260_), .Y(_09319_));
NAND_g _31376_ (.A(_11670_), .B(_09259_), .Y(_09320_));
NAND_g _31377_ (.A(_09319_), .B(_09320_), .Y(_01664_));
NAND_g _31378_ (.A(cpuregs_1[30]), .B(_09260_), .Y(_09321_));
NAND_g _31379_ (.A(_11683_), .B(_09259_), .Y(_09322_));
NAND_g _31380_ (.A(_09321_), .B(_09322_), .Y(_01665_));
NAND_g _31381_ (.A(cpuregs_1[31]), .B(_09260_), .Y(_09323_));
NAND_g _31382_ (.A(_11695_), .B(_09259_), .Y(_09324_));
NAND_g _31383_ (.A(_09323_), .B(_09324_), .Y(_01666_));
AND_g _31384_ (.A(_11697_), .B(_11765_), .Y(_09325_));
NAND_g _31385_ (.A(_11697_), .B(_11765_), .Y(_09326_));
NAND_g _31386_ (.A(_11301_), .B(_09325_), .Y(_09327_));
NAND_g _31387_ (.A(cpuregs_10[0]), .B(_09326_), .Y(_09328_));
NAND_g _31388_ (.A(_09327_), .B(_09328_), .Y(_01667_));
NAND_g _31389_ (.A(_11310_), .B(_09325_), .Y(_09329_));
NAND_g _31390_ (.A(cpuregs_10[1]), .B(_09326_), .Y(_09330_));
NAND_g _31391_ (.A(_09329_), .B(_09330_), .Y(_01668_));
NAND_g _31392_ (.A(_11319_), .B(_09325_), .Y(_09331_));
NAND_g _31393_ (.A(cpuregs_10[2]), .B(_09326_), .Y(_09332_));
NAND_g _31394_ (.A(_09331_), .B(_09332_), .Y(_01669_));
NAND_g _31395_ (.A(_11332_), .B(_09325_), .Y(_09333_));
NAND_g _31396_ (.A(cpuregs_10[3]), .B(_09326_), .Y(_09334_));
NAND_g _31397_ (.A(_09333_), .B(_09334_), .Y(_01670_));
NAND_g _31398_ (.A(_11345_), .B(_09325_), .Y(_09335_));
NAND_g _31399_ (.A(cpuregs_10[4]), .B(_09326_), .Y(_09336_));
NAND_g _31400_ (.A(_09335_), .B(_09336_), .Y(_01671_));
NAND_g _31401_ (.A(_11358_), .B(_09325_), .Y(_09337_));
NAND_g _31402_ (.A(cpuregs_10[5]), .B(_09326_), .Y(_09338_));
NAND_g _31403_ (.A(_09337_), .B(_09338_), .Y(_01672_));
NAND_g _31404_ (.A(_11371_), .B(_09325_), .Y(_09339_));
NAND_g _31405_ (.A(cpuregs_10[6]), .B(_09326_), .Y(_09340_));
NAND_g _31406_ (.A(_09339_), .B(_09340_), .Y(_01673_));
NAND_g _31407_ (.A(_11384_), .B(_09325_), .Y(_09341_));
NAND_g _31408_ (.A(cpuregs_10[7]), .B(_09326_), .Y(_09342_));
NAND_g _31409_ (.A(_09341_), .B(_09342_), .Y(_01674_));
NAND_g _31410_ (.A(_11397_), .B(_09325_), .Y(_09343_));
NAND_g _31411_ (.A(cpuregs_10[8]), .B(_09326_), .Y(_09344_));
NAND_g _31412_ (.A(_09343_), .B(_09344_), .Y(_01675_));
NAND_g _31413_ (.A(_11410_), .B(_09325_), .Y(_09345_));
NAND_g _31414_ (.A(cpuregs_10[9]), .B(_09326_), .Y(_09346_));
NAND_g _31415_ (.A(_09345_), .B(_09346_), .Y(_01676_));
NAND_g _31416_ (.A(_11423_), .B(_09325_), .Y(_09347_));
NAND_g _31417_ (.A(cpuregs_10[10]), .B(_09326_), .Y(_09348_));
NAND_g _31418_ (.A(_09347_), .B(_09348_), .Y(_01677_));
NAND_g _31419_ (.A(_11436_), .B(_09325_), .Y(_09349_));
NAND_g _31420_ (.A(cpuregs_10[11]), .B(_09326_), .Y(_09350_));
NAND_g _31421_ (.A(_09349_), .B(_09350_), .Y(_01678_));
NAND_g _31422_ (.A(_11449_), .B(_09325_), .Y(_09351_));
NAND_g _31423_ (.A(cpuregs_10[12]), .B(_09326_), .Y(_09352_));
NAND_g _31424_ (.A(_09351_), .B(_09352_), .Y(_01679_));
NAND_g _31425_ (.A(_11462_), .B(_09325_), .Y(_09353_));
NAND_g _31426_ (.A(cpuregs_10[13]), .B(_09326_), .Y(_09354_));
NAND_g _31427_ (.A(_09353_), .B(_09354_), .Y(_01680_));
NAND_g _31428_ (.A(_11475_), .B(_09325_), .Y(_09355_));
NAND_g _31429_ (.A(cpuregs_10[14]), .B(_09326_), .Y(_09356_));
NAND_g _31430_ (.A(_09355_), .B(_09356_), .Y(_01681_));
NAND_g _31431_ (.A(_11488_), .B(_09325_), .Y(_09357_));
NAND_g _31432_ (.A(cpuregs_10[15]), .B(_09326_), .Y(_09358_));
NAND_g _31433_ (.A(_09357_), .B(_09358_), .Y(_01682_));
NOR_g _31434_ (.A(cpuregs_10[16]), .B(_09325_), .Y(_09359_));
NOR_g _31435_ (.A(_11501_), .B(_09326_), .Y(_09360_));
NOR_g _31436_ (.A(_09359_), .B(_09360_), .Y(_01683_));
NAND_g _31437_ (.A(_11514_), .B(_09325_), .Y(_09361_));
NAND_g _31438_ (.A(cpuregs_10[17]), .B(_09326_), .Y(_09362_));
NAND_g _31439_ (.A(_09361_), .B(_09362_), .Y(_01684_));
NAND_g _31440_ (.A(_11527_), .B(_09325_), .Y(_09363_));
NAND_g _31441_ (.A(cpuregs_10[18]), .B(_09326_), .Y(_09364_));
NAND_g _31442_ (.A(_09363_), .B(_09364_), .Y(_01685_));
NAND_g _31443_ (.A(_11540_), .B(_09325_), .Y(_09365_));
NAND_g _31444_ (.A(cpuregs_10[19]), .B(_09326_), .Y(_09366_));
NAND_g _31445_ (.A(_09365_), .B(_09366_), .Y(_01686_));
NAND_g _31446_ (.A(_11553_), .B(_09325_), .Y(_09367_));
NAND_g _31447_ (.A(cpuregs_10[20]), .B(_09326_), .Y(_09368_));
NAND_g _31448_ (.A(_09367_), .B(_09368_), .Y(_01687_));
NAND_g _31449_ (.A(_11566_), .B(_09325_), .Y(_09369_));
NAND_g _31450_ (.A(cpuregs_10[21]), .B(_09326_), .Y(_09370_));
NAND_g _31451_ (.A(_09369_), .B(_09370_), .Y(_01688_));
NAND_g _31452_ (.A(_11579_), .B(_09325_), .Y(_09371_));
NAND_g _31453_ (.A(cpuregs_10[22]), .B(_09326_), .Y(_09372_));
NAND_g _31454_ (.A(_09371_), .B(_09372_), .Y(_01689_));
NAND_g _31455_ (.A(_11592_), .B(_09325_), .Y(_09373_));
NAND_g _31456_ (.A(cpuregs_10[23]), .B(_09326_), .Y(_09374_));
NAND_g _31457_ (.A(_09373_), .B(_09374_), .Y(_01690_));
NAND_g _31458_ (.A(_11605_), .B(_09325_), .Y(_09375_));
NAND_g _31459_ (.A(cpuregs_10[24]), .B(_09326_), .Y(_09376_));
NAND_g _31460_ (.A(_09375_), .B(_09376_), .Y(_01691_));
NAND_g _31461_ (.A(_11618_), .B(_09325_), .Y(_09377_));
NAND_g _31462_ (.A(cpuregs_10[25]), .B(_09326_), .Y(_09378_));
NAND_g _31463_ (.A(_09377_), .B(_09378_), .Y(_01692_));
NAND_g _31464_ (.A(_11631_), .B(_09325_), .Y(_09379_));
NAND_g _31465_ (.A(cpuregs_10[26]), .B(_09326_), .Y(_09380_));
NAND_g _31466_ (.A(_09379_), .B(_09380_), .Y(_01693_));
NAND_g _31467_ (.A(_11644_), .B(_09325_), .Y(_09381_));
NAND_g _31468_ (.A(cpuregs_10[27]), .B(_09326_), .Y(_09382_));
NAND_g _31469_ (.A(_09381_), .B(_09382_), .Y(_01694_));
NAND_g _31470_ (.A(_11657_), .B(_09325_), .Y(_09383_));
NAND_g _31471_ (.A(cpuregs_10[28]), .B(_09326_), .Y(_09384_));
NAND_g _31472_ (.A(_09383_), .B(_09384_), .Y(_01695_));
NAND_g _31473_ (.A(_11670_), .B(_09325_), .Y(_09385_));
NAND_g _31474_ (.A(cpuregs_10[29]), .B(_09326_), .Y(_09386_));
NAND_g _31475_ (.A(_09385_), .B(_09386_), .Y(_01696_));
NAND_g _31476_ (.A(_11683_), .B(_09325_), .Y(_09387_));
NAND_g _31477_ (.A(cpuregs_10[30]), .B(_09326_), .Y(_09388_));
NAND_g _31478_ (.A(_09387_), .B(_09388_), .Y(_01697_));
NAND_g _31479_ (.A(_11695_), .B(_09325_), .Y(_09389_));
NAND_g _31480_ (.A(cpuregs_10[31]), .B(_09326_), .Y(_09390_));
NAND_g _31481_ (.A(_09389_), .B(_09390_), .Y(_01698_));
NOR_g _31482_ (.A(instr_slt), .B(instr_slti), .Y(_09391_));
NAND_g _31483_ (.A(_10921_), .B(_09391_), .Y(_00007_));
NOR_g _31484_ (.A(instr_sltu), .B(instr_sltiu), .Y(_09392_));
NAND_g _31485_ (.A(_10919_), .B(_09392_), .Y(_00008_));
NAND_g _31486_ (.A(is_compare), .B(_02562_), .Y(_09393_));
NAND_g _31487_ (.A(_10907_), .B(_10914_), .Y(_09394_));
NOR_g _31488_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09394_), .Y(_09395_));
NOT_g _31489_ (.A(_09395_), .Y(_09396_));
NOR_g _31490_ (.A(instr_or), .B(instr_ori), .Y(_09397_));
NOR_g _31491_ (.A(instr_and), .B(instr_andi), .Y(_09398_));
NOR_g _31492_ (.A(_02425_), .B(_09398_), .Y(_09399_));
NAND_g _31493_ (.A(_02425_), .B(_09396_), .Y(_09400_));
AND_g _31494_ (.A(_09397_), .B(_09400_), .Y(_09401_));
NOR_g _31495_ (.A(_02424_), .B(_09401_), .Y(_09402_));
NOR_g _31496_ (.A(_09399_), .B(_09402_), .Y(_09403_));
NAND_g _31497_ (.A(_09393_), .B(_09403_), .Y(alu_out[0]));
NAND_g _31498_ (.A(_10910_), .B(_02425_), .Y(_09404_));
NAND_g _31499_ (.A(instr_sub), .B(_02427_), .Y(_09405_));
AND_g _31500_ (.A(_09404_), .B(_09405_), .Y(_09406_));
XNOR_g _31501_ (.A(_02423_), .B(_09406_), .Y(_09407_));
NAND_g _31502_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09407_), .Y(_09408_));
NAND_g _31503_ (.A(_02422_), .B(_09394_), .Y(_09409_));
NOR_g _31504_ (.A(_02419_), .B(_09397_), .Y(_09410_));
NOR_g _31505_ (.A(_02421_), .B(_09398_), .Y(_09411_));
NOR_g _31506_ (.A(_09410_), .B(_09411_), .Y(_09412_));
AND_g _31507_ (.A(_09409_), .B(_09412_), .Y(_09413_));
NAND_g _31508_ (.A(_09408_), .B(_09413_), .Y(alu_out[1]));
NOR_g _31509_ (.A(_10910_), .B(_02429_), .Y(_09414_));
NOR_g _31510_ (.A(_02419_), .B(_02425_), .Y(_09415_));
NOR_g _31511_ (.A(_02420_), .B(_09415_), .Y(_09416_));
NOR_g _31512_ (.A(instr_sub), .B(_09416_), .Y(_09417_));
NOR_g _31513_ (.A(_09414_), .B(_09417_), .Y(_09418_));
XNOR_g _31514_ (.A(_02416_), .B(_09418_), .Y(_09419_));
NAND_g _31515_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09419_), .Y(_09420_));
NAND_g _31516_ (.A(_02416_), .B(_09394_), .Y(_09421_));
NOR_g _31517_ (.A(_02413_), .B(_09397_), .Y(_09422_));
NOR_g _31518_ (.A(_02415_), .B(_09398_), .Y(_09423_));
NOR_g _31519_ (.A(_09422_), .B(_09423_), .Y(_09424_));
AND_g _31520_ (.A(_09421_), .B(_09424_), .Y(_09425_));
NAND_g _31521_ (.A(_09420_), .B(_09425_), .Y(alu_out[2]));
NOR_g _31522_ (.A(_02413_), .B(_09416_), .Y(_09426_));
NOR_g _31523_ (.A(_02414_), .B(_09426_), .Y(_09427_));
NAND_g _31524_ (.A(_10910_), .B(_09427_), .Y(_09428_));
NAND_g _31525_ (.A(instr_sub), .B(_02431_), .Y(_09429_));
AND_g _31526_ (.A(_09428_), .B(_09429_), .Y(_09430_));
XNOR_g _31527_ (.A(_02545_), .B(_09430_), .Y(_09431_));
NAND_g _31528_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09431_), .Y(_09432_));
NAND_g _31529_ (.A(_02544_), .B(_09394_), .Y(_09433_));
NOR_g _31530_ (.A(_02543_), .B(_09398_), .Y(_09434_));
NOR_g _31531_ (.A(_02541_), .B(_09397_), .Y(_09435_));
NOR_g _31532_ (.A(_09434_), .B(_09435_), .Y(_09436_));
AND_g _31533_ (.A(_09433_), .B(_09436_), .Y(_09437_));
NAND_g _31534_ (.A(_09432_), .B(_09437_), .Y(alu_out[3]));
NOR_g _31535_ (.A(_02541_), .B(_09427_), .Y(_09438_));
NOR_g _31536_ (.A(_02542_), .B(_09438_), .Y(_09439_));
NAND_g _31537_ (.A(_10910_), .B(_09439_), .Y(_09440_));
NAND_g _31538_ (.A(instr_sub), .B(_02435_), .Y(_09441_));
AND_g _31539_ (.A(_09440_), .B(_09441_), .Y(_09442_));
XNOR_g _31540_ (.A(_02411_), .B(_09442_), .Y(_09443_));
NAND_g _31541_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09443_), .Y(_09444_));
NAND_g _31542_ (.A(_02410_), .B(_09394_), .Y(_09445_));
NOR_g _31543_ (.A(_02409_), .B(_09398_), .Y(_09446_));
NOR_g _31544_ (.A(_02407_), .B(_09397_), .Y(_09447_));
NOR_g _31545_ (.A(_09446_), .B(_09447_), .Y(_09448_));
AND_g _31546_ (.A(_09445_), .B(_09448_), .Y(_09449_));
NAND_g _31547_ (.A(_09444_), .B(_09449_), .Y(alu_out[4]));
NAND_g _31548_ (.A(instr_sub), .B(_02438_), .Y(_09450_));
NOR_g _31549_ (.A(_02407_), .B(_09439_), .Y(_09451_));
NOR_g _31550_ (.A(_02408_), .B(_09451_), .Y(_09452_));
NAND_g _31551_ (.A(_10910_), .B(_09452_), .Y(_09453_));
AND_g _31552_ (.A(_09450_), .B(_09453_), .Y(_09454_));
XNOR_g _31553_ (.A(_02406_), .B(_09454_), .Y(_09455_));
NAND_g _31554_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09455_), .Y(_09456_));
NAND_g _31555_ (.A(_02405_), .B(_09394_), .Y(_09457_));
NOR_g _31556_ (.A(_02403_), .B(_09397_), .Y(_09458_));
NOR_g _31557_ (.A(_02404_), .B(_09398_), .Y(_09459_));
NOR_g _31558_ (.A(_09458_), .B(_09459_), .Y(_09460_));
AND_g _31559_ (.A(_09457_), .B(_09460_), .Y(_09461_));
NAND_g _31560_ (.A(_09456_), .B(_09461_), .Y(alu_out[5]));
AND_g _31561_ (.A(_02404_), .B(_09452_), .Y(_09462_));
NOR_g _31562_ (.A(_02403_), .B(_09462_), .Y(_09463_));
NOR_g _31563_ (.A(instr_sub), .B(_09463_), .Y(_09464_));
AND_g _31564_ (.A(instr_sub), .B(_02440_), .Y(_09465_));
NOR_g _31565_ (.A(_09464_), .B(_09465_), .Y(_09466_));
XNOR_g _31566_ (.A(_02400_), .B(_09466_), .Y(_09467_));
NAND_g _31567_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09467_), .Y(_09468_));
NAND_g _31568_ (.A(_02399_), .B(_09394_), .Y(_09469_));
NOR_g _31569_ (.A(_02398_), .B(_09398_), .Y(_09470_));
NOR_g _31570_ (.A(_02396_), .B(_09397_), .Y(_09471_));
NOR_g _31571_ (.A(_09470_), .B(_09471_), .Y(_09472_));
AND_g _31572_ (.A(_09469_), .B(_09472_), .Y(_09473_));
NAND_g _31573_ (.A(_09468_), .B(_09473_), .Y(alu_out[6]));
NAND_g _31574_ (.A(_02397_), .B(_09463_), .Y(_09474_));
AND_g _31575_ (.A(_02398_), .B(_09474_), .Y(_09475_));
NOR_g _31576_ (.A(instr_sub), .B(_09475_), .Y(_09476_));
NAND_g _31577_ (.A(_02400_), .B(_02440_), .Y(_09477_));
NAND_g _31578_ (.A(instr_sub), .B(_09477_), .Y(_09478_));
NOR_g _31579_ (.A(_02443_), .B(_09478_), .Y(_09479_));
NOR_g _31580_ (.A(_09476_), .B(_09479_), .Y(_09480_));
XNOR_g _31581_ (.A(_02394_), .B(_09480_), .Y(_09481_));
NAND_g _31582_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09481_), .Y(_09482_));
NAND_g _31583_ (.A(_02394_), .B(_09394_), .Y(_09483_));
NOR_g _31584_ (.A(_02392_), .B(_09397_), .Y(_09484_));
NOR_g _31585_ (.A(_02393_), .B(_09398_), .Y(_09485_));
NOR_g _31586_ (.A(_09484_), .B(_09485_), .Y(_09486_));
AND_g _31587_ (.A(_09483_), .B(_09486_), .Y(_09487_));
NAND_g _31588_ (.A(_09482_), .B(_09487_), .Y(alu_out[7]));
AND_g _31589_ (.A(_02393_), .B(_09475_), .Y(_09488_));
NOR_g _31590_ (.A(_02392_), .B(_09488_), .Y(_09489_));
NOR_g _31591_ (.A(instr_sub), .B(_09489_), .Y(_09490_));
AND_g _31592_ (.A(instr_sub), .B(_02446_), .Y(_09491_));
NOR_g _31593_ (.A(_09490_), .B(_09491_), .Y(_09492_));
XNOR_g _31594_ (.A(_02450_), .B(_09492_), .Y(_09493_));
NAND_g _31595_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09493_), .Y(_09494_));
NAND_g _31596_ (.A(_02449_), .B(_09394_), .Y(_09495_));
NOR_g _31597_ (.A(_02448_), .B(_09398_), .Y(_09496_));
NOR_g _31598_ (.A(_02447_), .B(_09397_), .Y(_09497_));
NOR_g _31599_ (.A(_09496_), .B(_09497_), .Y(_09498_));
AND_g _31600_ (.A(_09495_), .B(_09498_), .Y(_09499_));
NAND_g _31601_ (.A(_09494_), .B(_09499_), .Y(alu_out[8]));
NOR_g _31602_ (.A(_10910_), .B(_02458_), .Y(_09500_));
NAND_g _31603_ (.A(_02451_), .B(_09500_), .Y(_09501_));
NAND_g _31604_ (.A(_02449_), .B(_09489_), .Y(_09502_));
NAND_g _31605_ (.A(_02448_), .B(_09502_), .Y(_09503_));
NAND_g _31606_ (.A(_10910_), .B(_09503_), .Y(_09504_));
AND_g _31607_ (.A(_09501_), .B(_09504_), .Y(_09505_));
XNOR_g _31608_ (.A(_02390_), .B(_09505_), .Y(_09506_));
NAND_g _31609_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09506_), .Y(_09507_));
NAND_g _31610_ (.A(_02390_), .B(_09394_), .Y(_09508_));
NOR_g _31611_ (.A(_02389_), .B(_09398_), .Y(_09509_));
NOR_g _31612_ (.A(_02388_), .B(_09397_), .Y(_09510_));
NOR_g _31613_ (.A(_09509_), .B(_09510_), .Y(_09511_));
AND_g _31614_ (.A(_09508_), .B(_09511_), .Y(_09512_));
NAND_g _31615_ (.A(_09507_), .B(_09512_), .Y(alu_out[9]));
AND_g _31616_ (.A(_02389_), .B(_02448_), .Y(_09513_));
AND_g _31617_ (.A(_09502_), .B(_09513_), .Y(_09514_));
NOR_g _31618_ (.A(_02388_), .B(_09514_), .Y(_09515_));
NAND_g _31619_ (.A(_02454_), .B(_02460_), .Y(_09516_));
AND_g _31620_ (.A(instr_sub), .B(_09516_), .Y(_09517_));
NOR_g _31621_ (.A(instr_sub), .B(_09515_), .Y(_09518_));
NOR_g _31622_ (.A(_09517_), .B(_09518_), .Y(_09519_));
XNOR_g _31623_ (.A(_02386_), .B(_09519_), .Y(_09520_));
NAND_g _31624_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09520_), .Y(_09521_));
NAND_g _31625_ (.A(_02385_), .B(_09394_), .Y(_09522_));
NOR_g _31626_ (.A(_02384_), .B(_09398_), .Y(_09523_));
NOR_g _31627_ (.A(_02383_), .B(_09397_), .Y(_09524_));
NOR_g _31628_ (.A(_09523_), .B(_09524_), .Y(_09525_));
AND_g _31629_ (.A(_09522_), .B(_09525_), .Y(_09526_));
NAND_g _31630_ (.A(_09521_), .B(_09526_), .Y(alu_out[10]));
NAND_g _31631_ (.A(_02386_), .B(_09516_), .Y(_09527_));
NAND_g _31632_ (.A(_02456_), .B(_09527_), .Y(_09528_));
NAND_g _31633_ (.A(instr_sub), .B(_09528_), .Y(_09529_));
NAND_g _31634_ (.A(_02385_), .B(_09515_), .Y(_09530_));
AND_g _31635_ (.A(_10910_), .B(_02384_), .Y(_09531_));
NAND_g _31636_ (.A(_09530_), .B(_09531_), .Y(_09532_));
AND_g _31637_ (.A(_09529_), .B(_09532_), .Y(_09533_));
XNOR_g _31638_ (.A(_02382_), .B(_09533_), .Y(_09534_));
NAND_g _31639_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09534_), .Y(_09535_));
NAND_g _31640_ (.A(_02381_), .B(_09394_), .Y(_09536_));
NOR_g _31641_ (.A(_02379_), .B(_09397_), .Y(_09537_));
NOR_g _31642_ (.A(_02380_), .B(_09398_), .Y(_09538_));
NOR_g _31643_ (.A(_09537_), .B(_09538_), .Y(_09539_));
AND_g _31644_ (.A(_09536_), .B(_09539_), .Y(_09540_));
NAND_g _31645_ (.A(_09535_), .B(_09540_), .Y(alu_out[11]));
AND_g _31646_ (.A(_02380_), .B(_02384_), .Y(_09541_));
AND_g _31647_ (.A(_09530_), .B(_09541_), .Y(_09542_));
NOR_g _31648_ (.A(_02379_), .B(_09542_), .Y(_09543_));
NOR_g _31649_ (.A(instr_sub), .B(_09543_), .Y(_09544_));
AND_g _31650_ (.A(instr_sub), .B(_02467_), .Y(_09545_));
NOR_g _31651_ (.A(_09544_), .B(_09545_), .Y(_09546_));
XNOR_g _31652_ (.A(_02377_), .B(_09546_), .Y(_09547_));
NAND_g _31653_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09547_), .Y(_09548_));
NAND_g _31654_ (.A(_02376_), .B(_09394_), .Y(_09549_));
NOR_g _31655_ (.A(_02375_), .B(_09398_), .Y(_09550_));
NOR_g _31656_ (.A(_02374_), .B(_09397_), .Y(_09551_));
NOR_g _31657_ (.A(_09550_), .B(_09551_), .Y(_09552_));
AND_g _31658_ (.A(_09549_), .B(_09552_), .Y(_09553_));
NAND_g _31659_ (.A(_09548_), .B(_09553_), .Y(alu_out[12]));
NAND_g _31660_ (.A(_02468_), .B(_02474_), .Y(_09554_));
NAND_g _31661_ (.A(instr_sub), .B(_09554_), .Y(_09555_));
NAND_g _31662_ (.A(_02376_), .B(_09543_), .Y(_09556_));
AND_g _31663_ (.A(_10910_), .B(_02375_), .Y(_09557_));
NAND_g _31664_ (.A(_09556_), .B(_09557_), .Y(_09558_));
AND_g _31665_ (.A(_09555_), .B(_09558_), .Y(_09559_));
XNOR_g _31666_ (.A(_02373_), .B(_09559_), .Y(_09560_));
NAND_g _31667_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09560_), .Y(_09561_));
NAND_g _31668_ (.A(_02372_), .B(_09394_), .Y(_09562_));
NOR_g _31669_ (.A(_02370_), .B(_09397_), .Y(_09563_));
NOR_g _31670_ (.A(_02371_), .B(_09398_), .Y(_09564_));
NOR_g _31671_ (.A(_09563_), .B(_09564_), .Y(_09565_));
AND_g _31672_ (.A(_09562_), .B(_09565_), .Y(_09566_));
NAND_g _31673_ (.A(_09561_), .B(_09566_), .Y(alu_out[13]));
AND_g _31674_ (.A(_02371_), .B(_02375_), .Y(_09567_));
AND_g _31675_ (.A(_09556_), .B(_09567_), .Y(_09568_));
NOR_g _31676_ (.A(_02370_), .B(_09568_), .Y(_09569_));
NOR_g _31677_ (.A(instr_sub), .B(_09569_), .Y(_09570_));
NAND_g _31678_ (.A(_02469_), .B(_02476_), .Y(_09571_));
AND_g _31679_ (.A(instr_sub), .B(_09571_), .Y(_09572_));
NOR_g _31680_ (.A(_09570_), .B(_09572_), .Y(_09573_));
XNOR_g _31681_ (.A(_02368_), .B(_09573_), .Y(_09574_));
NAND_g _31682_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09574_), .Y(_09575_));
NAND_g _31683_ (.A(_02367_), .B(_09394_), .Y(_09576_));
NOR_g _31684_ (.A(_02366_), .B(_09398_), .Y(_09577_));
NOR_g _31685_ (.A(_02365_), .B(_09397_), .Y(_09578_));
NOR_g _31686_ (.A(_09577_), .B(_09578_), .Y(_09579_));
AND_g _31687_ (.A(_09576_), .B(_09579_), .Y(_09580_));
NAND_g _31688_ (.A(_09575_), .B(_09580_), .Y(alu_out[14]));
NAND_g _31689_ (.A(_02368_), .B(_09571_), .Y(_09581_));
NAND_g _31690_ (.A(_02480_), .B(_09581_), .Y(_09582_));
NAND_g _31691_ (.A(instr_sub), .B(_09582_), .Y(_09583_));
NAND_g _31692_ (.A(_02367_), .B(_09569_), .Y(_09584_));
AND_g _31693_ (.A(_10910_), .B(_02366_), .Y(_09585_));
NAND_g _31694_ (.A(_09584_), .B(_09585_), .Y(_09586_));
AND_g _31695_ (.A(_09583_), .B(_09586_), .Y(_09587_));
XNOR_g _31696_ (.A(_02364_), .B(_09587_), .Y(_09588_));
NAND_g _31697_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09588_), .Y(_09589_));
NAND_g _31698_ (.A(_02363_), .B(_09394_), .Y(_09590_));
NOR_g _31699_ (.A(_02362_), .B(_09398_), .Y(_09591_));
NOR_g _31700_ (.A(_02361_), .B(_09397_), .Y(_09592_));
NOR_g _31701_ (.A(_09591_), .B(_09592_), .Y(_09593_));
AND_g _31702_ (.A(_09590_), .B(_09593_), .Y(_09594_));
NAND_g _31703_ (.A(_09589_), .B(_09594_), .Y(alu_out[15]));
AND_g _31704_ (.A(_02362_), .B(_02366_), .Y(_09595_));
AND_g _31705_ (.A(_09584_), .B(_09595_), .Y(_09596_));
NOR_g _31706_ (.A(_02361_), .B(_09596_), .Y(_09597_));
NOR_g _31707_ (.A(instr_sub), .B(_09597_), .Y(_09598_));
AND_g _31708_ (.A(instr_sub), .B(_02485_), .Y(_09599_));
NOR_g _31709_ (.A(_09598_), .B(_09599_), .Y(_09600_));
XNOR_g _31710_ (.A(_02358_), .B(_09600_), .Y(_09601_));
NAND_g _31711_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09601_), .Y(_09602_));
NAND_g _31712_ (.A(_02357_), .B(_09394_), .Y(_09603_));
NOR_g _31713_ (.A(_02356_), .B(_09398_), .Y(_09604_));
NOR_g _31714_ (.A(_02355_), .B(_09397_), .Y(_09605_));
NOR_g _31715_ (.A(_09604_), .B(_09605_), .Y(_09606_));
AND_g _31716_ (.A(_09603_), .B(_09606_), .Y(_09607_));
NAND_g _31717_ (.A(_09602_), .B(_09607_), .Y(alu_out[16]));
AND_g _31718_ (.A(_02358_), .B(_02485_), .Y(_09608_));
NAND_g _31719_ (.A(_02358_), .B(_02485_), .Y(_09609_));
NAND_g _31720_ (.A(_02345_), .B(_09609_), .Y(_09610_));
NAND_g _31721_ (.A(instr_sub), .B(_09610_), .Y(_09611_));
NAND_g _31722_ (.A(_02357_), .B(_09597_), .Y(_09612_));
AND_g _31723_ (.A(_10910_), .B(_02356_), .Y(_09613_));
NAND_g _31724_ (.A(_09612_), .B(_09613_), .Y(_09614_));
AND_g _31725_ (.A(_09611_), .B(_09614_), .Y(_09615_));
XNOR_g _31726_ (.A(_02343_), .B(_09615_), .Y(_09616_));
NAND_g _31727_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09616_), .Y(_09617_));
NAND_g _31728_ (.A(_02342_), .B(_09394_), .Y(_09618_));
NOR_g _31729_ (.A(_02339_), .B(_09397_), .Y(_09619_));
NOR_g _31730_ (.A(_02341_), .B(_09398_), .Y(_09620_));
NOR_g _31731_ (.A(_09619_), .B(_09620_), .Y(_09621_));
AND_g _31732_ (.A(_09618_), .B(_09621_), .Y(_09622_));
NAND_g _31733_ (.A(_09617_), .B(_09622_), .Y(alu_out[17]));
NAND_g _31734_ (.A(_02343_), .B(_09608_), .Y(_09623_));
NAND_g _31735_ (.A(_02347_), .B(_09623_), .Y(_09624_));
NAND_g _31736_ (.A(instr_sub), .B(_09624_), .Y(_09625_));
AND_g _31737_ (.A(_02341_), .B(_02356_), .Y(_09626_));
NAND_g _31738_ (.A(_09612_), .B(_09626_), .Y(_09627_));
AND_g _31739_ (.A(_02340_), .B(_09627_), .Y(_09628_));
NAND_g _31740_ (.A(_02340_), .B(_09627_), .Y(_09629_));
NAND_g _31741_ (.A(_10910_), .B(_09629_), .Y(_09630_));
AND_g _31742_ (.A(_09625_), .B(_09630_), .Y(_09631_));
NAND_g _31743_ (.A(_02336_), .B(_09631_), .Y(_09632_));
NOR_g _31744_ (.A(_02336_), .B(_09631_), .Y(_09633_));
NOR_g _31745_ (.A(_11210_), .B(_09633_), .Y(_09634_));
NAND_g _31746_ (.A(_09632_), .B(_09634_), .Y(_09635_));
NAND_g _31747_ (.A(_02336_), .B(_09394_), .Y(_09636_));
NOR_g _31748_ (.A(_02335_), .B(_09398_), .Y(_09637_));
NOR_g _31749_ (.A(_02334_), .B(_09397_), .Y(_09638_));
NOR_g _31750_ (.A(_09637_), .B(_09638_), .Y(_09639_));
AND_g _31751_ (.A(_09636_), .B(_09639_), .Y(_09640_));
NAND_g _31752_ (.A(_09635_), .B(_09640_), .Y(alu_out[18]));
NAND_g _31753_ (.A(_02337_), .B(_09624_), .Y(_09641_));
NAND_g _31754_ (.A(_02333_), .B(_09641_), .Y(_09642_));
NAND_g _31755_ (.A(instr_sub), .B(_09642_), .Y(_09643_));
NAND_g _31756_ (.A(_02336_), .B(_09628_), .Y(_09644_));
AND_g _31757_ (.A(_10910_), .B(_02335_), .Y(_09645_));
NAND_g _31758_ (.A(_09644_), .B(_09645_), .Y(_09646_));
AND_g _31759_ (.A(_09643_), .B(_09646_), .Y(_09647_));
XNOR_g _31760_ (.A(_02332_), .B(_09647_), .Y(_09648_));
NAND_g _31761_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09648_), .Y(_09649_));
NAND_g _31762_ (.A(_02331_), .B(_09394_), .Y(_09650_));
NOR_g _31763_ (.A(_02329_), .B(_09397_), .Y(_09651_));
NOR_g _31764_ (.A(_02330_), .B(_09398_), .Y(_09652_));
NOR_g _31765_ (.A(_09651_), .B(_09652_), .Y(_09653_));
AND_g _31766_ (.A(_09650_), .B(_09653_), .Y(_09654_));
NAND_g _31767_ (.A(_09649_), .B(_09654_), .Y(alu_out[19]));
AND_g _31768_ (.A(_02330_), .B(_02335_), .Y(_09655_));
AND_g _31769_ (.A(_09644_), .B(_09655_), .Y(_09656_));
NOR_g _31770_ (.A(_02329_), .B(_09656_), .Y(_09657_));
NOR_g _31771_ (.A(instr_sub), .B(_09657_), .Y(_09658_));
AND_g _31772_ (.A(instr_sub), .B(_02487_), .Y(_09659_));
NOR_g _31773_ (.A(_09658_), .B(_09659_), .Y(_09660_));
XNOR_g _31774_ (.A(_02325_), .B(_09660_), .Y(_09661_));
NAND_g _31775_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09661_), .Y(_09662_));
NAND_g _31776_ (.A(_02324_), .B(_09394_), .Y(_09663_));
NOR_g _31777_ (.A(_02323_), .B(_09398_), .Y(_09664_));
NOR_g _31778_ (.A(_02322_), .B(_09397_), .Y(_09665_));
NOR_g _31779_ (.A(_09664_), .B(_09665_), .Y(_09666_));
AND_g _31780_ (.A(_09663_), .B(_09666_), .Y(_09667_));
NAND_g _31781_ (.A(_09662_), .B(_09667_), .Y(alu_out[20]));
NAND_g _31782_ (.A(_02325_), .B(_02487_), .Y(_09668_));
NAND_g _31783_ (.A(_02314_), .B(_09668_), .Y(_09669_));
NAND_g _31784_ (.A(instr_sub), .B(_09669_), .Y(_09670_));
NAND_g _31785_ (.A(_02324_), .B(_09657_), .Y(_09671_));
AND_g _31786_ (.A(_10910_), .B(_02323_), .Y(_09672_));
NAND_g _31787_ (.A(_09671_), .B(_09672_), .Y(_09673_));
AND_g _31788_ (.A(_09670_), .B(_09673_), .Y(_09674_));
XNOR_g _31789_ (.A(_02312_), .B(_09674_), .Y(_09675_));
NAND_g _31790_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09675_), .Y(_09676_));
NAND_g _31791_ (.A(_02311_), .B(_09394_), .Y(_09677_));
NOR_g _31792_ (.A(_02309_), .B(_09397_), .Y(_09678_));
NOR_g _31793_ (.A(_02310_), .B(_09398_), .Y(_09679_));
NOR_g _31794_ (.A(_09678_), .B(_09679_), .Y(_09680_));
AND_g _31795_ (.A(_09677_), .B(_09680_), .Y(_09681_));
NAND_g _31796_ (.A(_09676_), .B(_09681_), .Y(alu_out[21]));
NAND_g _31797_ (.A(_02312_), .B(_09669_), .Y(_09682_));
NAND_g _31798_ (.A(_02308_), .B(_09682_), .Y(_09683_));
AND_g _31799_ (.A(_02310_), .B(_02323_), .Y(_09684_));
AND_g _31800_ (.A(_09671_), .B(_09684_), .Y(_09685_));
NOR_g _31801_ (.A(_02309_), .B(_09685_), .Y(_09686_));
NOR_g _31802_ (.A(instr_sub), .B(_09686_), .Y(_09687_));
AND_g _31803_ (.A(instr_sub), .B(_09683_), .Y(_09688_));
NOR_g _31804_ (.A(_09687_), .B(_09688_), .Y(_09689_));
XNOR_g _31805_ (.A(_02307_), .B(_09689_), .Y(_09690_));
NAND_g _31806_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09690_), .Y(_09691_));
NAND_g _31807_ (.A(_02306_), .B(_09394_), .Y(_09692_));
NOR_g _31808_ (.A(_02305_), .B(_09398_), .Y(_09693_));
NOR_g _31809_ (.A(_02304_), .B(_09397_), .Y(_09694_));
NOR_g _31810_ (.A(_09693_), .B(_09694_), .Y(_09695_));
AND_g _31811_ (.A(_09692_), .B(_09695_), .Y(_09696_));
NAND_g _31812_ (.A(_09691_), .B(_09696_), .Y(alu_out[22]));
NAND_g _31813_ (.A(_02307_), .B(_09683_), .Y(_09697_));
NAND_g _31814_ (.A(_02303_), .B(_09697_), .Y(_09698_));
NAND_g _31815_ (.A(instr_sub), .B(_09698_), .Y(_09699_));
NAND_g _31816_ (.A(_02306_), .B(_09686_), .Y(_09700_));
AND_g _31817_ (.A(_10910_), .B(_02305_), .Y(_09701_));
NAND_g _31818_ (.A(_09700_), .B(_09701_), .Y(_09702_));
AND_g _31819_ (.A(_09699_), .B(_09702_), .Y(_09703_));
XNOR_g _31820_ (.A(_02302_), .B(_09703_), .Y(_09704_));
NAND_g _31821_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09704_), .Y(_09705_));
NAND_g _31822_ (.A(_02301_), .B(_09394_), .Y(_09706_));
NOR_g _31823_ (.A(_02299_), .B(_09397_), .Y(_09707_));
NOR_g _31824_ (.A(_02300_), .B(_09398_), .Y(_09708_));
NOR_g _31825_ (.A(_09707_), .B(_09708_), .Y(_09709_));
AND_g _31826_ (.A(_09706_), .B(_09709_), .Y(_09710_));
NAND_g _31827_ (.A(_09705_), .B(_09710_), .Y(alu_out[23]));
AND_g _31828_ (.A(_02300_), .B(_02305_), .Y(_09711_));
AND_g _31829_ (.A(_09700_), .B(_09711_), .Y(_09712_));
NOR_g _31830_ (.A(_02299_), .B(_09712_), .Y(_09713_));
NOR_g _31831_ (.A(instr_sub), .B(_09713_), .Y(_09714_));
AND_g _31832_ (.A(instr_sub), .B(_02489_), .Y(_09715_));
NOR_g _31833_ (.A(_09714_), .B(_09715_), .Y(_09716_));
XNOR_g _31834_ (.A(_02297_), .B(_09716_), .Y(_09717_));
NAND_g _31835_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09717_), .Y(_09718_));
NAND_g _31836_ (.A(_02296_), .B(_09394_), .Y(_09719_));
NOR_g _31837_ (.A(_02295_), .B(_09398_), .Y(_09720_));
NOR_g _31838_ (.A(_02294_), .B(_09397_), .Y(_09721_));
NOR_g _31839_ (.A(_09720_), .B(_09721_), .Y(_09722_));
AND_g _31840_ (.A(_09719_), .B(_09722_), .Y(_09723_));
NAND_g _31841_ (.A(_09718_), .B(_09723_), .Y(alu_out[24]));
NAND_g _31842_ (.A(_02290_), .B(_02491_), .Y(_09724_));
NAND_g _31843_ (.A(instr_sub), .B(_09724_), .Y(_09725_));
NAND_g _31844_ (.A(_02296_), .B(_09713_), .Y(_09726_));
AND_g _31845_ (.A(_10910_), .B(_02295_), .Y(_09727_));
NAND_g _31846_ (.A(_09726_), .B(_09727_), .Y(_09728_));
AND_g _31847_ (.A(_09725_), .B(_09728_), .Y(_09729_));
XNOR_g _31848_ (.A(_02288_), .B(_09729_), .Y(_09730_));
NAND_g _31849_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09730_), .Y(_09731_));
NAND_g _31850_ (.A(_02287_), .B(_09394_), .Y(_09732_));
NOR_g _31851_ (.A(_02285_), .B(_09397_), .Y(_09733_));
NOR_g _31852_ (.A(_02286_), .B(_09398_), .Y(_09734_));
NOR_g _31853_ (.A(_09733_), .B(_09734_), .Y(_09735_));
AND_g _31854_ (.A(_09732_), .B(_09735_), .Y(_09736_));
NAND_g _31855_ (.A(_09731_), .B(_09736_), .Y(alu_out[25]));
AND_g _31856_ (.A(_02286_), .B(_02295_), .Y(_09737_));
AND_g _31857_ (.A(_09726_), .B(_09737_), .Y(_09738_));
NOR_g _31858_ (.A(_02285_), .B(_09738_), .Y(_09739_));
NOR_g _31859_ (.A(instr_sub), .B(_09739_), .Y(_09740_));
AND_g _31860_ (.A(instr_sub), .B(_02493_), .Y(_09741_));
NOR_g _31861_ (.A(_09740_), .B(_09741_), .Y(_09742_));
XNOR_g _31862_ (.A(_02497_), .B(_09742_), .Y(_09743_));
NAND_g _31863_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09743_), .Y(_09744_));
NAND_g _31864_ (.A(_02496_), .B(_09394_), .Y(_09745_));
NOR_g _31865_ (.A(_02495_), .B(_09398_), .Y(_09746_));
NOR_g _31866_ (.A(_02494_), .B(_09397_), .Y(_09747_));
NOR_g _31867_ (.A(_09746_), .B(_09747_), .Y(_09748_));
AND_g _31868_ (.A(_09745_), .B(_09748_), .Y(_09749_));
NAND_g _31869_ (.A(_09744_), .B(_09749_), .Y(alu_out[26]));
NAND_g _31870_ (.A(_02280_), .B(_02498_), .Y(_09750_));
NAND_g _31871_ (.A(instr_sub), .B(_09750_), .Y(_09751_));
NAND_g _31872_ (.A(_02496_), .B(_09739_), .Y(_09752_));
AND_g _31873_ (.A(_10910_), .B(_02495_), .Y(_09753_));
NAND_g _31874_ (.A(_09752_), .B(_09753_), .Y(_09754_));
AND_g _31875_ (.A(_09751_), .B(_09754_), .Y(_09755_));
XNOR_g _31876_ (.A(_02278_), .B(_09755_), .Y(_09756_));
NAND_g _31877_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09756_), .Y(_09757_));
NAND_g _31878_ (.A(_02277_), .B(_09394_), .Y(_09758_));
NOR_g _31879_ (.A(_02276_), .B(_09398_), .Y(_09759_));
NOR_g _31880_ (.A(_02274_), .B(_09397_), .Y(_09760_));
NOR_g _31881_ (.A(_09759_), .B(_09760_), .Y(_09761_));
AND_g _31882_ (.A(_09758_), .B(_09761_), .Y(_09762_));
NAND_g _31883_ (.A(_09757_), .B(_09762_), .Y(alu_out[27]));
AND_g _31884_ (.A(_02276_), .B(_02495_), .Y(_09763_));
NAND_g _31885_ (.A(_09752_), .B(_09763_), .Y(_09764_));
NAND_g _31886_ (.A(_02275_), .B(_09764_), .Y(_09765_));
NAND_g _31887_ (.A(_10910_), .B(_09765_), .Y(_09766_));
NAND_g _31888_ (.A(instr_sub), .B(_02501_), .Y(_09767_));
AND_g _31889_ (.A(_09766_), .B(_09767_), .Y(_09768_));
XNOR_g _31890_ (.A(_02273_), .B(_09768_), .Y(_09769_));
NAND_g _31891_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09769_), .Y(_09770_));
NAND_g _31892_ (.A(_02272_), .B(_09394_), .Y(_09771_));
NOR_g _31893_ (.A(_02270_), .B(_09397_), .Y(_09772_));
NOR_g _31894_ (.A(_02271_), .B(_09398_), .Y(_09773_));
NOR_g _31895_ (.A(_09772_), .B(_09773_), .Y(_09774_));
AND_g _31896_ (.A(_09771_), .B(_09774_), .Y(_09775_));
NAND_g _31897_ (.A(_09770_), .B(_09775_), .Y(alu_out[28]));
AND_g _31898_ (.A(_02271_), .B(_09765_), .Y(_09776_));
NOR_g _31899_ (.A(_02270_), .B(_09776_), .Y(_09777_));
NAND_g _31900_ (.A(_10910_), .B(_09777_), .Y(_09778_));
NOR_g _31901_ (.A(_10910_), .B(_02266_), .Y(_09779_));
NAND_g _31902_ (.A(_02503_), .B(_09779_), .Y(_09780_));
AND_g _31903_ (.A(_09778_), .B(_09780_), .Y(_09781_));
XNOR_g _31904_ (.A(_02264_), .B(_09781_), .Y(_09782_));
NAND_g _31905_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09782_), .Y(_09783_));
NAND_g _31906_ (.A(_02264_), .B(_09394_), .Y(_09784_));
NOR_g _31907_ (.A(_02263_), .B(_09398_), .Y(_09785_));
NOR_g _31908_ (.A(_02261_), .B(_09397_), .Y(_09786_));
NOR_g _31909_ (.A(_09785_), .B(_09786_), .Y(_09787_));
AND_g _31910_ (.A(_09784_), .B(_09787_), .Y(_09788_));
NAND_g _31911_ (.A(_09783_), .B(_09788_), .Y(alu_out[29]));
NOR_g _31912_ (.A(_02262_), .B(_09777_), .Y(_09789_));
NOR_g _31913_ (.A(_02261_), .B(_09789_), .Y(_09790_));
NOR_g _31914_ (.A(instr_sub), .B(_09790_), .Y(_09791_));
AND_g _31915_ (.A(instr_sub), .B(_02505_), .Y(_09792_));
NOR_g _31916_ (.A(_09791_), .B(_09792_), .Y(_09793_));
XNOR_g _31917_ (.A(_02259_), .B(_09793_), .Y(_09794_));
NAND_g _31918_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09794_), .Y(_09795_));
NAND_g _31919_ (.A(_02258_), .B(_09394_), .Y(_09796_));
NOR_g _31920_ (.A(_02257_), .B(_09398_), .Y(_09797_));
NOR_g _31921_ (.A(_02256_), .B(_09397_), .Y(_09798_));
NOR_g _31922_ (.A(_09797_), .B(_09798_), .Y(_09799_));
AND_g _31923_ (.A(_09796_), .B(_09799_), .Y(_09800_));
NAND_g _31924_ (.A(_09795_), .B(_09800_), .Y(alu_out[30]));
NAND_g _31925_ (.A(instr_sub), .B(_02508_), .Y(_09801_));
NAND_g _31926_ (.A(_02258_), .B(_09790_), .Y(_09802_));
AND_g _31927_ (.A(_10910_), .B(_02257_), .Y(_09803_));
NAND_g _31928_ (.A(_09802_), .B(_09803_), .Y(_09804_));
AND_g _31929_ (.A(_09801_), .B(_09804_), .Y(_09805_));
XNOR_g _31930_ (.A(_02254_), .B(_09805_), .Y(_09806_));
NAND_g _31931_ (.A(is_lui_auipc_jal_jalr_addi_add_sub), .B(_09806_), .Y(_09807_));
NAND_g _31932_ (.A(_02253_), .B(_09394_), .Y(_09808_));
NOR_g _31933_ (.A(_02251_), .B(_09397_), .Y(_09809_));
NOR_g _31934_ (.A(_02252_), .B(_09398_), .Y(_09810_));
NOR_g _31935_ (.A(_09809_), .B(_09810_), .Y(_09811_));
AND_g _31936_ (.A(_09808_), .B(_09811_), .Y(_09812_));
NAND_g _31937_ (.A(_09807_), .B(_09812_), .Y(alu_out[31]));
AND_g _31938_ (.A(_11272_), .B(_13410_), .Y(_09813_));
NAND_g _31939_ (.A(_13413_), .B(_09813_), .Y(dbg_ascii_state[0]));
NAND_g _31940_ (.A(_11272_), .B(_13725_), .Y(dbg_ascii_state[1]));
AND_g _31941_ (.A(_13726_), .B(_02617_), .Y(_09814_));
NOT_g _31942_ (.A(_09814_), .Y(dbg_ascii_state[17]));
NAND_g _31943_ (.A(_13388_), .B(_09814_), .Y(dbg_ascii_state[4]));
NAND_g _31944_ (.A(_11272_), .B(_13412_), .Y(dbg_ascii_state[19]));
AND_g _31945_ (.A(_02618_), .B(_09814_), .Y(_09815_));
NOT_g _31946_ (.A(_09815_), .Y(dbg_ascii_state[20]));
NAND_g _31947_ (.A(_13413_), .B(_09815_), .Y(dbg_ascii_state[26]));
NAND_g _31948_ (.A(_13394_), .B(_09814_), .Y(dbg_ascii_state[28]));
AND_g _31949_ (.A(_13412_), .B(_02617_), .Y(_09816_));
NAND_g _31950_ (.A(_02618_), .B(_09816_), .Y(dbg_ascii_state[29]));
NAND_g _31951_ (.A(_04758_), .B(_09816_), .Y(dbg_ascii_state[30]));
NAND_g _31952_ (.A(_11263_), .B(_13411_), .Y(dbg_ascii_state[33]));
NAND_g _31953_ (.A(_13726_), .B(_02768_), .Y(dbg_ascii_state[34]));
AND_g _31954_ (.A(_11271_), .B(_11918_), .Y(_09817_));
NAND_g _31955_ (.A(_02564_), .B(_09817_), .Y(_09818_));
NAND_g _31956_ (.A(_11272_), .B(_11918_), .Y(_09819_));
AND_g _31957_ (.A(_02226_), .B(_09819_), .Y(_09820_));
NAND_g _31958_ (.A(_09818_), .B(_09820_), .Y(_00004_));
NAND_g _31959_ (.A(_10894_), .B(_10895_), .Y(_09821_));
NOR_g _31960_ (.A(latched_is_lb), .B(_09821_), .Y(_09822_));
NOT_g _31961_ (.A(_09822_), .Y(_09823_));
AND_g _31962_ (.A(dbg_ascii_state[35]), .B(_02225_), .Y(_09824_));
AND_g _31963_ (.A(_09823_), .B(_09824_), .Y(_09825_));
NAND_g _31964_ (.A(mem_rdata[16]), .B(_04054_), .Y(_09826_));
NAND_g _31965_ (.A(mem_rdata[0]), .B(mem_la_wstrb[0]), .Y(_09827_));
NAND_g _31966_ (.A(mem_rdata[24]), .B(_04059_), .Y(_09828_));
AND_g _31967_ (.A(_03928_), .B(_04045_), .Y(_09829_));
NAND_g _31968_ (.A(mem_rdata[8]), .B(_09829_), .Y(_09830_));
AND_g _31969_ (.A(_09828_), .B(_09830_), .Y(_09831_));
AND_g _31970_ (.A(_09827_), .B(_09831_), .Y(_09832_));
NAND_g _31971_ (.A(_09826_), .B(_09832_), .Y(_09833_));
NAND_g _31972_ (.A(_09825_), .B(_09833_), .Y(_09834_));
NAND_g _31973_ (.A(count_instr[0]), .B(instr_rdinstr), .Y(_09835_));
NAND_g _31974_ (.A(instr_rdcycleh), .B(count_cycle[32]), .Y(_09836_));
AND_g _31975_ (.A(_09835_), .B(_09836_), .Y(_09837_));
NAND_g _31976_ (.A(count_instr[32]), .B(instr_rdinstrh), .Y(_09838_));
NAND_g _31977_ (.A(instr_rdcycle), .B(count_cycle[0]), .Y(_09839_));
AND_g _31978_ (.A(_09838_), .B(_09839_), .Y(_09840_));
NAND_g _31979_ (.A(_09837_), .B(_09840_), .Y(_09841_));
NAND_g _31980_ (.A(_13409_), .B(_09841_), .Y(_09842_));
NAND_g _31981_ (.A(pcpi_rs1[0]), .B(_13416_), .Y(_09843_));
AND_g _31982_ (.A(_09842_), .B(_09843_), .Y(_09844_));
NAND_g _31983_ (.A(_09834_), .B(_09844_), .Y(_09845_));
NAND_g _31984_ (.A(resetn), .B(_09845_), .Y(_09846_));
AND_g _31985_ (.A(reg_next_pc[0]), .B(decoded_imm[0]), .Y(_09847_));
NAND_g _31986_ (.A(reg_next_pc[0]), .B(decoded_imm[0]), .Y(_09848_));
XOR_g _31987_ (.A(reg_next_pc[0]), .B(decoded_imm[0]), .Y(_09849_));
NAND_g _31988_ (.A(_02563_), .B(_09849_), .Y(_09850_));
NAND_g _31989_ (.A(_09846_), .B(_09850_), .Y(_00009_[0]));
NAND_g _31990_ (.A(mem_rdata[17]), .B(_04054_), .Y(_09851_));
NAND_g _31991_ (.A(mem_rdata[1]), .B(mem_la_wstrb[0]), .Y(_09852_));
NAND_g _31992_ (.A(mem_rdata[9]), .B(_09829_), .Y(_09853_));
NAND_g _31993_ (.A(mem_rdata[25]), .B(_04059_), .Y(_09854_));
AND_g _31994_ (.A(_09853_), .B(_09854_), .Y(_09855_));
AND_g _31995_ (.A(_09852_), .B(_09855_), .Y(_09856_));
NAND_g _31996_ (.A(_09851_), .B(_09856_), .Y(_09857_));
NAND_g _31997_ (.A(_09825_), .B(_09857_), .Y(_09858_));
NAND_g _31998_ (.A(pcpi_rs1[1]), .B(_13416_), .Y(_09859_));
NAND_g _31999_ (.A(reg_pc[1]), .B(decoded_imm[1]), .Y(_09860_));
XOR_g _32000_ (.A(reg_pc[1]), .B(decoded_imm[1]), .Y(_09861_));
XNOR_g _32001_ (.A(reg_pc[1]), .B(decoded_imm[1]), .Y(_09862_));
NAND_g _32002_ (.A(_09848_), .B(_09862_), .Y(_09863_));
NAND_g _32003_ (.A(_09847_), .B(_09861_), .Y(_09864_));
AND_g _32004_ (.A(_11271_), .B(_09863_), .Y(_09865_));
NAND_g _32005_ (.A(_09864_), .B(_09865_), .Y(_09866_));
NAND_g _32006_ (.A(count_instr[1]), .B(instr_rdinstr), .Y(_09867_));
NAND_g _32007_ (.A(instr_rdcycleh), .B(count_cycle[33]), .Y(_09868_));
AND_g _32008_ (.A(_09867_), .B(_09868_), .Y(_09869_));
NAND_g _32009_ (.A(instr_rdcycle), .B(count_cycle[1]), .Y(_09870_));
NAND_g _32010_ (.A(count_instr[33]), .B(instr_rdinstrh), .Y(_09871_));
AND_g _32011_ (.A(_09870_), .B(_09871_), .Y(_09872_));
NAND_g _32012_ (.A(_09869_), .B(_09872_), .Y(_09873_));
NAND_g _32013_ (.A(_13409_), .B(_09873_), .Y(_09874_));
AND_g _32014_ (.A(_09866_), .B(_09874_), .Y(_09875_));
AND_g _32015_ (.A(_09859_), .B(_09875_), .Y(_09876_));
NAND_g _32016_ (.A(_09858_), .B(_09876_), .Y(_09877_));
AND_g _32017_ (.A(resetn), .B(_09877_), .Y(_00009_[1]));
NAND_g _32018_ (.A(mem_rdata[18]), .B(_04054_), .Y(_09878_));
NAND_g _32019_ (.A(mem_rdata[26]), .B(_04059_), .Y(_09879_));
NAND_g _32020_ (.A(mem_rdata[10]), .B(_09829_), .Y(_09880_));
NAND_g _32021_ (.A(mem_rdata[2]), .B(mem_la_wstrb[0]), .Y(_09881_));
AND_g _32022_ (.A(_09880_), .B(_09881_), .Y(_09882_));
AND_g _32023_ (.A(_09879_), .B(_09882_), .Y(_09883_));
NAND_g _32024_ (.A(_09878_), .B(_09883_), .Y(_09884_));
NAND_g _32025_ (.A(_09825_), .B(_09884_), .Y(_09885_));
NAND_g _32026_ (.A(pcpi_rs1[2]), .B(_13416_), .Y(_09886_));
NAND_g _32027_ (.A(instr_rdcycle), .B(count_cycle[2]), .Y(_09887_));
NAND_g _32028_ (.A(count_instr[34]), .B(instr_rdinstrh), .Y(_09888_));
NAND_g _32029_ (.A(count_instr[2]), .B(instr_rdinstr), .Y(_09889_));
NAND_g _32030_ (.A(instr_rdcycleh), .B(count_cycle[34]), .Y(_09890_));
AND_g _32031_ (.A(_09888_), .B(_09890_), .Y(_09891_));
AND_g _32032_ (.A(_09887_), .B(_09889_), .Y(_09892_));
NAND_g _32033_ (.A(_09891_), .B(_09892_), .Y(_09893_));
NAND_g _32034_ (.A(_13409_), .B(_09893_), .Y(_09894_));
AND_g _32035_ (.A(_09886_), .B(_09894_), .Y(_09895_));
NAND_g _32036_ (.A(_09885_), .B(_09895_), .Y(_09896_));
NAND_g _32037_ (.A(resetn), .B(_09896_), .Y(_09897_));
NAND_g _32038_ (.A(_09860_), .B(_09864_), .Y(_09898_));
NAND_g _32039_ (.A(reg_pc[2]), .B(decoded_imm[2]), .Y(_09899_));
XOR_g _32040_ (.A(reg_pc[2]), .B(decoded_imm[2]), .Y(_09900_));
NAND_g _32041_ (.A(_09898_), .B(_09900_), .Y(_09901_));
XOR_g _32042_ (.A(_09898_), .B(_09900_), .Y(_09902_));
NAND_g _32043_ (.A(_02563_), .B(_09902_), .Y(_09903_));
NAND_g _32044_ (.A(_09897_), .B(_09903_), .Y(_00009_[2]));
NAND_g _32045_ (.A(mem_rdata[19]), .B(_04054_), .Y(_09904_));
NAND_g _32046_ (.A(mem_rdata[27]), .B(_04059_), .Y(_09905_));
NAND_g _32047_ (.A(mem_rdata[11]), .B(_09829_), .Y(_09906_));
NAND_g _32048_ (.A(mem_rdata[3]), .B(mem_la_wstrb[0]), .Y(_09907_));
AND_g _32049_ (.A(_09906_), .B(_09907_), .Y(_09908_));
AND_g _32050_ (.A(_09905_), .B(_09908_), .Y(_09909_));
NAND_g _32051_ (.A(_09904_), .B(_09909_), .Y(_09910_));
NAND_g _32052_ (.A(_09825_), .B(_09910_), .Y(_09911_));
NAND_g _32053_ (.A(pcpi_rs1[3]), .B(_13416_), .Y(_09912_));
NAND_g _32054_ (.A(count_instr[3]), .B(instr_rdinstr), .Y(_09913_));
NAND_g _32055_ (.A(instr_rdcycleh), .B(count_cycle[35]), .Y(_09914_));
AND_g _32056_ (.A(_09913_), .B(_09914_), .Y(_09915_));
NAND_g _32057_ (.A(count_instr[35]), .B(instr_rdinstrh), .Y(_09916_));
NAND_g _32058_ (.A(instr_rdcycle), .B(count_cycle[3]), .Y(_09917_));
AND_g _32059_ (.A(_09916_), .B(_09917_), .Y(_09918_));
NAND_g _32060_ (.A(_09915_), .B(_09918_), .Y(_09919_));
NAND_g _32061_ (.A(_13409_), .B(_09919_), .Y(_09920_));
AND_g _32062_ (.A(_09912_), .B(_09920_), .Y(_09921_));
NAND_g _32063_ (.A(_09899_), .B(_09901_), .Y(_09922_));
NAND_g _32064_ (.A(reg_pc[3]), .B(decoded_imm[3]), .Y(_09923_));
XOR_g _32065_ (.A(reg_pc[3]), .B(decoded_imm[3]), .Y(_09924_));
NAND_g _32066_ (.A(_09922_), .B(_09924_), .Y(_09925_));
XOR_g _32067_ (.A(_09922_), .B(_09924_), .Y(_09926_));
NAND_g _32068_ (.A(_11271_), .B(_09926_), .Y(_09927_));
AND_g _32069_ (.A(_09921_), .B(_09927_), .Y(_09928_));
NAND_g _32070_ (.A(_09911_), .B(_09928_), .Y(_09929_));
AND_g _32071_ (.A(resetn), .B(_09929_), .Y(_00009_[3]));
NAND_g _32072_ (.A(mem_rdata[20]), .B(_04054_), .Y(_09930_));
NAND_g _32073_ (.A(mem_rdata[28]), .B(_04059_), .Y(_09931_));
NAND_g _32074_ (.A(mem_rdata[4]), .B(mem_la_wstrb[0]), .Y(_09932_));
NAND_g _32075_ (.A(mem_rdata[12]), .B(_09829_), .Y(_09933_));
AND_g _32076_ (.A(_09932_), .B(_09933_), .Y(_09934_));
AND_g _32077_ (.A(_09931_), .B(_09934_), .Y(_09935_));
NAND_g _32078_ (.A(_09930_), .B(_09935_), .Y(_09936_));
NAND_g _32079_ (.A(_09825_), .B(_09936_), .Y(_09937_));
NAND_g _32080_ (.A(pcpi_rs1[4]), .B(_13416_), .Y(_09938_));
NAND_g _32081_ (.A(count_instr[4]), .B(instr_rdinstr), .Y(_09939_));
NAND_g _32082_ (.A(instr_rdcycleh), .B(count_cycle[36]), .Y(_09940_));
AND_g _32083_ (.A(_09939_), .B(_09940_), .Y(_09941_));
NAND_g _32084_ (.A(count_instr[36]), .B(instr_rdinstrh), .Y(_09942_));
NAND_g _32085_ (.A(instr_rdcycle), .B(count_cycle[4]), .Y(_09943_));
AND_g _32086_ (.A(_09942_), .B(_09943_), .Y(_09944_));
NAND_g _32087_ (.A(_09941_), .B(_09944_), .Y(_09945_));
NAND_g _32088_ (.A(_13409_), .B(_09945_), .Y(_09946_));
AND_g _32089_ (.A(_09938_), .B(_09946_), .Y(_09947_));
NAND_g _32090_ (.A(_09937_), .B(_09947_), .Y(_09948_));
NAND_g _32091_ (.A(_09923_), .B(_09925_), .Y(_09949_));
NAND_g _32092_ (.A(reg_pc[4]), .B(decoded_imm[4]), .Y(_09950_));
XOR_g _32093_ (.A(reg_pc[4]), .B(decoded_imm[4]), .Y(_09951_));
NAND_g _32094_ (.A(_09949_), .B(_09951_), .Y(_09952_));
XOR_g _32095_ (.A(_09949_), .B(_09951_), .Y(_09953_));
NAND_g _32096_ (.A(_02563_), .B(_09953_), .Y(_09954_));
NAND_g _32097_ (.A(resetn), .B(_09948_), .Y(_09955_));
NAND_g _32098_ (.A(_09954_), .B(_09955_), .Y(_00009_[4]));
NAND_g _32099_ (.A(mem_rdata[21]), .B(_04054_), .Y(_09956_));
NAND_g _32100_ (.A(mem_rdata[29]), .B(_04059_), .Y(_09957_));
NAND_g _32101_ (.A(mem_rdata[5]), .B(mem_la_wstrb[0]), .Y(_09958_));
NAND_g _32102_ (.A(mem_rdata[13]), .B(_09829_), .Y(_09959_));
AND_g _32103_ (.A(_09958_), .B(_09959_), .Y(_09960_));
AND_g _32104_ (.A(_09957_), .B(_09960_), .Y(_09961_));
NAND_g _32105_ (.A(_09956_), .B(_09961_), .Y(_09962_));
NAND_g _32106_ (.A(_09825_), .B(_09962_), .Y(_09963_));
NAND_g _32107_ (.A(pcpi_rs1[5]), .B(_13416_), .Y(_09964_));
NAND_g _32108_ (.A(count_instr[37]), .B(instr_rdinstrh), .Y(_09965_));
NAND_g _32109_ (.A(count_instr[5]), .B(instr_rdinstr), .Y(_09966_));
AND_g _32110_ (.A(_09965_), .B(_09966_), .Y(_09967_));
NAND_g _32111_ (.A(instr_rdcycle), .B(count_cycle[5]), .Y(_09968_));
NAND_g _32112_ (.A(instr_rdcycleh), .B(count_cycle[37]), .Y(_09969_));
AND_g _32113_ (.A(_09968_), .B(_09969_), .Y(_09970_));
NAND_g _32114_ (.A(_09967_), .B(_09970_), .Y(_09971_));
NAND_g _32115_ (.A(_13409_), .B(_09971_), .Y(_09972_));
AND_g _32116_ (.A(_09964_), .B(_09972_), .Y(_09973_));
NAND_g _32117_ (.A(_09963_), .B(_09973_), .Y(_09974_));
NAND_g _32118_ (.A(_09950_), .B(_09952_), .Y(_09975_));
NAND_g _32119_ (.A(reg_pc[5]), .B(decoded_imm[5]), .Y(_09976_));
XOR_g _32120_ (.A(reg_pc[5]), .B(decoded_imm[5]), .Y(_09977_));
NAND_g _32121_ (.A(_09975_), .B(_09977_), .Y(_09978_));
NAND_g _32122_ (.A(resetn), .B(_09974_), .Y(_09979_));
XOR_g _32123_ (.A(_09975_), .B(_09977_), .Y(_09980_));
NAND_g _32124_ (.A(_02563_), .B(_09980_), .Y(_09981_));
NAND_g _32125_ (.A(_09979_), .B(_09981_), .Y(_00009_[5]));
NAND_g _32126_ (.A(mem_rdata[22]), .B(_04054_), .Y(_09982_));
NAND_g _32127_ (.A(mem_rdata[6]), .B(mem_la_wstrb[0]), .Y(_09983_));
NAND_g _32128_ (.A(mem_rdata[14]), .B(_09829_), .Y(_09984_));
NAND_g _32129_ (.A(mem_rdata[30]), .B(_04059_), .Y(_09985_));
AND_g _32130_ (.A(_09984_), .B(_09985_), .Y(_09986_));
AND_g _32131_ (.A(_09983_), .B(_09986_), .Y(_09987_));
NAND_g _32132_ (.A(_09982_), .B(_09987_), .Y(_09988_));
NAND_g _32133_ (.A(_09825_), .B(_09988_), .Y(_09989_));
NAND_g _32134_ (.A(pcpi_rs1[6]), .B(_13416_), .Y(_09990_));
NAND_g _32135_ (.A(count_instr[6]), .B(instr_rdinstr), .Y(_09991_));
NAND_g _32136_ (.A(instr_rdcycleh), .B(count_cycle[38]), .Y(_09992_));
AND_g _32137_ (.A(_09991_), .B(_09992_), .Y(_09993_));
NAND_g _32138_ (.A(instr_rdcycle), .B(count_cycle[6]), .Y(_09994_));
NAND_g _32139_ (.A(count_instr[38]), .B(instr_rdinstrh), .Y(_09995_));
AND_g _32140_ (.A(_09994_), .B(_09995_), .Y(_09996_));
NAND_g _32141_ (.A(_09993_), .B(_09996_), .Y(_09997_));
NAND_g _32142_ (.A(_13409_), .B(_09997_), .Y(_09998_));
AND_g _32143_ (.A(_09990_), .B(_09998_), .Y(_09999_));
NAND_g _32144_ (.A(_09989_), .B(_09999_), .Y(_10000_));
NAND_g _32145_ (.A(resetn), .B(_10000_), .Y(_10001_));
AND_g _32146_ (.A(_09976_), .B(_09978_), .Y(_10002_));
NAND_g _32147_ (.A(_09976_), .B(_09978_), .Y(_10003_));
NAND_g _32148_ (.A(reg_pc[6]), .B(decoded_imm[6]), .Y(_10004_));
XOR_g _32149_ (.A(reg_pc[6]), .B(decoded_imm[6]), .Y(_10005_));
XNOR_g _32150_ (.A(reg_pc[6]), .B(decoded_imm[6]), .Y(_10006_));
NAND_g _32151_ (.A(_10002_), .B(_10006_), .Y(_10007_));
NAND_g _32152_ (.A(_10003_), .B(_10005_), .Y(_10008_));
AND_g _32153_ (.A(_02563_), .B(_10008_), .Y(_10009_));
NAND_g _32154_ (.A(_10007_), .B(_10009_), .Y(_10010_));
NAND_g _32155_ (.A(_10001_), .B(_10010_), .Y(_00009_[6]));
NAND_g _32156_ (.A(mem_rdata[23]), .B(_04054_), .Y(_10011_));
NAND_g _32157_ (.A(mem_rdata[31]), .B(_04059_), .Y(_10012_));
NAND_g _32158_ (.A(mem_rdata[15]), .B(_09829_), .Y(_10013_));
NAND_g _32159_ (.A(mem_rdata[7]), .B(mem_la_wstrb[0]), .Y(_10014_));
AND_g _32160_ (.A(_10013_), .B(_10014_), .Y(_10015_));
AND_g _32161_ (.A(_10012_), .B(_10015_), .Y(_10016_));
NAND_g _32162_ (.A(_10011_), .B(_10016_), .Y(_10017_));
NAND_g _32163_ (.A(_09825_), .B(_10017_), .Y(_10018_));
NAND_g _32164_ (.A(pcpi_rs1[7]), .B(_13416_), .Y(_10019_));
NAND_g _32165_ (.A(count_instr[7]), .B(instr_rdinstr), .Y(_10020_));
NAND_g _32166_ (.A(instr_rdcycleh), .B(count_cycle[39]), .Y(_10021_));
AND_g _32167_ (.A(_10020_), .B(_10021_), .Y(_10022_));
NAND_g _32168_ (.A(instr_rdcycle), .B(count_cycle[7]), .Y(_10023_));
NAND_g _32169_ (.A(count_instr[39]), .B(instr_rdinstrh), .Y(_10024_));
AND_g _32170_ (.A(_10023_), .B(_10024_), .Y(_10025_));
NAND_g _32171_ (.A(_10022_), .B(_10025_), .Y(_10026_));
NAND_g _32172_ (.A(_13409_), .B(_10026_), .Y(_10027_));
AND_g _32173_ (.A(_10019_), .B(_10027_), .Y(_10028_));
AND_g _32174_ (.A(_10004_), .B(_10008_), .Y(_10029_));
NAND_g _32175_ (.A(reg_pc[7]), .B(decoded_imm[7]), .Y(_10030_));
NOR_g _32176_ (.A(reg_pc[7]), .B(decoded_imm[7]), .Y(_10031_));
XNOR_g _32177_ (.A(reg_pc[7]), .B(decoded_imm[7]), .Y(_10032_));
NOR_g _32178_ (.A(_10029_), .B(_10032_), .Y(_10033_));
NAND_g _32179_ (.A(_10029_), .B(_10032_), .Y(_10034_));
NOR_g _32180_ (.A(_11272_), .B(_10033_), .Y(_10035_));
NAND_g _32181_ (.A(_10034_), .B(_10035_), .Y(_10036_));
AND_g _32182_ (.A(_10028_), .B(_10036_), .Y(_10037_));
NAND_g _32183_ (.A(_10018_), .B(_10037_), .Y(_10038_));
AND_g _32184_ (.A(resetn), .B(_10038_), .Y(_00009_[7]));
NAND_g _32185_ (.A(reg_pc[8]), .B(decoded_imm[8]), .Y(_10039_));
XOR_g _32186_ (.A(reg_pc[8]), .B(decoded_imm[8]), .Y(_10040_));
AND_g _32187_ (.A(_10029_), .B(_10030_), .Y(_10041_));
NOR_g _32188_ (.A(_10031_), .B(_10041_), .Y(_10042_));
NAND_g _32189_ (.A(_10040_), .B(_10042_), .Y(_10043_));
NOR_g _32190_ (.A(_10040_), .B(_10042_), .Y(_10044_));
NOR_g _32191_ (.A(_11272_), .B(_10044_), .Y(_10045_));
NAND_g _32192_ (.A(_10043_), .B(_10045_), .Y(_10046_));
NAND_g _32193_ (.A(latched_is_lb), .B(_10017_), .Y(_10047_));
NAND_g _32194_ (.A(mem_rdata[24]), .B(_04052_), .Y(_10048_));
NAND_g _32195_ (.A(mem_rdata[8]), .B(_04039_), .Y(_10049_));
NAND_g _32196_ (.A(_10048_), .B(_10049_), .Y(_10050_));
NAND_g _32197_ (.A(_09821_), .B(_10050_), .Y(_10051_));
NAND_g _32198_ (.A(_10047_), .B(_10051_), .Y(_10052_));
NAND_g _32199_ (.A(_09824_), .B(_10052_), .Y(_10053_));
NAND_g _32200_ (.A(pcpi_rs1[8]), .B(_13416_), .Y(_10054_));
NAND_g _32201_ (.A(count_instr[8]), .B(instr_rdinstr), .Y(_10055_));
NAND_g _32202_ (.A(instr_rdcycleh), .B(count_cycle[40]), .Y(_10056_));
AND_g _32203_ (.A(_10055_), .B(_10056_), .Y(_10057_));
NAND_g _32204_ (.A(instr_rdcycle), .B(count_cycle[8]), .Y(_10058_));
NAND_g _32205_ (.A(count_instr[40]), .B(instr_rdinstrh), .Y(_10059_));
AND_g _32206_ (.A(_10058_), .B(_10059_), .Y(_10060_));
NAND_g _32207_ (.A(_10057_), .B(_10060_), .Y(_10061_));
NAND_g _32208_ (.A(_13409_), .B(_10061_), .Y(_10062_));
AND_g _32209_ (.A(_10054_), .B(_10062_), .Y(_10063_));
AND_g _32210_ (.A(_10053_), .B(_10063_), .Y(_10064_));
NAND_g _32211_ (.A(_10046_), .B(_10064_), .Y(_10065_));
AND_g _32212_ (.A(resetn), .B(_10065_), .Y(_00009_[8]));
NAND_g _32213_ (.A(mem_rdata[25]), .B(_04052_), .Y(_10066_));
NAND_g _32214_ (.A(mem_rdata[9]), .B(_04039_), .Y(_10067_));
NAND_g _32215_ (.A(_10066_), .B(_10067_), .Y(_10068_));
NAND_g _32216_ (.A(_09821_), .B(_10068_), .Y(_10069_));
NAND_g _32217_ (.A(_10047_), .B(_10069_), .Y(_10070_));
NAND_g _32218_ (.A(_09824_), .B(_10070_), .Y(_10071_));
NAND_g _32219_ (.A(pcpi_rs1[9]), .B(_13416_), .Y(_10072_));
NAND_g _32220_ (.A(count_instr[9]), .B(instr_rdinstr), .Y(_10073_));
NAND_g _32221_ (.A(instr_rdcycleh), .B(count_cycle[41]), .Y(_10074_));
AND_g _32222_ (.A(_10073_), .B(_10074_), .Y(_10075_));
NAND_g _32223_ (.A(count_instr[41]), .B(instr_rdinstrh), .Y(_10076_));
NAND_g _32224_ (.A(instr_rdcycle), .B(count_cycle[9]), .Y(_10077_));
AND_g _32225_ (.A(_10076_), .B(_10077_), .Y(_10078_));
NAND_g _32226_ (.A(_10075_), .B(_10078_), .Y(_10079_));
NAND_g _32227_ (.A(_13409_), .B(_10079_), .Y(_10080_));
AND_g _32228_ (.A(_10072_), .B(_10080_), .Y(_10081_));
AND_g _32229_ (.A(_10071_), .B(_10081_), .Y(_10082_));
AND_g _32230_ (.A(_10039_), .B(_10043_), .Y(_10083_));
NAND_g _32231_ (.A(reg_pc[9]), .B(decoded_imm[9]), .Y(_10084_));
NOR_g _32232_ (.A(reg_pc[9]), .B(decoded_imm[9]), .Y(_10085_));
XOR_g _32233_ (.A(reg_pc[9]), .B(decoded_imm[9]), .Y(_10086_));
XNOR_g _32234_ (.A(_10083_), .B(_10086_), .Y(_10087_));
NAND_g _32235_ (.A(_11271_), .B(_10087_), .Y(_10088_));
NAND_g _32236_ (.A(_10082_), .B(_10088_), .Y(_10089_));
AND_g _32237_ (.A(resetn), .B(_10089_), .Y(_00009_[9]));
NAND_g _32238_ (.A(mem_rdata[26]), .B(_04052_), .Y(_10090_));
NAND_g _32239_ (.A(mem_rdata[10]), .B(_04039_), .Y(_10091_));
NAND_g _32240_ (.A(_10090_), .B(_10091_), .Y(_10092_));
NAND_g _32241_ (.A(_09821_), .B(_10092_), .Y(_10093_));
NAND_g _32242_ (.A(_10047_), .B(_10093_), .Y(_10094_));
NAND_g _32243_ (.A(_09824_), .B(_10094_), .Y(_10095_));
NAND_g _32244_ (.A(pcpi_rs1[10]), .B(_13416_), .Y(_10096_));
NAND_g _32245_ (.A(count_instr[10]), .B(instr_rdinstr), .Y(_10097_));
NAND_g _32246_ (.A(instr_rdcycleh), .B(count_cycle[42]), .Y(_10098_));
AND_g _32247_ (.A(_10097_), .B(_10098_), .Y(_10099_));
NAND_g _32248_ (.A(count_instr[42]), .B(instr_rdinstrh), .Y(_10100_));
NAND_g _32249_ (.A(instr_rdcycle), .B(count_cycle[10]), .Y(_10101_));
AND_g _32250_ (.A(_10100_), .B(_10101_), .Y(_10102_));
NAND_g _32251_ (.A(_10099_), .B(_10102_), .Y(_10103_));
NAND_g _32252_ (.A(_13409_), .B(_10103_), .Y(_10104_));
NAND_g _32253_ (.A(_10096_), .B(_10104_), .Y(_10105_));
NAND_g _32254_ (.A(reg_pc[10]), .B(decoded_imm[10]), .Y(_10106_));
XOR_g _32255_ (.A(reg_pc[10]), .B(decoded_imm[10]), .Y(_10107_));
AND_g _32256_ (.A(_10083_), .B(_10084_), .Y(_10108_));
NOR_g _32257_ (.A(_10085_), .B(_10108_), .Y(_10109_));
NOR_g _32258_ (.A(_10107_), .B(_10109_), .Y(_10110_));
NAND_g _32259_ (.A(_10107_), .B(_10109_), .Y(_10111_));
NAND_g _32260_ (.A(_11271_), .B(_10111_), .Y(_10112_));
NOR_g _32261_ (.A(_10110_), .B(_10112_), .Y(_10113_));
NOR_g _32262_ (.A(_10105_), .B(_10113_), .Y(_10114_));
NAND_g _32263_ (.A(_10095_), .B(_10114_), .Y(_10115_));
AND_g _32264_ (.A(resetn), .B(_10115_), .Y(_00009_[10]));
NAND_g _32265_ (.A(mem_rdata[27]), .B(_04052_), .Y(_10116_));
NAND_g _32266_ (.A(mem_rdata[11]), .B(_04039_), .Y(_10117_));
NAND_g _32267_ (.A(_10116_), .B(_10117_), .Y(_10118_));
NAND_g _32268_ (.A(_09821_), .B(_10118_), .Y(_10119_));
NAND_g _32269_ (.A(_10047_), .B(_10119_), .Y(_10120_));
NAND_g _32270_ (.A(_09824_), .B(_10120_), .Y(_10121_));
NAND_g _32271_ (.A(pcpi_rs1[11]), .B(_13416_), .Y(_10122_));
NAND_g _32272_ (.A(count_instr[11]), .B(instr_rdinstr), .Y(_10123_));
NAND_g _32273_ (.A(instr_rdcycleh), .B(count_cycle[43]), .Y(_10124_));
AND_g _32274_ (.A(_10123_), .B(_10124_), .Y(_10125_));
NAND_g _32275_ (.A(count_instr[43]), .B(instr_rdinstrh), .Y(_10126_));
NAND_g _32276_ (.A(instr_rdcycle), .B(count_cycle[11]), .Y(_10127_));
AND_g _32277_ (.A(_10126_), .B(_10127_), .Y(_10128_));
NAND_g _32278_ (.A(_10125_), .B(_10128_), .Y(_10129_));
NAND_g _32279_ (.A(_13409_), .B(_10129_), .Y(_10130_));
AND_g _32280_ (.A(_10122_), .B(_10130_), .Y(_10131_));
AND_g _32281_ (.A(_10121_), .B(_10131_), .Y(_10132_));
AND_g _32282_ (.A(_10106_), .B(_10111_), .Y(_10133_));
NAND_g _32283_ (.A(reg_pc[11]), .B(decoded_imm[11]), .Y(_10134_));
NOR_g _32284_ (.A(reg_pc[11]), .B(decoded_imm[11]), .Y(_10135_));
XOR_g _32285_ (.A(reg_pc[11]), .B(decoded_imm[11]), .Y(_10136_));
XNOR_g _32286_ (.A(_10133_), .B(_10136_), .Y(_10137_));
NAND_g _32287_ (.A(_11271_), .B(_10137_), .Y(_10138_));
NAND_g _32288_ (.A(_10132_), .B(_10138_), .Y(_10139_));
AND_g _32289_ (.A(resetn), .B(_10139_), .Y(_00009_[11]));
NAND_g _32290_ (.A(reg_pc[12]), .B(decoded_imm[12]), .Y(_10140_));
XOR_g _32291_ (.A(reg_pc[12]), .B(decoded_imm[12]), .Y(_10141_));
AND_g _32292_ (.A(_10133_), .B(_10134_), .Y(_10142_));
NOR_g _32293_ (.A(_10135_), .B(_10142_), .Y(_10143_));
NAND_g _32294_ (.A(_10141_), .B(_10143_), .Y(_10144_));
XOR_g _32295_ (.A(_10141_), .B(_10143_), .Y(_10145_));
NAND_g _32296_ (.A(_02563_), .B(_10145_), .Y(_10146_));
NAND_g _32297_ (.A(mem_rdata[28]), .B(_04052_), .Y(_10147_));
NAND_g _32298_ (.A(mem_rdata[12]), .B(_04039_), .Y(_10148_));
NAND_g _32299_ (.A(_10147_), .B(_10148_), .Y(_10149_));
NAND_g _32300_ (.A(_09821_), .B(_10149_), .Y(_10150_));
NAND_g _32301_ (.A(_10047_), .B(_10150_), .Y(_10151_));
NAND_g _32302_ (.A(_09824_), .B(_10151_), .Y(_10152_));
NAND_g _32303_ (.A(pcpi_rs1[12]), .B(_13416_), .Y(_10153_));
NAND_g _32304_ (.A(count_instr[12]), .B(instr_rdinstr), .Y(_10154_));
NAND_g _32305_ (.A(instr_rdcycleh), .B(count_cycle[44]), .Y(_10155_));
AND_g _32306_ (.A(_10154_), .B(_10155_), .Y(_10156_));
NAND_g _32307_ (.A(count_instr[44]), .B(instr_rdinstrh), .Y(_10157_));
NAND_g _32308_ (.A(instr_rdcycle), .B(count_cycle[12]), .Y(_10158_));
AND_g _32309_ (.A(_10157_), .B(_10158_), .Y(_10159_));
NAND_g _32310_ (.A(_10156_), .B(_10159_), .Y(_10160_));
NAND_g _32311_ (.A(_13409_), .B(_10160_), .Y(_10161_));
AND_g _32312_ (.A(_10152_), .B(_10161_), .Y(_10162_));
NAND_g _32313_ (.A(_10153_), .B(_10162_), .Y(_10163_));
NAND_g _32314_ (.A(resetn), .B(_10163_), .Y(_10164_));
NAND_g _32315_ (.A(_10146_), .B(_10164_), .Y(_00009_[12]));
AND_g _32316_ (.A(_10140_), .B(_10144_), .Y(_10165_));
NAND_g _32317_ (.A(reg_pc[13]), .B(decoded_imm[13]), .Y(_10166_));
NOR_g _32318_ (.A(reg_pc[13]), .B(decoded_imm[13]), .Y(_10167_));
XOR_g _32319_ (.A(reg_pc[13]), .B(decoded_imm[13]), .Y(_10168_));
XNOR_g _32320_ (.A(_10165_), .B(_10168_), .Y(_10169_));
NAND_g _32321_ (.A(_02563_), .B(_10169_), .Y(_10170_));
NAND_g _32322_ (.A(mem_rdata[29]), .B(_04052_), .Y(_10171_));
NAND_g _32323_ (.A(mem_rdata[13]), .B(_04039_), .Y(_10172_));
NAND_g _32324_ (.A(_10171_), .B(_10172_), .Y(_10173_));
NAND_g _32325_ (.A(_09821_), .B(_10173_), .Y(_10174_));
NAND_g _32326_ (.A(_10047_), .B(_10174_), .Y(_10175_));
NAND_g _32327_ (.A(_09824_), .B(_10175_), .Y(_10176_));
NAND_g _32328_ (.A(pcpi_rs1[13]), .B(_13416_), .Y(_10177_));
NAND_g _32329_ (.A(count_instr[13]), .B(instr_rdinstr), .Y(_10178_));
NAND_g _32330_ (.A(instr_rdcycleh), .B(count_cycle[45]), .Y(_10179_));
AND_g _32331_ (.A(_10178_), .B(_10179_), .Y(_10180_));
NAND_g _32332_ (.A(count_instr[45]), .B(instr_rdinstrh), .Y(_10181_));
NAND_g _32333_ (.A(instr_rdcycle), .B(count_cycle[13]), .Y(_10182_));
AND_g _32334_ (.A(_10181_), .B(_10182_), .Y(_10183_));
NAND_g _32335_ (.A(_10180_), .B(_10183_), .Y(_10184_));
NAND_g _32336_ (.A(_13409_), .B(_10184_), .Y(_10185_));
AND_g _32337_ (.A(_10176_), .B(_10185_), .Y(_10186_));
NAND_g _32338_ (.A(_10177_), .B(_10186_), .Y(_10187_));
NAND_g _32339_ (.A(resetn), .B(_10187_), .Y(_10188_));
NAND_g _32340_ (.A(_10170_), .B(_10188_), .Y(_00009_[13]));
NAND_g _32341_ (.A(reg_pc[14]), .B(decoded_imm[14]), .Y(_10189_));
XOR_g _32342_ (.A(reg_pc[14]), .B(decoded_imm[14]), .Y(_10190_));
AND_g _32343_ (.A(_10165_), .B(_10166_), .Y(_10191_));
NOR_g _32344_ (.A(_10167_), .B(_10191_), .Y(_10192_));
NAND_g _32345_ (.A(_10190_), .B(_10192_), .Y(_10193_));
XOR_g _32346_ (.A(_10190_), .B(_10192_), .Y(_10194_));
NAND_g _32347_ (.A(_02563_), .B(_10194_), .Y(_10195_));
NAND_g _32348_ (.A(mem_rdata[30]), .B(_04052_), .Y(_10196_));
NAND_g _32349_ (.A(mem_rdata[14]), .B(_04039_), .Y(_10197_));
NAND_g _32350_ (.A(_10196_), .B(_10197_), .Y(_10198_));
NAND_g _32351_ (.A(_09821_), .B(_10198_), .Y(_10199_));
NAND_g _32352_ (.A(_10047_), .B(_10199_), .Y(_10200_));
NAND_g _32353_ (.A(_09824_), .B(_10200_), .Y(_10201_));
NAND_g _32354_ (.A(pcpi_rs1[14]), .B(_13416_), .Y(_10202_));
NAND_g _32355_ (.A(count_instr[14]), .B(instr_rdinstr), .Y(_10203_));
NAND_g _32356_ (.A(instr_rdcycleh), .B(count_cycle[46]), .Y(_10204_));
AND_g _32357_ (.A(_10203_), .B(_10204_), .Y(_10205_));
NAND_g _32358_ (.A(count_instr[46]), .B(instr_rdinstrh), .Y(_10206_));
NAND_g _32359_ (.A(instr_rdcycle), .B(count_cycle[14]), .Y(_10207_));
AND_g _32360_ (.A(_10206_), .B(_10207_), .Y(_10208_));
NAND_g _32361_ (.A(_10205_), .B(_10208_), .Y(_10209_));
NAND_g _32362_ (.A(_13409_), .B(_10209_), .Y(_10210_));
AND_g _32363_ (.A(_10201_), .B(_10210_), .Y(_10211_));
NAND_g _32364_ (.A(_10202_), .B(_10211_), .Y(_10212_));
NAND_g _32365_ (.A(resetn), .B(_10212_), .Y(_10213_));
NAND_g _32366_ (.A(_10195_), .B(_10213_), .Y(_00009_[14]));
AND_g _32367_ (.A(_10189_), .B(_10193_), .Y(_10214_));
NAND_g _32368_ (.A(reg_pc[15]), .B(decoded_imm[15]), .Y(_10215_));
NOR_g _32369_ (.A(reg_pc[15]), .B(decoded_imm[15]), .Y(_10216_));
XOR_g _32370_ (.A(reg_pc[15]), .B(decoded_imm[15]), .Y(_10217_));
XNOR_g _32371_ (.A(_10214_), .B(_10217_), .Y(_10218_));
NAND_g _32372_ (.A(_02563_), .B(_10218_), .Y(_10219_));
NAND_g _32373_ (.A(mem_rdata[31]), .B(_04052_), .Y(_10220_));
NAND_g _32374_ (.A(mem_rdata[15]), .B(_04039_), .Y(_10221_));
NAND_g _32375_ (.A(_10220_), .B(_10221_), .Y(_10222_));
NAND_g _32376_ (.A(_09821_), .B(_10222_), .Y(_10223_));
NAND_g _32377_ (.A(_10047_), .B(_10223_), .Y(_10224_));
NAND_g _32378_ (.A(_09824_), .B(_10224_), .Y(_10225_));
NAND_g _32379_ (.A(pcpi_rs1[15]), .B(_13416_), .Y(_10226_));
NAND_g _32380_ (.A(count_instr[15]), .B(instr_rdinstr), .Y(_10227_));
NAND_g _32381_ (.A(instr_rdcycleh), .B(count_cycle[47]), .Y(_10228_));
AND_g _32382_ (.A(_10227_), .B(_10228_), .Y(_10229_));
NAND_g _32383_ (.A(instr_rdcycle), .B(count_cycle[15]), .Y(_10230_));
NAND_g _32384_ (.A(count_instr[47]), .B(instr_rdinstrh), .Y(_10231_));
AND_g _32385_ (.A(_10230_), .B(_10231_), .Y(_10232_));
NAND_g _32386_ (.A(_10229_), .B(_10232_), .Y(_10233_));
NAND_g _32387_ (.A(_13409_), .B(_10233_), .Y(_10234_));
AND_g _32388_ (.A(_10225_), .B(_10234_), .Y(_10235_));
NAND_g _32389_ (.A(_10226_), .B(_10235_), .Y(_10236_));
NAND_g _32390_ (.A(resetn), .B(_10236_), .Y(_10237_));
NAND_g _32391_ (.A(_10219_), .B(_10237_), .Y(_00009_[15]));
NAND_g _32392_ (.A(reg_pc[16]), .B(decoded_imm[16]), .Y(_10238_));
XOR_g _32393_ (.A(reg_pc[16]), .B(decoded_imm[16]), .Y(_10239_));
AND_g _32394_ (.A(_10214_), .B(_10215_), .Y(_10240_));
NOR_g _32395_ (.A(_10216_), .B(_10240_), .Y(_10241_));
NAND_g _32396_ (.A(_10239_), .B(_10241_), .Y(_10242_));
XOR_g _32397_ (.A(_10239_), .B(_10241_), .Y(_10243_));
NAND_g _32398_ (.A(_02563_), .B(_10243_), .Y(_10244_));
NAND_g _32399_ (.A(latched_is_lh), .B(_10222_), .Y(_10245_));
AND_g _32400_ (.A(_10047_), .B(_10245_), .Y(_10246_));
AND_g _32401_ (.A(latched_is_lu), .B(mem_rdata[16]), .Y(_10247_));
NAND_g _32402_ (.A(_03961_), .B(_10247_), .Y(_10248_));
NAND_g _32403_ (.A(_10246_), .B(_10248_), .Y(_10249_));
NAND_g _32404_ (.A(_09824_), .B(_10249_), .Y(_10250_));
NAND_g _32405_ (.A(pcpi_rs1[16]), .B(_13416_), .Y(_10251_));
NAND_g _32406_ (.A(count_instr[16]), .B(instr_rdinstr), .Y(_10252_));
NAND_g _32407_ (.A(instr_rdcycleh), .B(count_cycle[48]), .Y(_10253_));
AND_g _32408_ (.A(_10252_), .B(_10253_), .Y(_10254_));
NAND_g _32409_ (.A(instr_rdcycle), .B(count_cycle[16]), .Y(_10255_));
NAND_g _32410_ (.A(count_instr[48]), .B(instr_rdinstrh), .Y(_10256_));
AND_g _32411_ (.A(_10255_), .B(_10256_), .Y(_10257_));
NAND_g _32412_ (.A(_10254_), .B(_10257_), .Y(_10258_));
NAND_g _32413_ (.A(_13409_), .B(_10258_), .Y(_10259_));
AND_g _32414_ (.A(_10250_), .B(_10259_), .Y(_10260_));
NAND_g _32415_ (.A(_10251_), .B(_10260_), .Y(_10261_));
NAND_g _32416_ (.A(resetn), .B(_10261_), .Y(_10262_));
NAND_g _32417_ (.A(_10244_), .B(_10262_), .Y(_00009_[16]));
AND_g _32418_ (.A(_10238_), .B(_10242_), .Y(_10263_));
NAND_g _32419_ (.A(reg_pc[17]), .B(decoded_imm[17]), .Y(_10264_));
NOR_g _32420_ (.A(reg_pc[17]), .B(decoded_imm[17]), .Y(_10265_));
XNOR_g _32421_ (.A(reg_pc[17]), .B(decoded_imm[17]), .Y(_10266_));
NOR_g _32422_ (.A(_10263_), .B(_10266_), .Y(_10267_));
NAND_g _32423_ (.A(_10263_), .B(_10266_), .Y(_10268_));
NAND_g _32424_ (.A(_11271_), .B(_10268_), .Y(_10269_));
NOR_g _32425_ (.A(_10267_), .B(_10269_), .Y(_10270_));
AND_g _32426_ (.A(latched_is_lu), .B(mem_rdata[17]), .Y(_10271_));
NAND_g _32427_ (.A(_03961_), .B(_10271_), .Y(_10272_));
NAND_g _32428_ (.A(_10246_), .B(_10272_), .Y(_10273_));
NAND_g _32429_ (.A(_09824_), .B(_10273_), .Y(_10274_));
NAND_g _32430_ (.A(count_instr[17]), .B(instr_rdinstr), .Y(_10275_));
NAND_g _32431_ (.A(instr_rdcycleh), .B(count_cycle[49]), .Y(_10276_));
AND_g _32432_ (.A(_10275_), .B(_10276_), .Y(_10277_));
NAND_g _32433_ (.A(instr_rdcycle), .B(count_cycle[17]), .Y(_10278_));
NAND_g _32434_ (.A(count_instr[49]), .B(instr_rdinstrh), .Y(_10279_));
AND_g _32435_ (.A(_10278_), .B(_10279_), .Y(_10280_));
NAND_g _32436_ (.A(_10277_), .B(_10280_), .Y(_10281_));
NAND_g _32437_ (.A(_13409_), .B(_10281_), .Y(_10282_));
NAND_g _32438_ (.A(pcpi_rs1[17]), .B(_13416_), .Y(_10283_));
AND_g _32439_ (.A(_10282_), .B(_10283_), .Y(_10284_));
NAND_g _32440_ (.A(_10274_), .B(_10284_), .Y(_10285_));
NOR_g _32441_ (.A(_10270_), .B(_10285_), .Y(_10286_));
NOR_g _32442_ (.A(_10963_), .B(_10286_), .Y(_00009_[17]));
NAND_g _32443_ (.A(reg_pc[18]), .B(decoded_imm[18]), .Y(_10287_));
XOR_g _32444_ (.A(reg_pc[18]), .B(decoded_imm[18]), .Y(_10288_));
AND_g _32445_ (.A(_10263_), .B(_10264_), .Y(_10289_));
NOR_g _32446_ (.A(_10265_), .B(_10289_), .Y(_10290_));
NAND_g _32447_ (.A(_10288_), .B(_10290_), .Y(_10291_));
NOR_g _32448_ (.A(_10288_), .B(_10290_), .Y(_10292_));
NOR_g _32449_ (.A(_11272_), .B(_10292_), .Y(_10293_));
NAND_g _32450_ (.A(_10291_), .B(_10293_), .Y(_10294_));
AND_g _32451_ (.A(latched_is_lu), .B(mem_rdata[18]), .Y(_10295_));
NAND_g _32452_ (.A(_03961_), .B(_10295_), .Y(_10296_));
NAND_g _32453_ (.A(_10246_), .B(_10296_), .Y(_10297_));
NAND_g _32454_ (.A(_09824_), .B(_10297_), .Y(_10298_));
NAND_g _32455_ (.A(count_instr[18]), .B(instr_rdinstr), .Y(_10299_));
NAND_g _32456_ (.A(instr_rdcycleh), .B(count_cycle[50]), .Y(_10300_));
AND_g _32457_ (.A(_10299_), .B(_10300_), .Y(_10301_));
NAND_g _32458_ (.A(instr_rdcycle), .B(count_cycle[18]), .Y(_10302_));
NAND_g _32459_ (.A(count_instr[50]), .B(instr_rdinstrh), .Y(_10303_));
AND_g _32460_ (.A(_10302_), .B(_10303_), .Y(_10304_));
NAND_g _32461_ (.A(_10301_), .B(_10304_), .Y(_10305_));
NAND_g _32462_ (.A(_13409_), .B(_10305_), .Y(_10306_));
NAND_g _32463_ (.A(pcpi_rs1[18]), .B(_13416_), .Y(_10307_));
AND_g _32464_ (.A(_10306_), .B(_10307_), .Y(_10308_));
AND_g _32465_ (.A(_10298_), .B(_10308_), .Y(_10309_));
NAND_g _32466_ (.A(_10294_), .B(_10309_), .Y(_10310_));
AND_g _32467_ (.A(resetn), .B(_10310_), .Y(_00009_[18]));
AND_g _32468_ (.A(_10287_), .B(_10291_), .Y(_10311_));
NAND_g _32469_ (.A(reg_pc[19]), .B(decoded_imm[19]), .Y(_10312_));
NOR_g _32470_ (.A(reg_pc[19]), .B(decoded_imm[19]), .Y(_10313_));
XNOR_g _32471_ (.A(reg_pc[19]), .B(decoded_imm[19]), .Y(_10314_));
NOR_g _32472_ (.A(_10311_), .B(_10314_), .Y(_10315_));
NAND_g _32473_ (.A(_10311_), .B(_10314_), .Y(_10316_));
NAND_g _32474_ (.A(_11271_), .B(_10316_), .Y(_10317_));
NOR_g _32475_ (.A(_10315_), .B(_10317_), .Y(_10318_));
AND_g _32476_ (.A(latched_is_lu), .B(mem_rdata[19]), .Y(_10319_));
NAND_g _32477_ (.A(_03961_), .B(_10319_), .Y(_10320_));
NAND_g _32478_ (.A(_10246_), .B(_10320_), .Y(_10321_));
NAND_g _32479_ (.A(_09824_), .B(_10321_), .Y(_10322_));
NAND_g _32480_ (.A(count_instr[19]), .B(instr_rdinstr), .Y(_10323_));
NAND_g _32481_ (.A(instr_rdcycleh), .B(count_cycle[51]), .Y(_10324_));
AND_g _32482_ (.A(_10323_), .B(_10324_), .Y(_10325_));
NAND_g _32483_ (.A(count_instr[51]), .B(instr_rdinstrh), .Y(_10326_));
NAND_g _32484_ (.A(instr_rdcycle), .B(count_cycle[19]), .Y(_10327_));
AND_g _32485_ (.A(_10326_), .B(_10327_), .Y(_10328_));
NAND_g _32486_ (.A(_10325_), .B(_10328_), .Y(_10329_));
NAND_g _32487_ (.A(_13409_), .B(_10329_), .Y(_10330_));
NAND_g _32488_ (.A(pcpi_rs1[19]), .B(_13416_), .Y(_10331_));
AND_g _32489_ (.A(_10330_), .B(_10331_), .Y(_10332_));
NAND_g _32490_ (.A(_10322_), .B(_10332_), .Y(_10333_));
NOR_g _32491_ (.A(_10318_), .B(_10333_), .Y(_10334_));
NOR_g _32492_ (.A(_10963_), .B(_10334_), .Y(_00009_[19]));
NAND_g _32493_ (.A(reg_pc[20]), .B(decoded_imm[20]), .Y(_10335_));
XOR_g _32494_ (.A(reg_pc[20]), .B(decoded_imm[20]), .Y(_10336_));
AND_g _32495_ (.A(_10311_), .B(_10312_), .Y(_10337_));
NOR_g _32496_ (.A(_10313_), .B(_10337_), .Y(_10338_));
NAND_g _32497_ (.A(_10336_), .B(_10338_), .Y(_10339_));
NOR_g _32498_ (.A(_10336_), .B(_10338_), .Y(_10340_));
NOR_g _32499_ (.A(_11272_), .B(_10340_), .Y(_10341_));
NAND_g _32500_ (.A(_10339_), .B(_10341_), .Y(_10342_));
AND_g _32501_ (.A(latched_is_lu), .B(mem_rdata[20]), .Y(_10343_));
NAND_g _32502_ (.A(_03961_), .B(_10343_), .Y(_10344_));
NAND_g _32503_ (.A(_10246_), .B(_10344_), .Y(_10345_));
NAND_g _32504_ (.A(_09824_), .B(_10345_), .Y(_10346_));
NAND_g _32505_ (.A(pcpi_rs1[20]), .B(_13416_), .Y(_10347_));
NAND_g _32506_ (.A(count_instr[20]), .B(instr_rdinstr), .Y(_10348_));
NAND_g _32507_ (.A(instr_rdcycleh), .B(count_cycle[52]), .Y(_10349_));
AND_g _32508_ (.A(_10348_), .B(_10349_), .Y(_10350_));
NAND_g _32509_ (.A(instr_rdcycle), .B(count_cycle[20]), .Y(_10351_));
NAND_g _32510_ (.A(count_instr[52]), .B(instr_rdinstrh), .Y(_10352_));
AND_g _32511_ (.A(_10351_), .B(_10352_), .Y(_10353_));
NAND_g _32512_ (.A(_10350_), .B(_10353_), .Y(_10354_));
NAND_g _32513_ (.A(_13409_), .B(_10354_), .Y(_10355_));
AND_g _32514_ (.A(_10347_), .B(_10355_), .Y(_10356_));
AND_g _32515_ (.A(_10346_), .B(_10356_), .Y(_10357_));
NAND_g _32516_ (.A(_10342_), .B(_10357_), .Y(_10358_));
AND_g _32517_ (.A(resetn), .B(_10358_), .Y(_00009_[20]));
AND_g _32518_ (.A(_10335_), .B(_10339_), .Y(_10359_));
NAND_g _32519_ (.A(reg_pc[21]), .B(decoded_imm[21]), .Y(_10360_));
NOR_g _32520_ (.A(reg_pc[21]), .B(decoded_imm[21]), .Y(_10361_));
XNOR_g _32521_ (.A(reg_pc[21]), .B(decoded_imm[21]), .Y(_10362_));
NOR_g _32522_ (.A(_10359_), .B(_10362_), .Y(_10363_));
NAND_g _32523_ (.A(_10359_), .B(_10362_), .Y(_10364_));
AND_g _32524_ (.A(latched_is_lu), .B(mem_rdata[21]), .Y(_10365_));
NAND_g _32525_ (.A(_03961_), .B(_10365_), .Y(_10366_));
NAND_g _32526_ (.A(_10246_), .B(_10366_), .Y(_10367_));
NAND_g _32527_ (.A(_09824_), .B(_10367_), .Y(_10368_));
NAND_g _32528_ (.A(pcpi_rs1[21]), .B(_13416_), .Y(_10369_));
NAND_g _32529_ (.A(count_instr[21]), .B(instr_rdinstr), .Y(_10370_));
NAND_g _32530_ (.A(instr_rdcycleh), .B(count_cycle[53]), .Y(_10371_));
AND_g _32531_ (.A(_10370_), .B(_10371_), .Y(_10372_));
NAND_g _32532_ (.A(count_instr[53]), .B(instr_rdinstrh), .Y(_10373_));
NAND_g _32533_ (.A(instr_rdcycle), .B(count_cycle[21]), .Y(_10374_));
AND_g _32534_ (.A(_10373_), .B(_10374_), .Y(_10375_));
NAND_g _32535_ (.A(_10372_), .B(_10375_), .Y(_10376_));
NAND_g _32536_ (.A(_13409_), .B(_10376_), .Y(_10377_));
AND_g _32537_ (.A(_10369_), .B(_10377_), .Y(_10378_));
NOR_g _32538_ (.A(_11272_), .B(_10363_), .Y(_10379_));
NAND_g _32539_ (.A(_10364_), .B(_10379_), .Y(_10380_));
AND_g _32540_ (.A(_10378_), .B(_10380_), .Y(_10381_));
NAND_g _32541_ (.A(_10368_), .B(_10381_), .Y(_10382_));
AND_g _32542_ (.A(resetn), .B(_10382_), .Y(_00009_[21]));
NAND_g _32543_ (.A(reg_pc[22]), .B(decoded_imm[22]), .Y(_10383_));
XOR_g _32544_ (.A(reg_pc[22]), .B(decoded_imm[22]), .Y(_10384_));
AND_g _32545_ (.A(_10359_), .B(_10360_), .Y(_10385_));
NOR_g _32546_ (.A(_10361_), .B(_10385_), .Y(_10386_));
NAND_g _32547_ (.A(_10384_), .B(_10386_), .Y(_10387_));
NOR_g _32548_ (.A(_10384_), .B(_10386_), .Y(_10388_));
NOR_g _32549_ (.A(_11272_), .B(_10388_), .Y(_10389_));
NAND_g _32550_ (.A(_10387_), .B(_10389_), .Y(_10390_));
AND_g _32551_ (.A(latched_is_lu), .B(mem_rdata[22]), .Y(_10391_));
NAND_g _32552_ (.A(_03961_), .B(_10391_), .Y(_10392_));
NAND_g _32553_ (.A(_10246_), .B(_10392_), .Y(_10393_));
NAND_g _32554_ (.A(_09824_), .B(_10393_), .Y(_10394_));
NAND_g _32555_ (.A(pcpi_rs1[22]), .B(_13416_), .Y(_10395_));
NAND_g _32556_ (.A(count_instr[22]), .B(instr_rdinstr), .Y(_10396_));
NAND_g _32557_ (.A(instr_rdcycleh), .B(count_cycle[54]), .Y(_10397_));
AND_g _32558_ (.A(_10396_), .B(_10397_), .Y(_10398_));
NAND_g _32559_ (.A(instr_rdcycle), .B(count_cycle[22]), .Y(_10399_));
NAND_g _32560_ (.A(count_instr[54]), .B(instr_rdinstrh), .Y(_10400_));
AND_g _32561_ (.A(_10399_), .B(_10400_), .Y(_10401_));
NAND_g _32562_ (.A(_10398_), .B(_10401_), .Y(_10402_));
NAND_g _32563_ (.A(_13409_), .B(_10402_), .Y(_10403_));
AND_g _32564_ (.A(_10395_), .B(_10403_), .Y(_10404_));
AND_g _32565_ (.A(_10394_), .B(_10404_), .Y(_10405_));
NAND_g _32566_ (.A(_10390_), .B(_10405_), .Y(_10406_));
AND_g _32567_ (.A(resetn), .B(_10406_), .Y(_00009_[22]));
AND_g _32568_ (.A(latched_is_lu), .B(mem_rdata[23]), .Y(_10407_));
NAND_g _32569_ (.A(_03961_), .B(_10407_), .Y(_10408_));
NAND_g _32570_ (.A(_10246_), .B(_10408_), .Y(_10409_));
NAND_g _32571_ (.A(_09824_), .B(_10409_), .Y(_10410_));
NAND_g _32572_ (.A(count_instr[23]), .B(instr_rdinstr), .Y(_10411_));
NAND_g _32573_ (.A(instr_rdcycleh), .B(count_cycle[55]), .Y(_10412_));
AND_g _32574_ (.A(_10411_), .B(_10412_), .Y(_10413_));
NAND_g _32575_ (.A(instr_rdcycle), .B(count_cycle[23]), .Y(_10414_));
NAND_g _32576_ (.A(count_instr[55]), .B(instr_rdinstrh), .Y(_10415_));
AND_g _32577_ (.A(_10414_), .B(_10415_), .Y(_10416_));
NAND_g _32578_ (.A(_10413_), .B(_10416_), .Y(_10417_));
NAND_g _32579_ (.A(_13409_), .B(_10417_), .Y(_10418_));
NAND_g _32580_ (.A(pcpi_rs1[23]), .B(_13416_), .Y(_10419_));
AND_g _32581_ (.A(_10418_), .B(_10419_), .Y(_10420_));
AND_g _32582_ (.A(_10383_), .B(_10387_), .Y(_10421_));
NAND_g _32583_ (.A(reg_pc[23]), .B(decoded_imm[23]), .Y(_10422_));
NOR_g _32584_ (.A(reg_pc[23]), .B(decoded_imm[23]), .Y(_10423_));
XNOR_g _32585_ (.A(reg_pc[23]), .B(decoded_imm[23]), .Y(_10424_));
NOR_g _32586_ (.A(_10421_), .B(_10424_), .Y(_10425_));
NAND_g _32587_ (.A(_10421_), .B(_10424_), .Y(_10426_));
NOR_g _32588_ (.A(_11272_), .B(_10425_), .Y(_10427_));
NAND_g _32589_ (.A(_10426_), .B(_10427_), .Y(_10428_));
AND_g _32590_ (.A(_10420_), .B(_10428_), .Y(_10429_));
NAND_g _32591_ (.A(_10410_), .B(_10429_), .Y(_10430_));
AND_g _32592_ (.A(resetn), .B(_10430_), .Y(_00009_[23]));
NAND_g _32593_ (.A(reg_pc[24]), .B(decoded_imm[24]), .Y(_10431_));
XOR_g _32594_ (.A(reg_pc[24]), .B(decoded_imm[24]), .Y(_10432_));
AND_g _32595_ (.A(_10421_), .B(_10422_), .Y(_10433_));
NOR_g _32596_ (.A(_10423_), .B(_10433_), .Y(_10434_));
NAND_g _32597_ (.A(_10432_), .B(_10434_), .Y(_10435_));
NOR_g _32598_ (.A(_10432_), .B(_10434_), .Y(_10436_));
NOR_g _32599_ (.A(_11272_), .B(_10436_), .Y(_10437_));
NAND_g _32600_ (.A(_10435_), .B(_10437_), .Y(_10438_));
AND_g _32601_ (.A(latched_is_lu), .B(mem_rdata[24]), .Y(_10439_));
NAND_g _32602_ (.A(_03961_), .B(_10439_), .Y(_10440_));
NAND_g _32603_ (.A(_10246_), .B(_10440_), .Y(_10441_));
NAND_g _32604_ (.A(_09824_), .B(_10441_), .Y(_10442_));
NAND_g _32605_ (.A(count_instr[24]), .B(instr_rdinstr), .Y(_10443_));
NAND_g _32606_ (.A(instr_rdcycleh), .B(count_cycle[56]), .Y(_10444_));
AND_g _32607_ (.A(_10443_), .B(_10444_), .Y(_10445_));
NAND_g _32608_ (.A(instr_rdcycle), .B(count_cycle[24]), .Y(_10446_));
NAND_g _32609_ (.A(count_instr[56]), .B(instr_rdinstrh), .Y(_10447_));
AND_g _32610_ (.A(_10446_), .B(_10447_), .Y(_10448_));
NAND_g _32611_ (.A(_10445_), .B(_10448_), .Y(_10449_));
NAND_g _32612_ (.A(_13409_), .B(_10449_), .Y(_10450_));
NAND_g _32613_ (.A(pcpi_rs1[24]), .B(_13416_), .Y(_10451_));
AND_g _32614_ (.A(_10450_), .B(_10451_), .Y(_10452_));
AND_g _32615_ (.A(_10442_), .B(_10452_), .Y(_10453_));
NAND_g _32616_ (.A(_10438_), .B(_10453_), .Y(_10454_));
AND_g _32617_ (.A(resetn), .B(_10454_), .Y(_00009_[24]));
AND_g _32618_ (.A(_10431_), .B(_10435_), .Y(_10455_));
NAND_g _32619_ (.A(reg_pc[25]), .B(decoded_imm[25]), .Y(_10456_));
NOR_g _32620_ (.A(reg_pc[25]), .B(decoded_imm[25]), .Y(_10457_));
XNOR_g _32621_ (.A(reg_pc[25]), .B(decoded_imm[25]), .Y(_10458_));
NOR_g _32622_ (.A(_10455_), .B(_10458_), .Y(_10459_));
NAND_g _32623_ (.A(_10455_), .B(_10458_), .Y(_10460_));
NAND_g _32624_ (.A(_11271_), .B(_10460_), .Y(_10461_));
NOR_g _32625_ (.A(_10459_), .B(_10461_), .Y(_10462_));
AND_g _32626_ (.A(latched_is_lu), .B(mem_rdata[25]), .Y(_10463_));
NAND_g _32627_ (.A(_03961_), .B(_10463_), .Y(_10464_));
NAND_g _32628_ (.A(_10246_), .B(_10464_), .Y(_10465_));
NAND_g _32629_ (.A(_09824_), .B(_10465_), .Y(_10466_));
NAND_g _32630_ (.A(count_instr[25]), .B(instr_rdinstr), .Y(_10467_));
NAND_g _32631_ (.A(instr_rdcycleh), .B(count_cycle[57]), .Y(_10468_));
AND_g _32632_ (.A(_10467_), .B(_10468_), .Y(_10469_));
NAND_g _32633_ (.A(count_instr[57]), .B(instr_rdinstrh), .Y(_10470_));
NAND_g _32634_ (.A(instr_rdcycle), .B(count_cycle[25]), .Y(_10471_));
AND_g _32635_ (.A(_10470_), .B(_10471_), .Y(_10472_));
NAND_g _32636_ (.A(_10469_), .B(_10472_), .Y(_10473_));
NAND_g _32637_ (.A(_13409_), .B(_10473_), .Y(_10474_));
NAND_g _32638_ (.A(pcpi_rs1[25]), .B(_13416_), .Y(_10475_));
AND_g _32639_ (.A(_10474_), .B(_10475_), .Y(_10476_));
NAND_g _32640_ (.A(_10466_), .B(_10476_), .Y(_10477_));
NOR_g _32641_ (.A(_10462_), .B(_10477_), .Y(_10478_));
NOR_g _32642_ (.A(_10963_), .B(_10478_), .Y(_00009_[25]));
NAND_g _32643_ (.A(reg_pc[26]), .B(decoded_imm[26]), .Y(_10479_));
XOR_g _32644_ (.A(reg_pc[26]), .B(decoded_imm[26]), .Y(_10480_));
AND_g _32645_ (.A(_10455_), .B(_10456_), .Y(_10481_));
NOR_g _32646_ (.A(_10457_), .B(_10481_), .Y(_10482_));
NAND_g _32647_ (.A(_10480_), .B(_10482_), .Y(_10483_));
NOR_g _32648_ (.A(_10480_), .B(_10482_), .Y(_10484_));
NOR_g _32649_ (.A(_11272_), .B(_10484_), .Y(_10485_));
NAND_g _32650_ (.A(_10483_), .B(_10485_), .Y(_10486_));
AND_g _32651_ (.A(latched_is_lu), .B(mem_rdata[26]), .Y(_10487_));
NAND_g _32652_ (.A(_03961_), .B(_10487_), .Y(_10488_));
NAND_g _32653_ (.A(_10246_), .B(_10488_), .Y(_10489_));
NAND_g _32654_ (.A(_09824_), .B(_10489_), .Y(_10490_));
NAND_g _32655_ (.A(count_instr[26]), .B(instr_rdinstr), .Y(_10491_));
NAND_g _32656_ (.A(instr_rdcycleh), .B(count_cycle[58]), .Y(_10492_));
AND_g _32657_ (.A(_10491_), .B(_10492_), .Y(_10493_));
NAND_g _32658_ (.A(instr_rdcycle), .B(count_cycle[26]), .Y(_10494_));
NAND_g _32659_ (.A(count_instr[58]), .B(instr_rdinstrh), .Y(_10495_));
AND_g _32660_ (.A(_10494_), .B(_10495_), .Y(_10496_));
NAND_g _32661_ (.A(_10493_), .B(_10496_), .Y(_10497_));
NAND_g _32662_ (.A(_13409_), .B(_10497_), .Y(_10498_));
NAND_g _32663_ (.A(pcpi_rs1[26]), .B(_13416_), .Y(_10499_));
AND_g _32664_ (.A(_10498_), .B(_10499_), .Y(_10500_));
AND_g _32665_ (.A(_10490_), .B(_10500_), .Y(_10501_));
NAND_g _32666_ (.A(_10486_), .B(_10501_), .Y(_10502_));
AND_g _32667_ (.A(resetn), .B(_10502_), .Y(_00009_[26]));
AND_g _32668_ (.A(_10479_), .B(_10483_), .Y(_10503_));
NAND_g _32669_ (.A(reg_pc[27]), .B(decoded_imm[27]), .Y(_10504_));
NOR_g _32670_ (.A(reg_pc[27]), .B(decoded_imm[27]), .Y(_10505_));
XOR_g _32671_ (.A(reg_pc[27]), .B(decoded_imm[27]), .Y(_10506_));
XNOR_g _32672_ (.A(_10503_), .B(_10506_), .Y(_10507_));
NAND_g _32673_ (.A(_02563_), .B(_10507_), .Y(_10508_));
AND_g _32674_ (.A(latched_is_lu), .B(mem_rdata[27]), .Y(_10509_));
NAND_g _32675_ (.A(_03961_), .B(_10509_), .Y(_10510_));
NAND_g _32676_ (.A(_10246_), .B(_10510_), .Y(_10511_));
NAND_g _32677_ (.A(_09824_), .B(_10511_), .Y(_10512_));
NAND_g _32678_ (.A(pcpi_rs1[27]), .B(_13416_), .Y(_10513_));
NAND_g _32679_ (.A(count_instr[27]), .B(instr_rdinstr), .Y(_10514_));
NAND_g _32680_ (.A(instr_rdcycleh), .B(count_cycle[59]), .Y(_10515_));
AND_g _32681_ (.A(_10514_), .B(_10515_), .Y(_10516_));
NAND_g _32682_ (.A(instr_rdcycle), .B(count_cycle[27]), .Y(_10517_));
NAND_g _32683_ (.A(count_instr[59]), .B(instr_rdinstrh), .Y(_10518_));
AND_g _32684_ (.A(_10517_), .B(_10518_), .Y(_10519_));
NAND_g _32685_ (.A(_10516_), .B(_10519_), .Y(_10520_));
NAND_g _32686_ (.A(_13409_), .B(_10520_), .Y(_10521_));
AND_g _32687_ (.A(_10512_), .B(_10521_), .Y(_10522_));
NAND_g _32688_ (.A(_10513_), .B(_10522_), .Y(_10523_));
NAND_g _32689_ (.A(resetn), .B(_10523_), .Y(_10524_));
NAND_g _32690_ (.A(_10508_), .B(_10524_), .Y(_00009_[27]));
NAND_g _32691_ (.A(reg_pc[28]), .B(decoded_imm[28]), .Y(_10525_));
XOR_g _32692_ (.A(reg_pc[28]), .B(decoded_imm[28]), .Y(_10526_));
AND_g _32693_ (.A(_10503_), .B(_10504_), .Y(_10527_));
NOR_g _32694_ (.A(_10505_), .B(_10527_), .Y(_10528_));
NAND_g _32695_ (.A(_10526_), .B(_10528_), .Y(_10529_));
NOR_g _32696_ (.A(_10526_), .B(_10528_), .Y(_10530_));
NOR_g _32697_ (.A(_11272_), .B(_10530_), .Y(_10531_));
NAND_g _32698_ (.A(_10529_), .B(_10531_), .Y(_10532_));
AND_g _32699_ (.A(latched_is_lu), .B(mem_rdata[28]), .Y(_10533_));
NAND_g _32700_ (.A(_03961_), .B(_10533_), .Y(_10534_));
NAND_g _32701_ (.A(_10246_), .B(_10534_), .Y(_10535_));
NAND_g _32702_ (.A(_09824_), .B(_10535_), .Y(_10536_));
NAND_g _32703_ (.A(pcpi_rs1[28]), .B(_13416_), .Y(_10537_));
NAND_g _32704_ (.A(count_instr[28]), .B(instr_rdinstr), .Y(_10538_));
NAND_g _32705_ (.A(instr_rdcycleh), .B(count_cycle[60]), .Y(_10539_));
AND_g _32706_ (.A(_10538_), .B(_10539_), .Y(_10540_));
NAND_g _32707_ (.A(count_instr[60]), .B(instr_rdinstrh), .Y(_10541_));
NAND_g _32708_ (.A(instr_rdcycle), .B(count_cycle[28]), .Y(_10542_));
AND_g _32709_ (.A(_10541_), .B(_10542_), .Y(_10543_));
NAND_g _32710_ (.A(_10540_), .B(_10543_), .Y(_10544_));
NAND_g _32711_ (.A(_13409_), .B(_10544_), .Y(_10545_));
AND_g _32712_ (.A(_10537_), .B(_10545_), .Y(_10546_));
AND_g _32713_ (.A(_10536_), .B(_10546_), .Y(_10547_));
NAND_g _32714_ (.A(_10532_), .B(_10547_), .Y(_10548_));
AND_g _32715_ (.A(resetn), .B(_10548_), .Y(_00009_[28]));
AND_g _32716_ (.A(latched_is_lu), .B(mem_rdata[29]), .Y(_10549_));
NAND_g _32717_ (.A(_03961_), .B(_10549_), .Y(_10550_));
NAND_g _32718_ (.A(_10246_), .B(_10550_), .Y(_10551_));
NAND_g _32719_ (.A(_09824_), .B(_10551_), .Y(_10552_));
NAND_g _32720_ (.A(count_instr[29]), .B(instr_rdinstr), .Y(_10553_));
NAND_g _32721_ (.A(instr_rdcycleh), .B(count_cycle[61]), .Y(_10554_));
AND_g _32722_ (.A(_10553_), .B(_10554_), .Y(_10555_));
NAND_g _32723_ (.A(instr_rdcycle), .B(count_cycle[29]), .Y(_10556_));
NAND_g _32724_ (.A(count_instr[61]), .B(instr_rdinstrh), .Y(_10557_));
AND_g _32725_ (.A(_10556_), .B(_10557_), .Y(_10558_));
NAND_g _32726_ (.A(_10555_), .B(_10558_), .Y(_10559_));
NAND_g _32727_ (.A(_13409_), .B(_10559_), .Y(_10560_));
NAND_g _32728_ (.A(pcpi_rs1[29]), .B(_13416_), .Y(_10561_));
AND_g _32729_ (.A(_10560_), .B(_10561_), .Y(_10562_));
NAND_g _32730_ (.A(_10552_), .B(_10562_), .Y(_10563_));
NAND_g _32731_ (.A(resetn), .B(_10563_), .Y(_10564_));
AND_g _32732_ (.A(_10525_), .B(_10529_), .Y(_10565_));
NAND_g _32733_ (.A(_10525_), .B(_10529_), .Y(_10566_));
NAND_g _32734_ (.A(reg_pc[29]), .B(decoded_imm[29]), .Y(_10567_));
XOR_g _32735_ (.A(reg_pc[29]), .B(decoded_imm[29]), .Y(_10568_));
XNOR_g _32736_ (.A(reg_pc[29]), .B(decoded_imm[29]), .Y(_10569_));
NAND_g _32737_ (.A(_10565_), .B(_10569_), .Y(_10570_));
NAND_g _32738_ (.A(_10566_), .B(_10568_), .Y(_10571_));
AND_g _32739_ (.A(_02563_), .B(_10571_), .Y(_10572_));
NAND_g _32740_ (.A(_10570_), .B(_10572_), .Y(_10573_));
NAND_g _32741_ (.A(_10564_), .B(_10573_), .Y(_00009_[29]));
AND_g _32742_ (.A(_10567_), .B(_10571_), .Y(_10574_));
NAND_g _32743_ (.A(_10567_), .B(_10571_), .Y(_10575_));
NAND_g _32744_ (.A(reg_pc[30]), .B(decoded_imm[30]), .Y(_10576_));
XOR_g _32745_ (.A(reg_pc[30]), .B(decoded_imm[30]), .Y(_10577_));
XNOR_g _32746_ (.A(reg_pc[30]), .B(decoded_imm[30]), .Y(_10578_));
NAND_g _32747_ (.A(_10575_), .B(_10577_), .Y(_10579_));
NAND_g _32748_ (.A(_10574_), .B(_10578_), .Y(_10580_));
AND_g _32749_ (.A(_11271_), .B(_10580_), .Y(_10581_));
NAND_g _32750_ (.A(_10579_), .B(_10581_), .Y(_10582_));
AND_g _32751_ (.A(latched_is_lu), .B(mem_rdata[30]), .Y(_10583_));
NAND_g _32752_ (.A(_03961_), .B(_10583_), .Y(_10584_));
NAND_g _32753_ (.A(_10246_), .B(_10584_), .Y(_10585_));
NAND_g _32754_ (.A(_09824_), .B(_10585_), .Y(_10586_));
NAND_g _32755_ (.A(count_instr[30]), .B(instr_rdinstr), .Y(_10587_));
NAND_g _32756_ (.A(instr_rdcycleh), .B(count_cycle[62]), .Y(_10588_));
AND_g _32757_ (.A(_10587_), .B(_10588_), .Y(_10589_));
NAND_g _32758_ (.A(count_instr[62]), .B(instr_rdinstrh), .Y(_10590_));
NAND_g _32759_ (.A(instr_rdcycle), .B(count_cycle[30]), .Y(_10591_));
AND_g _32760_ (.A(_10590_), .B(_10591_), .Y(_10592_));
NAND_g _32761_ (.A(_10589_), .B(_10592_), .Y(_10593_));
NAND_g _32762_ (.A(_13409_), .B(_10593_), .Y(_10594_));
NAND_g _32763_ (.A(pcpi_rs1[30]), .B(_13416_), .Y(_10595_));
AND_g _32764_ (.A(_10594_), .B(_10595_), .Y(_10596_));
AND_g _32765_ (.A(_10586_), .B(_10596_), .Y(_10597_));
NAND_g _32766_ (.A(_10582_), .B(_10597_), .Y(_10598_));
AND_g _32767_ (.A(resetn), .B(_10598_), .Y(_00009_[30]));
AND_g _32768_ (.A(_10576_), .B(_10579_), .Y(_10599_));
NAND_g _32769_ (.A(_10576_), .B(_10579_), .Y(_10600_));
XNOR_g _32770_ (.A(reg_pc[31]), .B(decoded_imm[31]), .Y(_10601_));
XOR_g _32771_ (.A(reg_pc[31]), .B(decoded_imm[31]), .Y(_10602_));
NAND_g _32772_ (.A(_10599_), .B(_10601_), .Y(_10603_));
NAND_g _32773_ (.A(_10600_), .B(_10602_), .Y(_10604_));
AND_g _32774_ (.A(_11271_), .B(_10604_), .Y(_10605_));
NAND_g _32775_ (.A(_10603_), .B(_10605_), .Y(_10606_));
AND_g _32776_ (.A(latched_is_lu), .B(mem_rdata[31]), .Y(_10607_));
NAND_g _32777_ (.A(_03961_), .B(_10607_), .Y(_10608_));
NAND_g _32778_ (.A(_10246_), .B(_10608_), .Y(_10609_));
NAND_g _32779_ (.A(_09824_), .B(_10609_), .Y(_10610_));
NAND_g _32780_ (.A(count_instr[31]), .B(instr_rdinstr), .Y(_10611_));
NAND_g _32781_ (.A(instr_rdcycleh), .B(count_cycle[63]), .Y(_10612_));
AND_g _32782_ (.A(_10611_), .B(_10612_), .Y(_10613_));
NAND_g _32783_ (.A(count_instr[63]), .B(instr_rdinstrh), .Y(_10614_));
NAND_g _32784_ (.A(instr_rdcycle), .B(count_cycle[31]), .Y(_10615_));
AND_g _32785_ (.A(_10614_), .B(_10615_), .Y(_10616_));
NAND_g _32786_ (.A(_10613_), .B(_10616_), .Y(_10617_));
NAND_g _32787_ (.A(_13409_), .B(_10617_), .Y(_10618_));
NAND_g _32788_ (.A(pcpi_rs1[31]), .B(_13416_), .Y(_10619_));
AND_g _32789_ (.A(_10618_), .B(_10619_), .Y(_10620_));
AND_g _32790_ (.A(_10610_), .B(_10620_), .Y(_10621_));
NAND_g _32791_ (.A(_10606_), .B(_10621_), .Y(_10622_));
AND_g _32792_ (.A(resetn), .B(_10622_), .Y(_00009_[31]));
XNOR_g _32793_ (.A(_11207_), .B(_13382_), .Y(_10623_));
NAND_g _32794_ (.A(_13389_), .B(_10623_), .Y(_10624_));
NAND_g _32795_ (.A(decoded_imm_j[11]), .B(_04777_), .Y(_10625_));
NAND_g _32796_ (.A(_10624_), .B(_10625_), .Y(_10626_));
NAND_g _32797_ (.A(resetn), .B(_10626_), .Y(_10627_));
NAND_g _32798_ (.A(_13835_), .B(_04805_), .Y(_10628_));
NAND_g _32799_ (.A(resetn), .B(_13840_), .Y(_10629_));
AND_g _32800_ (.A(_10628_), .B(_10629_), .Y(_10630_));
NAND_g _32801_ (.A(_10627_), .B(_10630_), .Y(_00010_[0]));
NAND_g _32802_ (.A(decoded_imm_j[1]), .B(_04777_), .Y(_10631_));
AND_g _32803_ (.A(reg_sh[1]), .B(_13384_), .Y(_10632_));
NAND_g _32804_ (.A(_13387_), .B(_10632_), .Y(_10633_));
AND_g _32805_ (.A(_10631_), .B(_10633_), .Y(_10634_));
AND_g _32806_ (.A(_13942_), .B(_10634_), .Y(_10635_));
NAND_g _32807_ (.A(_13941_), .B(_10635_), .Y(_10636_));
AND_g _32808_ (.A(resetn), .B(_10636_), .Y(_00010_[1]));
NAND_g _32809_ (.A(decoded_imm_j[2]), .B(_04777_), .Y(_10637_));
NOR_g _32810_ (.A(reg_sh[2]), .B(_13382_), .Y(_10638_));
NAND_g _32811_ (.A(_13387_), .B(_10638_), .Y(_10639_));
AND_g _32812_ (.A(_10637_), .B(_10639_), .Y(_10640_));
AND_g _32813_ (.A(_14047_), .B(_10640_), .Y(_10641_));
NAND_g _32814_ (.A(_14046_), .B(_10641_), .Y(_10642_));
AND_g _32815_ (.A(resetn), .B(_10642_), .Y(_00010_[2]));
NAND_g _32816_ (.A(reg_sh[2]), .B(reg_sh[3]), .Y(_10643_));
NAND_g _32817_ (.A(reg_sh[4]), .B(_13381_), .Y(_10644_));
NAND_g _32818_ (.A(_10643_), .B(_10644_), .Y(_10645_));
NAND_g _32819_ (.A(_13387_), .B(_10645_), .Y(_10646_));
NAND_g _32820_ (.A(decoded_imm_j[3]), .B(_04777_), .Y(_10647_));
NAND_g _32821_ (.A(_10646_), .B(_10647_), .Y(_10648_));
NAND_g _32822_ (.A(resetn), .B(_10648_), .Y(_10649_));
NAND_g _32823_ (.A(_14149_), .B(_04805_), .Y(_10650_));
NAND_g _32824_ (.A(resetn), .B(_14154_), .Y(_10651_));
AND_g _32825_ (.A(_10649_), .B(_10651_), .Y(_10652_));
NAND_g _32826_ (.A(_10650_), .B(_10652_), .Y(_00010_[3]));
NAND_g _32827_ (.A(_14253_), .B(_04805_), .Y(_10653_));
NOR_g _32828_ (.A(_11208_), .B(_13381_), .Y(_10654_));
NAND_g _32829_ (.A(_13387_), .B(_10654_), .Y(_10655_));
NAND_g _32830_ (.A(decoded_imm_j[4]), .B(_04777_), .Y(_10656_));
AND_g _32831_ (.A(_10655_), .B(_10656_), .Y(_10657_));
NAND_g _32832_ (.A(_14258_), .B(_10657_), .Y(_10658_));
NAND_g _32833_ (.A(resetn), .B(_10658_), .Y(_10659_));
NAND_g _32834_ (.A(_10653_), .B(_10659_), .Y(_00010_[4]));
NAND_g _32835_ (.A(dbg_rs2val_valid), .B(_11264_), .Y(_10660_));
AND_g _32836_ (.A(resetn), .B(_14358_), .Y(_10661_));
NOT_g _32837_ (.A(_10661_), .Y(_10662_));
NAND_g _32838_ (.A(_10660_), .B(_10662_), .Y(_00003_));
NAND_g _32839_ (.A(dbg_rs1val_valid), .B(_11264_), .Y(_10663_));
AND_g _32840_ (.A(resetn), .B(_05765_), .Y(_10664_));
NOT_g _32841_ (.A(_10664_), .Y(_10665_));
NAND_g _32842_ (.A(_10663_), .B(_10665_), .Y(_00001_));
AND_g _32843_ (.A(dbg_rs2val[0]), .B(_11264_), .Y(_10666_));
NAND_g _32844_ (.A(_13834_), .B(_04805_), .Y(_10667_));
NAND_g _32845_ (.A(_13727_), .B(_10667_), .Y(_10668_));
NAND_g _32846_ (.A(_10666_), .B(_10668_), .Y(_10669_));
NAND_g _32847_ (.A(_10630_), .B(_10669_), .Y(_00002_[0]));
AND_g _32848_ (.A(dbg_rs2val[1]), .B(_11264_), .Y(_10670_));
NAND_g _32849_ (.A(_13834_), .B(_10670_), .Y(_10671_));
NAND_g _32850_ (.A(_13948_), .B(_10671_), .Y(_10672_));
NAND_g _32851_ (.A(_04805_), .B(_10672_), .Y(_10673_));
NAND_g _32852_ (.A(resetn), .B(_13943_), .Y(_10674_));
NAND_g _32853_ (.A(_13728_), .B(_10670_), .Y(_10675_));
AND_g _32854_ (.A(_10673_), .B(_10675_), .Y(_10676_));
NAND_g _32855_ (.A(_10674_), .B(_10676_), .Y(_00002_[1]));
AND_g _32856_ (.A(dbg_rs2val[2]), .B(_11264_), .Y(_10677_));
NAND_g _32857_ (.A(_10668_), .B(_10677_), .Y(_10678_));
NOR_g _32858_ (.A(_10963_), .B(_14047_), .Y(_10679_));
AND_g _32859_ (.A(_13833_), .B(_04805_), .Y(_10680_));
AND_g _32860_ (.A(_14045_), .B(_10680_), .Y(_10681_));
NOR_g _32861_ (.A(_10679_), .B(_10681_), .Y(_10682_));
NAND_g _32862_ (.A(_10678_), .B(_10682_), .Y(_00002_[2]));
AND_g _32863_ (.A(dbg_rs2val[3]), .B(_11264_), .Y(_10683_));
NAND_g _32864_ (.A(_10668_), .B(_10683_), .Y(_10684_));
AND_g _32865_ (.A(_10650_), .B(_10651_), .Y(_10685_));
NAND_g _32866_ (.A(_10684_), .B(_10685_), .Y(_00002_[3]));
AND_g _32867_ (.A(dbg_rs2val[4]), .B(_11264_), .Y(_10686_));
NAND_g _32868_ (.A(_10668_), .B(_10686_), .Y(_10687_));
NAND_g _32869_ (.A(resetn), .B(_14259_), .Y(_10688_));
AND_g _32870_ (.A(_10653_), .B(_10688_), .Y(_10689_));
NAND_g _32871_ (.A(_10687_), .B(_10689_), .Y(_00002_[4]));
AND_g _32872_ (.A(dbg_rs2val[5]), .B(_11264_), .Y(_10690_));
NAND_g _32873_ (.A(_10668_), .B(_10690_), .Y(_10691_));
NAND_g _32874_ (.A(_14357_), .B(_10661_), .Y(_10692_));
NAND_g _32875_ (.A(_10691_), .B(_10692_), .Y(_00002_[5]));
AND_g _32876_ (.A(dbg_rs2val[6]), .B(_11264_), .Y(_10693_));
NAND_g _32877_ (.A(_10668_), .B(_10693_), .Y(_10694_));
NAND_g _32878_ (.A(_14459_), .B(_10661_), .Y(_10695_));
NAND_g _32879_ (.A(_10694_), .B(_10695_), .Y(_00002_[6]));
AND_g _32880_ (.A(dbg_rs2val[7]), .B(_11264_), .Y(_10696_));
NAND_g _32881_ (.A(_10668_), .B(_10696_), .Y(_10697_));
NAND_g _32882_ (.A(_14560_), .B(_10661_), .Y(_10698_));
NAND_g _32883_ (.A(_10697_), .B(_10698_), .Y(_00002_[7]));
AND_g _32884_ (.A(dbg_rs2val[8]), .B(_11264_), .Y(_10699_));
NAND_g _32885_ (.A(_10668_), .B(_10699_), .Y(_10700_));
NAND_g _32886_ (.A(_14661_), .B(_10661_), .Y(_10701_));
NAND_g _32887_ (.A(_10700_), .B(_10701_), .Y(_00002_[8]));
AND_g _32888_ (.A(dbg_rs2val[9]), .B(_11264_), .Y(_10702_));
NAND_g _32889_ (.A(_10668_), .B(_10702_), .Y(_10703_));
NAND_g _32890_ (.A(_14761_), .B(_10661_), .Y(_10704_));
NAND_g _32891_ (.A(_10703_), .B(_10704_), .Y(_00002_[9]));
AND_g _32892_ (.A(dbg_rs2val[10]), .B(_11264_), .Y(_10705_));
NAND_g _32893_ (.A(_10668_), .B(_10705_), .Y(_10706_));
NOR_g _32894_ (.A(_10963_), .B(_14867_), .Y(_10707_));
NOR_g _32895_ (.A(_14863_), .B(_04806_), .Y(_10708_));
NOR_g _32896_ (.A(_10707_), .B(_10708_), .Y(_10709_));
NAND_g _32897_ (.A(_10706_), .B(_10709_), .Y(_00002_[10]));
AND_g _32898_ (.A(dbg_rs2val[11]), .B(_11264_), .Y(_10710_));
NAND_g _32899_ (.A(_10668_), .B(_10710_), .Y(_10711_));
NAND_g _32900_ (.A(_14964_), .B(_10661_), .Y(_10712_));
NAND_g _32901_ (.A(_10711_), .B(_10712_), .Y(_00002_[11]));
AND_g _32902_ (.A(dbg_rs2val[12]), .B(_11264_), .Y(_10713_));
NAND_g _32903_ (.A(_10668_), .B(_10713_), .Y(_10714_));
NAND_g _32904_ (.A(_15064_), .B(_10661_), .Y(_10715_));
NAND_g _32905_ (.A(_10714_), .B(_10715_), .Y(_00002_[12]));
AND_g _32906_ (.A(dbg_rs2val[13]), .B(_11264_), .Y(_10716_));
NAND_g _32907_ (.A(_10668_), .B(_10716_), .Y(_10717_));
AND_g _32908_ (.A(resetn), .B(_15169_), .Y(_10718_));
NOR_g _32909_ (.A(_15165_), .B(_04806_), .Y(_10719_));
NOR_g _32910_ (.A(_10718_), .B(_10719_), .Y(_10720_));
NAND_g _32911_ (.A(_10717_), .B(_10720_), .Y(_00002_[13]));
AND_g _32912_ (.A(dbg_rs2val[14]), .B(_11264_), .Y(_10721_));
NAND_g _32913_ (.A(_10668_), .B(_10721_), .Y(_10722_));
NAND_g _32914_ (.A(_15267_), .B(_10661_), .Y(_10723_));
NAND_g _32915_ (.A(_10722_), .B(_10723_), .Y(_00002_[14]));
AND_g _32916_ (.A(dbg_rs2val[15]), .B(_11264_), .Y(_10724_));
NAND_g _32917_ (.A(_10668_), .B(_10724_), .Y(_10725_));
NAND_g _32918_ (.A(_15368_), .B(_10661_), .Y(_10726_));
NAND_g _32919_ (.A(_10725_), .B(_10726_), .Y(_00002_[15]));
AND_g _32920_ (.A(dbg_rs2val[16]), .B(_11264_), .Y(_10727_));
NAND_g _32921_ (.A(_10668_), .B(_10727_), .Y(_10728_));
NAND_g _32922_ (.A(_15468_), .B(_10661_), .Y(_10729_));
NAND_g _32923_ (.A(_10728_), .B(_10729_), .Y(_00002_[16]));
AND_g _32924_ (.A(dbg_rs2val[17]), .B(_11264_), .Y(_10730_));
NAND_g _32925_ (.A(_10668_), .B(_10730_), .Y(_10731_));
NAND_g _32926_ (.A(_15569_), .B(_10661_), .Y(_10732_));
NAND_g _32927_ (.A(_10731_), .B(_10732_), .Y(_00002_[17]));
AND_g _32928_ (.A(dbg_rs2val[18]), .B(_11264_), .Y(_10733_));
NAND_g _32929_ (.A(_10668_), .B(_10733_), .Y(_10734_));
NAND_g _32930_ (.A(_15669_), .B(_10661_), .Y(_10735_));
NAND_g _32931_ (.A(_10734_), .B(_10735_), .Y(_00002_[18]));
AND_g _32932_ (.A(dbg_rs2val[19]), .B(_11264_), .Y(_10736_));
NAND_g _32933_ (.A(_10668_), .B(_10736_), .Y(_10737_));
NAND_g _32934_ (.A(_15770_), .B(_10661_), .Y(_10738_));
NAND_g _32935_ (.A(_10737_), .B(_10738_), .Y(_00002_[19]));
AND_g _32936_ (.A(dbg_rs2val[20]), .B(_11264_), .Y(_10739_));
NAND_g _32937_ (.A(_10668_), .B(_10739_), .Y(_10740_));
NAND_g _32938_ (.A(_15870_), .B(_10661_), .Y(_10741_));
NAND_g _32939_ (.A(_10740_), .B(_10741_), .Y(_00002_[20]));
AND_g _32940_ (.A(dbg_rs2val[21]), .B(_11264_), .Y(_10742_));
NAND_g _32941_ (.A(_10668_), .B(_10742_), .Y(_10743_));
NAND_g _32942_ (.A(_15970_), .B(_10661_), .Y(_10744_));
NAND_g _32943_ (.A(_10743_), .B(_10744_), .Y(_00002_[21]));
AND_g _32944_ (.A(dbg_rs2val[22]), .B(_11264_), .Y(_10745_));
NAND_g _32945_ (.A(_13834_), .B(_10745_), .Y(_10746_));
NAND_g _32946_ (.A(_16072_), .B(_10746_), .Y(_10747_));
NAND_g _32947_ (.A(_04805_), .B(_10747_), .Y(_10748_));
NAND_g _32948_ (.A(resetn), .B(_16076_), .Y(_10749_));
NAND_g _32949_ (.A(_13728_), .B(_10745_), .Y(_10750_));
AND_g _32950_ (.A(_10749_), .B(_10750_), .Y(_10751_));
NAND_g _32951_ (.A(_10748_), .B(_10751_), .Y(_00002_[22]));
AND_g _32952_ (.A(dbg_rs2val[23]), .B(_11264_), .Y(_10752_));
NAND_g _32953_ (.A(_10668_), .B(_10752_), .Y(_10753_));
NAND_g _32954_ (.A(_16173_), .B(_10661_), .Y(_10754_));
NAND_g _32955_ (.A(_10753_), .B(_10754_), .Y(_00002_[23]));
AND_g _32956_ (.A(dbg_rs2val[24]), .B(_11264_), .Y(_10755_));
NAND_g _32957_ (.A(_10668_), .B(_10755_), .Y(_10756_));
NAND_g _32958_ (.A(_16273_), .B(_10661_), .Y(_10757_));
NAND_g _32959_ (.A(_10756_), .B(_10757_), .Y(_00002_[24]));
AND_g _32960_ (.A(dbg_rs2val[25]), .B(_11264_), .Y(_10758_));
NAND_g _32961_ (.A(_13834_), .B(_10758_), .Y(_10759_));
NAND_g _32962_ (.A(_16374_), .B(_10759_), .Y(_10760_));
NAND_g _32963_ (.A(_04805_), .B(_10760_), .Y(_10761_));
NAND_g _32964_ (.A(resetn), .B(_16378_), .Y(_10762_));
NAND_g _32965_ (.A(_13728_), .B(_10758_), .Y(_10763_));
AND_g _32966_ (.A(_10762_), .B(_10763_), .Y(_10764_));
NAND_g _32967_ (.A(_10761_), .B(_10764_), .Y(_00002_[25]));
AND_g _32968_ (.A(dbg_rs2val[26]), .B(_11264_), .Y(_10765_));
NAND_g _32969_ (.A(_10668_), .B(_10765_), .Y(_10766_));
NAND_g _32970_ (.A(_01714_), .B(_10661_), .Y(_10767_));
NAND_g _32971_ (.A(_10766_), .B(_10767_), .Y(_00002_[26]));
AND_g _32972_ (.A(dbg_rs2val[27]), .B(_11264_), .Y(_10768_));
NAND_g _32973_ (.A(_10668_), .B(_10768_), .Y(_10769_));
NAND_g _32974_ (.A(_01815_), .B(_10661_), .Y(_10770_));
NAND_g _32975_ (.A(_10769_), .B(_10770_), .Y(_00002_[27]));
AND_g _32976_ (.A(dbg_rs2val[28]), .B(_11264_), .Y(_10771_));
NAND_g _32977_ (.A(_10668_), .B(_10771_), .Y(_10772_));
NAND_g _32978_ (.A(_01915_), .B(_10661_), .Y(_10773_));
NAND_g _32979_ (.A(_10772_), .B(_10773_), .Y(_00002_[28]));
AND_g _32980_ (.A(dbg_rs2val[29]), .B(_11264_), .Y(_10774_));
NAND_g _32981_ (.A(_13834_), .B(_10774_), .Y(_10775_));
NAND_g _32982_ (.A(_02016_), .B(_10775_), .Y(_10776_));
NAND_g _32983_ (.A(_04805_), .B(_10776_), .Y(_10777_));
NAND_g _32984_ (.A(resetn), .B(_02020_), .Y(_10778_));
NAND_g _32985_ (.A(_13728_), .B(_10774_), .Y(_10779_));
AND_g _32986_ (.A(_10778_), .B(_10779_), .Y(_10780_));
NAND_g _32987_ (.A(_10777_), .B(_10780_), .Y(_00002_[29]));
AND_g _32988_ (.A(dbg_rs2val[30]), .B(_11264_), .Y(_10781_));
NAND_g _32989_ (.A(_10668_), .B(_10781_), .Y(_10782_));
NOR_g _32990_ (.A(_10963_), .B(_02122_), .Y(_10783_));
NOR_g _32991_ (.A(_02118_), .B(_04806_), .Y(_10784_));
NOR_g _32992_ (.A(_10783_), .B(_10784_), .Y(_10785_));
NAND_g _32993_ (.A(_10782_), .B(_10785_), .Y(_00002_[30]));
AND_g _32994_ (.A(dbg_rs2val[31]), .B(_11264_), .Y(_10786_));
NAND_g _32995_ (.A(_10668_), .B(_10786_), .Y(_10787_));
NAND_g _32996_ (.A(_02219_), .B(_10661_), .Y(_10788_));
NAND_g _32997_ (.A(_10787_), .B(_10788_), .Y(_00002_[31]));
NAND_g _32998_ (.A(resetn), .B(_04971_), .Y(_10789_));
NOR_g _32999_ (.A(launch_next_insn), .B(_10664_), .Y(_10790_));
NAND_g _33000_ (.A(dbg_rs1val[0]), .B(_10790_), .Y(_10791_));
NAND_g _33001_ (.A(_10789_), .B(_10791_), .Y(_00000_[0]));
NAND_g _33002_ (.A(resetn), .B(_05079_), .Y(_10792_));
NAND_g _33003_ (.A(dbg_rs1val[1]), .B(_10790_), .Y(_10793_));
NAND_g _33004_ (.A(_10792_), .B(_10793_), .Y(_00000_[1]));
NAND_g _33005_ (.A(resetn), .B(_05190_), .Y(_10794_));
NAND_g _33006_ (.A(dbg_rs1val[2]), .B(_10790_), .Y(_10795_));
NAND_g _33007_ (.A(_10794_), .B(_10795_), .Y(_00000_[2]));
NAND_g _33008_ (.A(resetn), .B(_05301_), .Y(_10796_));
NAND_g _33009_ (.A(dbg_rs1val[3]), .B(_10790_), .Y(_10797_));
NAND_g _33010_ (.A(_10796_), .B(_10797_), .Y(_00000_[3]));
NAND_g _33011_ (.A(dbg_rs1val[4]), .B(_10790_), .Y(_10798_));
NAND_g _33012_ (.A(resetn), .B(_05413_), .Y(_10799_));
NAND_g _33013_ (.A(_10798_), .B(_10799_), .Y(_00000_[4]));
NAND_g _33014_ (.A(dbg_rs1val[5]), .B(_10790_), .Y(_10800_));
NAND_g _33015_ (.A(resetn), .B(_05525_), .Y(_10801_));
NAND_g _33016_ (.A(_10800_), .B(_10801_), .Y(_00000_[5]));
NAND_g _33017_ (.A(resetn), .B(_05636_), .Y(_10802_));
NAND_g _33018_ (.A(dbg_rs1val[6]), .B(_10790_), .Y(_10803_));
NAND_g _33019_ (.A(_10802_), .B(_10803_), .Y(_00000_[6]));
NAND_g _33020_ (.A(dbg_rs1val[7]), .B(_10790_), .Y(_10804_));
NAND_g _33021_ (.A(resetn), .B(_05750_), .Y(_10805_));
NAND_g _33022_ (.A(_10804_), .B(_10805_), .Y(_00000_[7]));
NAND_g _33023_ (.A(dbg_rs1val[8]), .B(_10790_), .Y(_10806_));
NAND_g _33024_ (.A(_05860_), .B(_10664_), .Y(_10807_));
NAND_g _33025_ (.A(_10806_), .B(_10807_), .Y(_00000_[8]));
NAND_g _33026_ (.A(dbg_rs1val[9]), .B(_10790_), .Y(_10808_));
NAND_g _33027_ (.A(resetn), .B(_05976_), .Y(_10809_));
NAND_g _33028_ (.A(_10808_), .B(_10809_), .Y(_00000_[9]));
NAND_g _33029_ (.A(dbg_rs1val[10]), .B(_10790_), .Y(_10810_));
NAND_g _33030_ (.A(_06097_), .B(_10664_), .Y(_10811_));
NAND_g _33031_ (.A(_10810_), .B(_10811_), .Y(_00000_[10]));
NAND_g _33032_ (.A(resetn), .B(_06201_), .Y(_10812_));
NAND_g _33033_ (.A(dbg_rs1val[11]), .B(_10790_), .Y(_10813_));
NAND_g _33034_ (.A(_10812_), .B(_10813_), .Y(_00000_[11]));
NAND_g _33035_ (.A(dbg_rs1val[12]), .B(_10790_), .Y(_10814_));
NAND_g _33036_ (.A(_06312_), .B(_10664_), .Y(_10815_));
NAND_g _33037_ (.A(_10814_), .B(_10815_), .Y(_00000_[12]));
NAND_g _33038_ (.A(dbg_rs1val[13]), .B(_10790_), .Y(_10816_));
NAND_g _33039_ (.A(_06436_), .B(_10664_), .Y(_10817_));
NAND_g _33040_ (.A(_10816_), .B(_10817_), .Y(_00000_[13]));
NAND_g _33041_ (.A(dbg_rs1val[14]), .B(_10790_), .Y(_10818_));
NAND_g _33042_ (.A(resetn), .B(_06535_), .Y(_10819_));
NAND_g _33043_ (.A(_10818_), .B(_10819_), .Y(_00000_[14]));
NAND_g _33044_ (.A(dbg_rs1val[15]), .B(_10790_), .Y(_10820_));
NAND_g _33045_ (.A(_06659_), .B(_10664_), .Y(_10821_));
NAND_g _33046_ (.A(_10820_), .B(_10821_), .Y(_00000_[15]));
NAND_g _33047_ (.A(dbg_rs1val[16]), .B(_10790_), .Y(_10822_));
NAND_g _33048_ (.A(_06770_), .B(_10664_), .Y(_10823_));
NAND_g _33049_ (.A(_10822_), .B(_10823_), .Y(_00000_[16]));
NAND_g _33050_ (.A(resetn), .B(_06869_), .Y(_10824_));
NAND_g _33051_ (.A(dbg_rs1val[17]), .B(_10790_), .Y(_10825_));
NAND_g _33052_ (.A(_10824_), .B(_10825_), .Y(_00000_[17]));
NAND_g _33053_ (.A(dbg_rs1val[18]), .B(_10790_), .Y(_10826_));
NAND_g _33054_ (.A(_06991_), .B(_10664_), .Y(_10827_));
NAND_g _33055_ (.A(_10826_), .B(_10827_), .Y(_00000_[18]));
NAND_g _33056_ (.A(dbg_rs1val[19]), .B(_10790_), .Y(_10828_));
NAND_g _33057_ (.A(_04805_), .B(_07094_), .Y(_10829_));
NAND_g _33058_ (.A(_10828_), .B(_10829_), .Y(_00000_[19]));
NAND_g _33059_ (.A(dbg_rs1val[20]), .B(_10790_), .Y(_10830_));
NAND_g _33060_ (.A(_07215_), .B(_10664_), .Y(_10831_));
NAND_g _33061_ (.A(_10830_), .B(_10831_), .Y(_00000_[20]));
NAND_g _33062_ (.A(dbg_rs1val[21]), .B(_10790_), .Y(_10832_));
NAND_g _33063_ (.A(_07327_), .B(_10664_), .Y(_10833_));
NAND_g _33064_ (.A(_10832_), .B(_10833_), .Y(_00000_[21]));
NAND_g _33065_ (.A(dbg_rs1val[22]), .B(_10790_), .Y(_10834_));
NAND_g _33066_ (.A(_07429_), .B(_10664_), .Y(_10835_));
NAND_g _33067_ (.A(_10834_), .B(_10835_), .Y(_00000_[22]));
NAND_g _33068_ (.A(dbg_rs1val[23]), .B(_10790_), .Y(_10836_));
NAND_g _33069_ (.A(resetn), .B(_07539_), .Y(_10837_));
NAND_g _33070_ (.A(_10836_), .B(_10837_), .Y(_00000_[23]));
NAND_g _33071_ (.A(dbg_rs1val[24]), .B(_10790_), .Y(_10838_));
NAND_g _33072_ (.A(resetn), .B(_07651_), .Y(_10839_));
NAND_g _33073_ (.A(_10838_), .B(_10839_), .Y(_00000_[24]));
NAND_g _33074_ (.A(dbg_rs1val[25]), .B(_10790_), .Y(_10840_));
NAND_g _33075_ (.A(_07772_), .B(_10664_), .Y(_10841_));
NAND_g _33076_ (.A(_10840_), .B(_10841_), .Y(_00000_[25]));
NAND_g _33077_ (.A(dbg_rs1val[26]), .B(_10790_), .Y(_10842_));
NAND_g _33078_ (.A(resetn), .B(_07877_), .Y(_10843_));
NAND_g _33079_ (.A(_10842_), .B(_10843_), .Y(_00000_[26]));
NAND_g _33080_ (.A(dbg_rs1val[27]), .B(_10790_), .Y(_10844_));
NAND_g _33081_ (.A(_08000_), .B(_10664_), .Y(_10845_));
NAND_g _33082_ (.A(_10844_), .B(_10845_), .Y(_00000_[27]));
NAND_g _33083_ (.A(dbg_rs1val[28]), .B(_10790_), .Y(_10846_));
NAND_g _33084_ (.A(resetn), .B(_08099_), .Y(_10847_));
NAND_g _33085_ (.A(_10846_), .B(_10847_), .Y(_00000_[28]));
NAND_g _33086_ (.A(resetn), .B(_08212_), .Y(_10848_));
NAND_g _33087_ (.A(dbg_rs1val[29]), .B(_10790_), .Y(_10849_));
NAND_g _33088_ (.A(_10848_), .B(_10849_), .Y(_00000_[29]));
NAND_g _33089_ (.A(dbg_rs1val[30]), .B(_10790_), .Y(_10850_));
NAND_g _33090_ (.A(_04805_), .B(_08318_), .Y(_10851_));
NAND_g _33091_ (.A(_10850_), .B(_10851_), .Y(_00000_[30]));
NAND_g _33092_ (.A(dbg_rs1val[31]), .B(_10790_), .Y(_10852_));
NAND_g _33093_ (.A(resetn), .B(_13718_), .Y(_10853_));
NAND_g _33094_ (.A(_10852_), .B(_10853_), .Y(_00000_[31]));
BUF_g _33095_ (.A(cpuregs_0[0]), .Y(_01238_));
BUF_g _33096_ (.A(cpuregs_0[1]), .Y(_01239_));
BUF_g _33097_ (.A(cpuregs_0[2]), .Y(_01240_));
BUF_g _33098_ (.A(cpuregs_0[3]), .Y(_01241_));
BUF_g _33099_ (.A(cpuregs_0[4]), .Y(_01242_));
BUF_g _33100_ (.A(cpuregs_0[5]), .Y(_01243_));
BUF_g _33101_ (.A(cpuregs_0[6]), .Y(_01244_));
BUF_g _33102_ (.A(cpuregs_0[7]), .Y(_01245_));
BUF_g _33103_ (.A(cpuregs_0[8]), .Y(_01246_));
BUF_g _33104_ (.A(cpuregs_0[9]), .Y(_01247_));
BUF_g _33105_ (.A(cpuregs_0[10]), .Y(_01248_));
BUF_g _33106_ (.A(cpuregs_0[11]), .Y(_01249_));
BUF_g _33107_ (.A(cpuregs_0[12]), .Y(_01250_));
BUF_g _33108_ (.A(cpuregs_0[13]), .Y(_01251_));
BUF_g _33109_ (.A(cpuregs_0[14]), .Y(_01252_));
BUF_g _33110_ (.A(cpuregs_0[15]), .Y(_01253_));
BUF_g _33111_ (.A(cpuregs_0[16]), .Y(_01254_));
BUF_g _33112_ (.A(cpuregs_0[17]), .Y(_01255_));
BUF_g _33113_ (.A(cpuregs_0[18]), .Y(_01256_));
BUF_g _33114_ (.A(cpuregs_0[19]), .Y(_01257_));
BUF_g _33115_ (.A(cpuregs_0[20]), .Y(_01258_));
BUF_g _33116_ (.A(cpuregs_0[21]), .Y(_01259_));
BUF_g _33117_ (.A(cpuregs_0[22]), .Y(_01260_));
BUF_g _33118_ (.A(cpuregs_0[23]), .Y(_01261_));
BUF_g _33119_ (.A(cpuregs_0[24]), .Y(_01262_));
BUF_g _33120_ (.A(cpuregs_0[25]), .Y(_01263_));
BUF_g _33121_ (.A(cpuregs_0[26]), .Y(_01264_));
BUF_g _33122_ (.A(cpuregs_0[27]), .Y(_01265_));
BUF_g _33123_ (.A(cpuregs_0[28]), .Y(_01266_));
BUF_g _33124_ (.A(cpuregs_0[29]), .Y(_01267_));
BUF_g _33125_ (.A(cpuregs_0[30]), .Y(_01268_));
BUF_g _33126_ (.A(cpuregs_0[31]), .Y(_01269_));
NAND_g _33127_ (.A(_02964_), .B(_02993_), .Y(dbg_ascii_instr[8]));
NAND_g _33128_ (.A(_02994_), .B(_03011_), .Y(dbg_ascii_instr[9]));
NAND_g _33129_ (.A(_03012_), .B(_03032_), .Y(dbg_ascii_instr[10]));
NAND_g _33130_ (.A(_03033_), .B(_03058_), .Y(dbg_ascii_instr[11]));
NAND_g _33131_ (.A(_03059_), .B(_03085_), .Y(dbg_ascii_instr[12]));
NOR_g _33132_ (.A(_03086_), .B(_03090_), .Y(dbg_ascii_instr[14]));
NAND_g _33133_ (.A(_03091_), .B(_03107_), .Y(dbg_ascii_instr[16]));
NAND_g _33134_ (.A(_03108_), .B(_03128_), .Y(dbg_ascii_instr[17]));
NAND_g _33135_ (.A(_03129_), .B(_03145_), .Y(dbg_ascii_instr[18]));
NAND_g _33136_ (.A(_03146_), .B(_03164_), .Y(dbg_ascii_instr[19]));
NAND_g _33137_ (.A(_03165_), .B(_03178_), .Y(dbg_ascii_instr[20]));
NAND_g _33138_ (.A(_03179_), .B(_03192_), .Y(dbg_ascii_instr[22]));
NAND_g _33139_ (.A(_03193_), .B(_03207_), .Y(dbg_ascii_instr[24]));
NAND_g _33140_ (.A(_03208_), .B(_03223_), .Y(dbg_ascii_instr[25]));
NAND_g _33141_ (.A(_03224_), .B(_03235_), .Y(dbg_ascii_instr[26]));
NAND_g _33142_ (.A(_03236_), .B(_03248_), .Y(dbg_ascii_instr[27]));
NAND_g _33143_ (.A(_03249_), .B(_03265_), .Y(dbg_ascii_instr[28]));
NAND_g _33144_ (.A(_03266_), .B(_03280_), .Y(dbg_ascii_instr[30]));
NAND_g _33145_ (.A(_03281_), .B(_03289_), .Y(dbg_ascii_instr[32]));
NAND_g _33146_ (.A(_03290_), .B(_03299_), .Y(dbg_ascii_instr[33]));
NAND_g _33147_ (.A(_03301_), .B(_03303_), .Y(dbg_ascii_instr[35]));
NAND_g _33148_ (.A(_03304_), .B(_03309_), .Y(dbg_ascii_instr[36]));
NAND_g _33149_ (.A(_03310_), .B(_03314_), .Y(dbg_ascii_instr[38]));
NOR_g _33150_ (.A(_03317_), .B(_03318_), .Y(dbg_ascii_instr[41]));
NAND_g _33151_ (.A(_03321_), .B(_03322_), .Y(dbg_ascii_instr[43]));
NOR_g _33152_ (.A(_03325_), .B(_03326_), .Y(dbg_ascii_instr[52]));
NOR_g _33153_ (.A(_03329_), .B(_03331_), .Y(dbg_ascii_instr[54]));
NOR_g _33154_ (.A(_03334_), .B(_03335_), .Y(dbg_ascii_instr[62]));
NAND_g _33155_ (.A(_08418_), .B(_08419_), .Y(_00018_));
NAND_g _33156_ (.A(_08420_), .B(_08421_), .Y(_00019_));
NAND_g _33157_ (.A(_08422_), .B(_08423_), .Y(_00020_));
NAND_g _33158_ (.A(_08414_), .B(_08415_), .Y(_00021_));
NAND_g _33159_ (.A(_08416_), .B(_08417_), .Y(_00022_));
NAND_g _33160_ (.A(_12476_), .B(_12477_), .Y(_00013_));
NAND_g _33161_ (.A(_12492_), .B(_12493_), .Y(_00014_));
NAND_g _33162_ (.A(_12496_), .B(_12497_), .Y(_00015_));
NAND_g _33163_ (.A(_12480_), .B(_12481_), .Y(_00016_));
NAND_g _33164_ (.A(_08339_), .B(_08340_), .Y(_00017_));
NOR_g _33165_ (.A(_03498_), .B(_03500_), .Y(dbg_insn_rd[0]));
NOR_g _33166_ (.A(_03503_), .B(_03505_), .Y(dbg_insn_rd[1]));
NOR_g _33167_ (.A(_03508_), .B(_03510_), .Y(dbg_insn_rd[2]));
NOR_g _33168_ (.A(_03513_), .B(_03515_), .Y(dbg_insn_rd[3]));
NOR_g _33169_ (.A(_03518_), .B(_03520_), .Y(dbg_insn_rd[4]));
NOR_g _33170_ (.A(_02780_), .B(_02782_), .Y(dbg_insn_rs2[0]));
NOR_g _33171_ (.A(_02785_), .B(_02787_), .Y(dbg_insn_rs2[1]));
NOR_g _33172_ (.A(_02790_), .B(_02792_), .Y(dbg_insn_rs2[2]));
NOR_g _33173_ (.A(_02795_), .B(_02797_), .Y(dbg_insn_rs2[3]));
NOR_g _33174_ (.A(_02800_), .B(_02802_), .Y(dbg_insn_rs2[4]));
NOR_g _33175_ (.A(_03523_), .B(_03525_), .Y(dbg_insn_rs1[0]));
NOR_g _33176_ (.A(_03528_), .B(_03530_), .Y(dbg_insn_rs1[1]));
NOR_g _33177_ (.A(_03533_), .B(_03535_), .Y(dbg_insn_rs1[2]));
NOR_g _33178_ (.A(_03538_), .B(_03540_), .Y(dbg_insn_rs1[3]));
NOR_g _33179_ (.A(_03543_), .B(_03545_), .Y(dbg_insn_rs1[4]));
NOR_g _33180_ (.A(_03338_), .B(_03340_), .Y(dbg_insn_imm[0]));
NOR_g _33181_ (.A(_03343_), .B(_03345_), .Y(dbg_insn_imm[1]));
NOR_g _33182_ (.A(_03348_), .B(_03350_), .Y(dbg_insn_imm[2]));
NOR_g _33183_ (.A(_03353_), .B(_03355_), .Y(dbg_insn_imm[3]));
NOR_g _33184_ (.A(_03358_), .B(_03360_), .Y(dbg_insn_imm[4]));
NOR_g _33185_ (.A(_03363_), .B(_03365_), .Y(dbg_insn_imm[5]));
NOR_g _33186_ (.A(_03368_), .B(_03370_), .Y(dbg_insn_imm[6]));
NOR_g _33187_ (.A(_03373_), .B(_03375_), .Y(dbg_insn_imm[7]));
NOR_g _33188_ (.A(_03378_), .B(_03380_), .Y(dbg_insn_imm[8]));
NOR_g _33189_ (.A(_03383_), .B(_03385_), .Y(dbg_insn_imm[9]));
NOR_g _33190_ (.A(_03388_), .B(_03390_), .Y(dbg_insn_imm[10]));
NOR_g _33191_ (.A(_03393_), .B(_03395_), .Y(dbg_insn_imm[11]));
NOR_g _33192_ (.A(_03398_), .B(_03400_), .Y(dbg_insn_imm[12]));
NOR_g _33193_ (.A(_03403_), .B(_03405_), .Y(dbg_insn_imm[13]));
NOR_g _33194_ (.A(_03408_), .B(_03410_), .Y(dbg_insn_imm[14]));
NOR_g _33195_ (.A(_03413_), .B(_03415_), .Y(dbg_insn_imm[15]));
NOR_g _33196_ (.A(_03418_), .B(_03420_), .Y(dbg_insn_imm[16]));
NOR_g _33197_ (.A(_03423_), .B(_03425_), .Y(dbg_insn_imm[17]));
NOR_g _33198_ (.A(_03428_), .B(_03430_), .Y(dbg_insn_imm[18]));
NOR_g _33199_ (.A(_03433_), .B(_03435_), .Y(dbg_insn_imm[19]));
NOR_g _33200_ (.A(_03438_), .B(_03440_), .Y(dbg_insn_imm[20]));
NOR_g _33201_ (.A(_03443_), .B(_03445_), .Y(dbg_insn_imm[21]));
NOR_g _33202_ (.A(_03448_), .B(_03450_), .Y(dbg_insn_imm[22]));
NOR_g _33203_ (.A(_03453_), .B(_03455_), .Y(dbg_insn_imm[23]));
NOR_g _33204_ (.A(_03458_), .B(_03460_), .Y(dbg_insn_imm[24]));
NOR_g _33205_ (.A(_03463_), .B(_03465_), .Y(dbg_insn_imm[25]));
NOR_g _33206_ (.A(_03468_), .B(_03470_), .Y(dbg_insn_imm[26]));
NOR_g _33207_ (.A(_03473_), .B(_03475_), .Y(dbg_insn_imm[27]));
NOR_g _33208_ (.A(_03478_), .B(_03480_), .Y(dbg_insn_imm[28]));
NOR_g _33209_ (.A(_03483_), .B(_03485_), .Y(dbg_insn_imm[29]));
NOR_g _33210_ (.A(_03488_), .B(_03490_), .Y(dbg_insn_imm[30]));
NOR_g _33211_ (.A(_03493_), .B(_03495_), .Y(dbg_insn_imm[31]));
NAND_g _33212_ (.A(_02815_), .B(_02851_), .Y(dbg_ascii_instr[0]));
NAND_g _33213_ (.A(_02852_), .B(_02887_), .Y(dbg_ascii_instr[1]));
NAND_g _33214_ (.A(_02888_), .B(_02912_), .Y(dbg_ascii_instr[2]));
NAND_g _33215_ (.A(_02913_), .B(_02942_), .Y(dbg_ascii_instr[3]));
NAND_g _33216_ (.A(_02943_), .B(_02963_), .Y(dbg_ascii_instr[4]));
DFFcell _33217_ (.C(clk), .D(_00023_), .Q(cpuregs_29[0]));
DFFcell _33218_ (.C(clk), .D(_00024_), .Q(cpuregs_29[1]));
DFFcell _33219_ (.C(clk), .D(_00025_), .Q(cpuregs_29[2]));
DFFcell _33220_ (.C(clk), .D(_00026_), .Q(cpuregs_29[3]));
DFFcell _33221_ (.C(clk), .D(_00027_), .Q(cpuregs_29[4]));
DFFcell _33222_ (.C(clk), .D(_00028_), .Q(cpuregs_29[5]));
DFFcell _33223_ (.C(clk), .D(_00029_), .Q(cpuregs_29[6]));
DFFcell _33224_ (.C(clk), .D(_00030_), .Q(cpuregs_29[7]));
DFFcell _33225_ (.C(clk), .D(_00031_), .Q(cpuregs_29[8]));
DFFcell _33226_ (.C(clk), .D(_00032_), .Q(cpuregs_29[9]));
DFFcell _33227_ (.C(clk), .D(_00033_), .Q(cpuregs_29[10]));
DFFcell _33228_ (.C(clk), .D(_00034_), .Q(cpuregs_29[11]));
DFFcell _33229_ (.C(clk), .D(_00035_), .Q(cpuregs_29[12]));
DFFcell _33230_ (.C(clk), .D(_00036_), .Q(cpuregs_29[13]));
DFFcell _33231_ (.C(clk), .D(_00037_), .Q(cpuregs_29[14]));
DFFcell _33232_ (.C(clk), .D(_00038_), .Q(cpuregs_29[15]));
DFFcell _33233_ (.C(clk), .D(_00039_), .Q(cpuregs_29[16]));
DFFcell _33234_ (.C(clk), .D(_00040_), .Q(cpuregs_29[17]));
DFFcell _33235_ (.C(clk), .D(_00041_), .Q(cpuregs_29[18]));
DFFcell _33236_ (.C(clk), .D(_00042_), .Q(cpuregs_29[19]));
DFFcell _33237_ (.C(clk), .D(_00043_), .Q(cpuregs_29[20]));
DFFcell _33238_ (.C(clk), .D(_00044_), .Q(cpuregs_29[21]));
DFFcell _33239_ (.C(clk), .D(_00045_), .Q(cpuregs_29[22]));
DFFcell _33240_ (.C(clk), .D(_00046_), .Q(cpuregs_29[23]));
DFFcell _33241_ (.C(clk), .D(_00047_), .Q(cpuregs_29[24]));
DFFcell _33242_ (.C(clk), .D(_00048_), .Q(cpuregs_29[25]));
DFFcell _33243_ (.C(clk), .D(_00049_), .Q(cpuregs_29[26]));
DFFcell _33244_ (.C(clk), .D(_00050_), .Q(cpuregs_29[27]));
DFFcell _33245_ (.C(clk), .D(_00051_), .Q(cpuregs_29[28]));
DFFcell _33246_ (.C(clk), .D(_00052_), .Q(cpuregs_29[29]));
DFFcell _33247_ (.C(clk), .D(_00053_), .Q(cpuregs_29[30]));
DFFcell _33248_ (.C(clk), .D(_00054_), .Q(cpuregs_29[31]));
DFFcell _33249_ (.C(clk), .D(_00055_), .Q(cpuregs_9[0]));
DFFcell _33250_ (.C(clk), .D(_00056_), .Q(cpuregs_9[1]));
DFFcell _33251_ (.C(clk), .D(_00057_), .Q(cpuregs_9[2]));
DFFcell _33252_ (.C(clk), .D(_00058_), .Q(cpuregs_9[3]));
DFFcell _33253_ (.C(clk), .D(_00059_), .Q(cpuregs_9[4]));
DFFcell _33254_ (.C(clk), .D(_00060_), .Q(cpuregs_9[5]));
DFFcell _33255_ (.C(clk), .D(_00061_), .Q(cpuregs_9[6]));
DFFcell _33256_ (.C(clk), .D(_00062_), .Q(cpuregs_9[7]));
DFFcell _33257_ (.C(clk), .D(_00063_), .Q(cpuregs_9[8]));
DFFcell _33258_ (.C(clk), .D(_00064_), .Q(cpuregs_9[9]));
DFFcell _33259_ (.C(clk), .D(_00065_), .Q(cpuregs_9[10]));
DFFcell _33260_ (.C(clk), .D(_00066_), .Q(cpuregs_9[11]));
DFFcell _33261_ (.C(clk), .D(_00067_), .Q(cpuregs_9[12]));
DFFcell _33262_ (.C(clk), .D(_00068_), .Q(cpuregs_9[13]));
DFFcell _33263_ (.C(clk), .D(_00069_), .Q(cpuregs_9[14]));
DFFcell _33264_ (.C(clk), .D(_00070_), .Q(cpuregs_9[15]));
DFFcell _33265_ (.C(clk), .D(_00071_), .Q(cpuregs_9[16]));
DFFcell _33266_ (.C(clk), .D(_00072_), .Q(cpuregs_9[17]));
DFFcell _33267_ (.C(clk), .D(_00073_), .Q(cpuregs_9[18]));
DFFcell _33268_ (.C(clk), .D(_00074_), .Q(cpuregs_9[19]));
DFFcell _33269_ (.C(clk), .D(_00075_), .Q(cpuregs_9[20]));
DFFcell _33270_ (.C(clk), .D(_00076_), .Q(cpuregs_9[21]));
DFFcell _33271_ (.C(clk), .D(_00077_), .Q(cpuregs_9[22]));
DFFcell _33272_ (.C(clk), .D(_00078_), .Q(cpuregs_9[23]));
DFFcell _33273_ (.C(clk), .D(_00079_), .Q(cpuregs_9[24]));
DFFcell _33274_ (.C(clk), .D(_00080_), .Q(cpuregs_9[25]));
DFFcell _33275_ (.C(clk), .D(_00081_), .Q(cpuregs_9[26]));
DFFcell _33276_ (.C(clk), .D(_00082_), .Q(cpuregs_9[27]));
DFFcell _33277_ (.C(clk), .D(_00083_), .Q(cpuregs_9[28]));
DFFcell _33278_ (.C(clk), .D(_00084_), .Q(cpuregs_9[29]));
DFFcell _33279_ (.C(clk), .D(_00085_), .Q(cpuregs_9[30]));
DFFcell _33280_ (.C(clk), .D(_00086_), .Q(cpuregs_9[31]));
DFFcell _33281_ (.C(clk), .D(_00087_), .Q(cpuregs_6[0]));
DFFcell _33282_ (.C(clk), .D(_00088_), .Q(cpuregs_6[1]));
DFFcell _33283_ (.C(clk), .D(_00089_), .Q(cpuregs_6[2]));
DFFcell _33284_ (.C(clk), .D(_00090_), .Q(cpuregs_6[3]));
DFFcell _33285_ (.C(clk), .D(_00091_), .Q(cpuregs_6[4]));
DFFcell _33286_ (.C(clk), .D(_00092_), .Q(cpuregs_6[5]));
DFFcell _33287_ (.C(clk), .D(_00093_), .Q(cpuregs_6[6]));
DFFcell _33288_ (.C(clk), .D(_00094_), .Q(cpuregs_6[7]));
DFFcell _33289_ (.C(clk), .D(_00095_), .Q(cpuregs_6[8]));
DFFcell _33290_ (.C(clk), .D(_00096_), .Q(cpuregs_6[9]));
DFFcell _33291_ (.C(clk), .D(_00097_), .Q(cpuregs_6[10]));
DFFcell _33292_ (.C(clk), .D(_00098_), .Q(cpuregs_6[11]));
DFFcell _33293_ (.C(clk), .D(_00099_), .Q(cpuregs_6[12]));
DFFcell _33294_ (.C(clk), .D(_00100_), .Q(cpuregs_6[13]));
DFFcell _33295_ (.C(clk), .D(_00101_), .Q(cpuregs_6[14]));
DFFcell _33296_ (.C(clk), .D(_00102_), .Q(cpuregs_6[15]));
DFFcell _33297_ (.C(clk), .D(_00103_), .Q(cpuregs_6[16]));
DFFcell _33298_ (.C(clk), .D(_00104_), .Q(cpuregs_6[17]));
DFFcell _33299_ (.C(clk), .D(_00105_), .Q(cpuregs_6[18]));
DFFcell _33300_ (.C(clk), .D(_00106_), .Q(cpuregs_6[19]));
DFFcell _33301_ (.C(clk), .D(_00107_), .Q(cpuregs_6[20]));
DFFcell _33302_ (.C(clk), .D(_00108_), .Q(cpuregs_6[21]));
DFFcell _33303_ (.C(clk), .D(_00109_), .Q(cpuregs_6[22]));
DFFcell _33304_ (.C(clk), .D(_00110_), .Q(cpuregs_6[23]));
DFFcell _33305_ (.C(clk), .D(_00111_), .Q(cpuregs_6[24]));
DFFcell _33306_ (.C(clk), .D(_00112_), .Q(cpuregs_6[25]));
DFFcell _33307_ (.C(clk), .D(_00113_), .Q(cpuregs_6[26]));
DFFcell _33308_ (.C(clk), .D(_00114_), .Q(cpuregs_6[27]));
DFFcell _33309_ (.C(clk), .D(_00115_), .Q(cpuregs_6[28]));
DFFcell _33310_ (.C(clk), .D(_00116_), .Q(cpuregs_6[29]));
DFFcell _33311_ (.C(clk), .D(_00117_), .Q(cpuregs_6[30]));
DFFcell _33312_ (.C(clk), .D(_00118_), .Q(cpuregs_6[31]));
DFFcell _33313_ (.C(clk), .D(_00119_), .Q(cpuregs_18[0]));
DFFcell _33314_ (.C(clk), .D(_00120_), .Q(cpuregs_18[1]));
DFFcell _33315_ (.C(clk), .D(_00121_), .Q(cpuregs_18[2]));
DFFcell _33316_ (.C(clk), .D(_00122_), .Q(cpuregs_18[3]));
DFFcell _33317_ (.C(clk), .D(_00123_), .Q(cpuregs_18[4]));
DFFcell _33318_ (.C(clk), .D(_00124_), .Q(cpuregs_18[5]));
DFFcell _33319_ (.C(clk), .D(_00125_), .Q(cpuregs_18[6]));
DFFcell _33320_ (.C(clk), .D(_00126_), .Q(cpuregs_18[7]));
DFFcell _33321_ (.C(clk), .D(_00127_), .Q(cpuregs_18[8]));
DFFcell _33322_ (.C(clk), .D(_00128_), .Q(cpuregs_18[9]));
DFFcell _33323_ (.C(clk), .D(_00129_), .Q(cpuregs_18[10]));
DFFcell _33324_ (.C(clk), .D(_00130_), .Q(cpuregs_18[11]));
DFFcell _33325_ (.C(clk), .D(_00131_), .Q(cpuregs_18[12]));
DFFcell _33326_ (.C(clk), .D(_00132_), .Q(cpuregs_18[13]));
DFFcell _33327_ (.C(clk), .D(_00133_), .Q(cpuregs_18[14]));
DFFcell _33328_ (.C(clk), .D(_00134_), .Q(cpuregs_18[15]));
DFFcell _33329_ (.C(clk), .D(_00135_), .Q(cpuregs_18[16]));
DFFcell _33330_ (.C(clk), .D(_00136_), .Q(cpuregs_18[17]));
DFFcell _33331_ (.C(clk), .D(_00137_), .Q(cpuregs_18[18]));
DFFcell _33332_ (.C(clk), .D(_00138_), .Q(cpuregs_18[19]));
DFFcell _33333_ (.C(clk), .D(_00139_), .Q(cpuregs_18[20]));
DFFcell _33334_ (.C(clk), .D(_00140_), .Q(cpuregs_18[21]));
DFFcell _33335_ (.C(clk), .D(_00141_), .Q(cpuregs_18[22]));
DFFcell _33336_ (.C(clk), .D(_00142_), .Q(cpuregs_18[23]));
DFFcell _33337_ (.C(clk), .D(_00143_), .Q(cpuregs_18[24]));
DFFcell _33338_ (.C(clk), .D(_00144_), .Q(cpuregs_18[25]));
DFFcell _33339_ (.C(clk), .D(_00145_), .Q(cpuregs_18[26]));
DFFcell _33340_ (.C(clk), .D(_00146_), .Q(cpuregs_18[27]));
DFFcell _33341_ (.C(clk), .D(_00147_), .Q(cpuregs_18[28]));
DFFcell _33342_ (.C(clk), .D(_00148_), .Q(cpuregs_18[29]));
DFFcell _33343_ (.C(clk), .D(_00149_), .Q(cpuregs_18[30]));
DFFcell _33344_ (.C(clk), .D(_00150_), .Q(cpuregs_18[31]));
DFFcell _33345_ (.C(clk), .D(_00151_), .Q(decoded_imm_j[5]));
DFFcell _33346_ (.C(clk), .D(_00152_), .Q(decoded_imm_j[8]));
DFFcell _33347_ (.C(clk), .D(_00153_), .Q(decoded_imm_j[9]));
DFFcell _33348_ (.C(clk), .D(_00154_), .Q(cpuregs_11[0]));
DFFcell _33349_ (.C(clk), .D(_00155_), .Q(cpuregs_11[1]));
DFFcell _33350_ (.C(clk), .D(_00156_), .Q(cpuregs_11[2]));
DFFcell _33351_ (.C(clk), .D(_00157_), .Q(cpuregs_11[3]));
DFFcell _33352_ (.C(clk), .D(_00158_), .Q(cpuregs_11[4]));
DFFcell _33353_ (.C(clk), .D(_00159_), .Q(cpuregs_11[5]));
DFFcell _33354_ (.C(clk), .D(_00160_), .Q(cpuregs_11[6]));
DFFcell _33355_ (.C(clk), .D(_00161_), .Q(cpuregs_11[7]));
DFFcell _33356_ (.C(clk), .D(_00162_), .Q(cpuregs_11[8]));
DFFcell _33357_ (.C(clk), .D(_00163_), .Q(cpuregs_11[9]));
DFFcell _33358_ (.C(clk), .D(_00164_), .Q(cpuregs_11[10]));
DFFcell _33359_ (.C(clk), .D(_00165_), .Q(cpuregs_11[11]));
DFFcell _33360_ (.C(clk), .D(_00166_), .Q(cpuregs_11[12]));
DFFcell _33361_ (.C(clk), .D(_00167_), .Q(cpuregs_11[13]));
DFFcell _33362_ (.C(clk), .D(_00168_), .Q(cpuregs_11[14]));
DFFcell _33363_ (.C(clk), .D(_00169_), .Q(cpuregs_11[15]));
DFFcell _33364_ (.C(clk), .D(_00170_), .Q(cpuregs_11[16]));
DFFcell _33365_ (.C(clk), .D(_00171_), .Q(cpuregs_11[17]));
DFFcell _33366_ (.C(clk), .D(_00172_), .Q(cpuregs_11[18]));
DFFcell _33367_ (.C(clk), .D(_00173_), .Q(cpuregs_11[19]));
DFFcell _33368_ (.C(clk), .D(_00174_), .Q(cpuregs_11[20]));
DFFcell _33369_ (.C(clk), .D(_00175_), .Q(cpuregs_11[21]));
DFFcell _33370_ (.C(clk), .D(_00176_), .Q(cpuregs_11[22]));
DFFcell _33371_ (.C(clk), .D(_00177_), .Q(cpuregs_11[23]));
DFFcell _33372_ (.C(clk), .D(_00178_), .Q(cpuregs_11[24]));
DFFcell _33373_ (.C(clk), .D(_00179_), .Q(cpuregs_11[25]));
DFFcell _33374_ (.C(clk), .D(_00180_), .Q(cpuregs_11[26]));
DFFcell _33375_ (.C(clk), .D(_00181_), .Q(cpuregs_11[27]));
DFFcell _33376_ (.C(clk), .D(_00182_), .Q(cpuregs_11[28]));
DFFcell _33377_ (.C(clk), .D(_00183_), .Q(cpuregs_11[29]));
DFFcell _33378_ (.C(clk), .D(_00184_), .Q(cpuregs_11[30]));
DFFcell _33379_ (.C(clk), .D(_00185_), .Q(cpuregs_11[31]));
DFFcell _33380_ (.C(clk), .D(_00186_), .Q(cpuregs_25[0]));
DFFcell _33381_ (.C(clk), .D(_00187_), .Q(cpuregs_25[1]));
DFFcell _33382_ (.C(clk), .D(_00188_), .Q(cpuregs_25[2]));
DFFcell _33383_ (.C(clk), .D(_00189_), .Q(cpuregs_25[3]));
DFFcell _33384_ (.C(clk), .D(_00190_), .Q(cpuregs_25[4]));
DFFcell _33385_ (.C(clk), .D(_00191_), .Q(cpuregs_25[5]));
DFFcell _33386_ (.C(clk), .D(_00192_), .Q(cpuregs_25[6]));
DFFcell _33387_ (.C(clk), .D(_00193_), .Q(cpuregs_25[7]));
DFFcell _33388_ (.C(clk), .D(_00194_), .Q(cpuregs_25[8]));
DFFcell _33389_ (.C(clk), .D(_00195_), .Q(cpuregs_25[9]));
DFFcell _33390_ (.C(clk), .D(_00196_), .Q(cpuregs_25[10]));
DFFcell _33391_ (.C(clk), .D(_00197_), .Q(cpuregs_25[11]));
DFFcell _33392_ (.C(clk), .D(_00198_), .Q(cpuregs_25[12]));
DFFcell _33393_ (.C(clk), .D(_00199_), .Q(cpuregs_25[13]));
DFFcell _33394_ (.C(clk), .D(_00200_), .Q(cpuregs_25[14]));
DFFcell _33395_ (.C(clk), .D(_00201_), .Q(cpuregs_25[15]));
DFFcell _33396_ (.C(clk), .D(_00202_), .Q(cpuregs_25[16]));
DFFcell _33397_ (.C(clk), .D(_00203_), .Q(cpuregs_25[17]));
DFFcell _33398_ (.C(clk), .D(_00204_), .Q(cpuregs_25[18]));
DFFcell _33399_ (.C(clk), .D(_00205_), .Q(cpuregs_25[19]));
DFFcell _33400_ (.C(clk), .D(_00206_), .Q(cpuregs_25[20]));
DFFcell _33401_ (.C(clk), .D(_00207_), .Q(cpuregs_25[21]));
DFFcell _33402_ (.C(clk), .D(_00208_), .Q(cpuregs_25[22]));
DFFcell _33403_ (.C(clk), .D(_00209_), .Q(cpuregs_25[23]));
DFFcell _33404_ (.C(clk), .D(_00210_), .Q(cpuregs_25[24]));
DFFcell _33405_ (.C(clk), .D(_00211_), .Q(cpuregs_25[25]));
DFFcell _33406_ (.C(clk), .D(_00212_), .Q(cpuregs_25[26]));
DFFcell _33407_ (.C(clk), .D(_00213_), .Q(cpuregs_25[27]));
DFFcell _33408_ (.C(clk), .D(_00214_), .Q(cpuregs_25[28]));
DFFcell _33409_ (.C(clk), .D(_00215_), .Q(cpuregs_25[29]));
DFFcell _33410_ (.C(clk), .D(_00216_), .Q(cpuregs_25[30]));
DFFcell _33411_ (.C(clk), .D(_00217_), .Q(cpuregs_25[31]));
DFFcell _33412_ (.C(clk), .D(_00218_), .Q(cpuregs_4[0]));
DFFcell _33413_ (.C(clk), .D(_00219_), .Q(cpuregs_4[1]));
DFFcell _33414_ (.C(clk), .D(_00220_), .Q(cpuregs_4[2]));
DFFcell _33415_ (.C(clk), .D(_00221_), .Q(cpuregs_4[3]));
DFFcell _33416_ (.C(clk), .D(_00222_), .Q(cpuregs_4[4]));
DFFcell _33417_ (.C(clk), .D(_00223_), .Q(cpuregs_4[5]));
DFFcell _33418_ (.C(clk), .D(_00224_), .Q(cpuregs_4[6]));
DFFcell _33419_ (.C(clk), .D(_00225_), .Q(cpuregs_4[7]));
DFFcell _33420_ (.C(clk), .D(_00226_), .Q(cpuregs_4[8]));
DFFcell _33421_ (.C(clk), .D(_00227_), .Q(cpuregs_4[9]));
DFFcell _33422_ (.C(clk), .D(_00228_), .Q(cpuregs_4[10]));
DFFcell _33423_ (.C(clk), .D(_00229_), .Q(cpuregs_4[11]));
DFFcell _33424_ (.C(clk), .D(_00230_), .Q(cpuregs_4[12]));
DFFcell _33425_ (.C(clk), .D(_00231_), .Q(cpuregs_4[13]));
DFFcell _33426_ (.C(clk), .D(_00232_), .Q(cpuregs_4[14]));
DFFcell _33427_ (.C(clk), .D(_00233_), .Q(cpuregs_4[15]));
DFFcell _33428_ (.C(clk), .D(_00234_), .Q(cpuregs_4[16]));
DFFcell _33429_ (.C(clk), .D(_00235_), .Q(cpuregs_4[17]));
DFFcell _33430_ (.C(clk), .D(_00236_), .Q(cpuregs_4[18]));
DFFcell _33431_ (.C(clk), .D(_00237_), .Q(cpuregs_4[19]));
DFFcell _33432_ (.C(clk), .D(_00238_), .Q(cpuregs_4[20]));
DFFcell _33433_ (.C(clk), .D(_00239_), .Q(cpuregs_4[21]));
DFFcell _33434_ (.C(clk), .D(_00240_), .Q(cpuregs_4[22]));
DFFcell _33435_ (.C(clk), .D(_00241_), .Q(cpuregs_4[23]));
DFFcell _33436_ (.C(clk), .D(_00242_), .Q(cpuregs_4[24]));
DFFcell _33437_ (.C(clk), .D(_00243_), .Q(cpuregs_4[25]));
DFFcell _33438_ (.C(clk), .D(_00244_), .Q(cpuregs_4[26]));
DFFcell _33439_ (.C(clk), .D(_00245_), .Q(cpuregs_4[27]));
DFFcell _33440_ (.C(clk), .D(_00246_), .Q(cpuregs_4[28]));
DFFcell _33441_ (.C(clk), .D(_00247_), .Q(cpuregs_4[29]));
DFFcell _33442_ (.C(clk), .D(_00248_), .Q(cpuregs_4[30]));
DFFcell _33443_ (.C(clk), .D(_00249_), .Q(cpuregs_4[31]));
DFFcell _33444_ (.C(clk), .D(_00018_), .Q(_00012_[0]));
DFFcell _33445_ (.C(clk), .D(_00019_), .Q(_00012_[1]));
DFFcell _33446_ (.C(clk), .D(_00020_), .Q(_00012_[2]));
DFFcell _33447_ (.C(clk), .D(_00021_), .Q(_00012_[3]));
DFFcell _33448_ (.C(clk), .D(_00022_), .Q(_00012_[4]));
DFFcell _33449_ (.C(clk), .D(_00250_), .Q(cpuregs_17[0]));
DFFcell _33450_ (.C(clk), .D(_00251_), .Q(cpuregs_17[1]));
DFFcell _33451_ (.C(clk), .D(_00252_), .Q(cpuregs_17[2]));
DFFcell _33452_ (.C(clk), .D(_00253_), .Q(cpuregs_17[3]));
DFFcell _33453_ (.C(clk), .D(_00254_), .Q(cpuregs_17[4]));
DFFcell _33454_ (.C(clk), .D(_00255_), .Q(cpuregs_17[5]));
DFFcell _33455_ (.C(clk), .D(_00256_), .Q(cpuregs_17[6]));
DFFcell _33456_ (.C(clk), .D(_00257_), .Q(cpuregs_17[7]));
DFFcell _33457_ (.C(clk), .D(_00258_), .Q(cpuregs_17[8]));
DFFcell _33458_ (.C(clk), .D(_00259_), .Q(cpuregs_17[9]));
DFFcell _33459_ (.C(clk), .D(_00260_), .Q(cpuregs_17[10]));
DFFcell _33460_ (.C(clk), .D(_00261_), .Q(cpuregs_17[11]));
DFFcell _33461_ (.C(clk), .D(_00262_), .Q(cpuregs_17[12]));
DFFcell _33462_ (.C(clk), .D(_00263_), .Q(cpuregs_17[13]));
DFFcell _33463_ (.C(clk), .D(_00264_), .Q(cpuregs_17[14]));
DFFcell _33464_ (.C(clk), .D(_00265_), .Q(cpuregs_17[15]));
DFFcell _33465_ (.C(clk), .D(_00266_), .Q(cpuregs_17[16]));
DFFcell _33466_ (.C(clk), .D(_00267_), .Q(cpuregs_17[17]));
DFFcell _33467_ (.C(clk), .D(_00268_), .Q(cpuregs_17[18]));
DFFcell _33468_ (.C(clk), .D(_00269_), .Q(cpuregs_17[19]));
DFFcell _33469_ (.C(clk), .D(_00270_), .Q(cpuregs_17[20]));
DFFcell _33470_ (.C(clk), .D(_00271_), .Q(cpuregs_17[21]));
DFFcell _33471_ (.C(clk), .D(_00272_), .Q(cpuregs_17[22]));
DFFcell _33472_ (.C(clk), .D(_00273_), .Q(cpuregs_17[23]));
DFFcell _33473_ (.C(clk), .D(_00274_), .Q(cpuregs_17[24]));
DFFcell _33474_ (.C(clk), .D(_00275_), .Q(cpuregs_17[25]));
DFFcell _33475_ (.C(clk), .D(_00276_), .Q(cpuregs_17[26]));
DFFcell _33476_ (.C(clk), .D(_00277_), .Q(cpuregs_17[27]));
DFFcell _33477_ (.C(clk), .D(_00278_), .Q(cpuregs_17[28]));
DFFcell _33478_ (.C(clk), .D(_00279_), .Q(cpuregs_17[29]));
DFFcell _33479_ (.C(clk), .D(_00280_), .Q(cpuregs_17[30]));
DFFcell _33480_ (.C(clk), .D(_00281_), .Q(cpuregs_17[31]));
DFFcell _33481_ (.C(clk), .D(_00013_), .Q(_00011_[0]));
DFFcell _33482_ (.C(clk), .D(_00014_), .Q(_00011_[1]));
DFFcell _33483_ (.C(clk), .D(_00015_), .Q(_00011_[2]));
DFFcell _33484_ (.C(clk), .D(_00016_), .Q(_00011_[3]));
DFFcell _33485_ (.C(clk), .D(_00017_), .Q(_00011_[4]));
DFFcell _33486_ (.C(clk), .D(_00282_), .Q(cpuregs_27[0]));
DFFcell _33487_ (.C(clk), .D(_00283_), .Q(cpuregs_27[1]));
DFFcell _33488_ (.C(clk), .D(_00284_), .Q(cpuregs_27[2]));
DFFcell _33489_ (.C(clk), .D(_00285_), .Q(cpuregs_27[3]));
DFFcell _33490_ (.C(clk), .D(_00286_), .Q(cpuregs_27[4]));
DFFcell _33491_ (.C(clk), .D(_00287_), .Q(cpuregs_27[5]));
DFFcell _33492_ (.C(clk), .D(_00288_), .Q(cpuregs_27[6]));
DFFcell _33493_ (.C(clk), .D(_00289_), .Q(cpuregs_27[7]));
DFFcell _33494_ (.C(clk), .D(_00290_), .Q(cpuregs_27[8]));
DFFcell _33495_ (.C(clk), .D(_00291_), .Q(cpuregs_27[9]));
DFFcell _33496_ (.C(clk), .D(_00292_), .Q(cpuregs_27[10]));
DFFcell _33497_ (.C(clk), .D(_00293_), .Q(cpuregs_27[11]));
DFFcell _33498_ (.C(clk), .D(_00294_), .Q(cpuregs_27[12]));
DFFcell _33499_ (.C(clk), .D(_00295_), .Q(cpuregs_27[13]));
DFFcell _33500_ (.C(clk), .D(_00296_), .Q(cpuregs_27[14]));
DFFcell _33501_ (.C(clk), .D(_00297_), .Q(cpuregs_27[15]));
DFFcell _33502_ (.C(clk), .D(_00298_), .Q(cpuregs_27[16]));
DFFcell _33503_ (.C(clk), .D(_00299_), .Q(cpuregs_27[17]));
DFFcell _33504_ (.C(clk), .D(_00300_), .Q(cpuregs_27[18]));
DFFcell _33505_ (.C(clk), .D(_00301_), .Q(cpuregs_27[19]));
DFFcell _33506_ (.C(clk), .D(_00302_), .Q(cpuregs_27[20]));
DFFcell _33507_ (.C(clk), .D(_00303_), .Q(cpuregs_27[21]));
DFFcell _33508_ (.C(clk), .D(_00304_), .Q(cpuregs_27[22]));
DFFcell _33509_ (.C(clk), .D(_00305_), .Q(cpuregs_27[23]));
DFFcell _33510_ (.C(clk), .D(_00306_), .Q(cpuregs_27[24]));
DFFcell _33511_ (.C(clk), .D(_00307_), .Q(cpuregs_27[25]));
DFFcell _33512_ (.C(clk), .D(_00308_), .Q(cpuregs_27[26]));
DFFcell _33513_ (.C(clk), .D(_00309_), .Q(cpuregs_27[27]));
DFFcell _33514_ (.C(clk), .D(_00310_), .Q(cpuregs_27[28]));
DFFcell _33515_ (.C(clk), .D(_00311_), .Q(cpuregs_27[29]));
DFFcell _33516_ (.C(clk), .D(_00312_), .Q(cpuregs_27[30]));
DFFcell _33517_ (.C(clk), .D(_00313_), .Q(cpuregs_27[31]));
DFFcell _33518_ (.C(clk), .D(_00314_), .Q(instr_jalr));
DFFcell _33519_ (.C(clk), .D(_00315_), .Q(instr_auipc));
DFFcell _33520_ (.C(clk), .D(_00316_), .Q(instr_jal));
DFFcell _33521_ (.C(clk), .D(_00317_), .Q(instr_beq));
DFFcell _33522_ (.C(clk), .D(_00318_), .Q(instr_bne));
DFFcell _33523_ (.C(clk), .D(_00319_), .Q(instr_blt));
DFFcell _33524_ (.C(clk), .D(_00320_), .Q(instr_bge));
DFFcell _33525_ (.C(clk), .D(_00321_), .Q(instr_bltu));
DFFcell _33526_ (.C(clk), .D(_00322_), .Q(instr_bgeu));
DFFcell _33527_ (.C(clk), .D(_00323_), .Q(is_sll_srl_sra));
DFFcell _33528_ (.C(clk), .D(_00324_), .Q(instr_lb));
DFFcell _33529_ (.C(clk), .D(_00325_), .Q(instr_lh));
DFFcell _33530_ (.C(clk), .D(_00326_), .Q(instr_lw));
DFFcell _33531_ (.C(clk), .D(_00327_), .Q(instr_lbu));
DFFcell _33532_ (.C(clk), .D(_00328_), .Q(instr_lhu));
DFFcell _33533_ (.C(clk), .D(_00329_), .Q(instr_sb));
DFFcell _33534_ (.C(clk), .D(_00330_), .Q(instr_sh));
DFFcell _33535_ (.C(clk), .D(_00331_), .Q(instr_addi));
DFFcell _33536_ (.C(clk), .D(_00332_), .Q(instr_slti));
DFFcell _33537_ (.C(clk), .D(_00333_), .Q(instr_sltiu));
DFFcell _33538_ (.C(clk), .D(_00334_), .Q(instr_xori));
DFFcell _33539_ (.C(clk), .D(_00335_), .Q(instr_ori));
DFFcell _33540_ (.C(clk), .D(_00336_), .Q(instr_andi));
DFFcell _33541_ (.C(clk), .D(_00337_), .Q(instr_sw));
DFFcell _33542_ (.C(clk), .D(_00338_), .Q(instr_slli));
DFFcell _33543_ (.C(clk), .D(_00339_), .Q(instr_srli));
DFFcell _33544_ (.C(clk), .D(_00340_), .Q(instr_add));
DFFcell _33545_ (.C(clk), .D(_00341_), .Q(instr_sub));
DFFcell _33546_ (.C(clk), .D(_00342_), .Q(instr_sll));
DFFcell _33547_ (.C(clk), .D(_00343_), .Q(instr_slt));
DFFcell _33548_ (.C(clk), .D(_00344_), .Q(instr_sltu));
DFFcell _33549_ (.C(clk), .D(_00345_), .Q(instr_xor));
DFFcell _33550_ (.C(clk), .D(_00346_), .Q(instr_srl));
DFFcell _33551_ (.C(clk), .D(_00347_), .Q(instr_sra));
DFFcell _33552_ (.C(clk), .D(_00348_), .Q(instr_or));
DFFcell _33553_ (.C(clk), .D(_00349_), .Q(instr_and));
DFFcell _33554_ (.C(clk), .D(_00350_), .Q(instr_srai));
DFFcell _33555_ (.C(clk), .D(_00351_), .Q(instr_rdcycle));
DFFcell _33556_ (.C(clk), .D(_00352_), .Q(instr_rdcycleh));
DFFcell _33557_ (.C(clk), .D(_00353_), .Q(instr_rdinstr));
DFFcell _33558_ (.C(clk), .D(_00354_), .Q(instr_rdinstrh));
DFFcell _33559_ (.C(clk), .D(_00355_), .Q(decoded_rd[0]));
DFFcell _33560_ (.C(clk), .D(_00356_), .Q(decoded_rd[1]));
DFFcell _33561_ (.C(clk), .D(_00357_), .Q(decoded_rd[2]));
DFFcell _33562_ (.C(clk), .D(_00358_), .Q(decoded_rd[3]));
DFFcell _33563_ (.C(clk), .D(_00359_), .Q(decoded_rd[4]));
DFFcell _33564_ (.C(clk), .D(_00360_), .Q(decoded_imm_j[11]));
DFFcell _33565_ (.C(clk), .D(_00361_), .Q(decoded_imm_j[3]));
DFFcell _33566_ (.C(clk), .D(_00362_), .Q(decoded_imm[0]));
DFFcell _33567_ (.C(clk), .D(_00363_), .Q(decoded_imm_j[1]));
DFFcell _33568_ (.C(clk), .D(_00364_), .Q(decoded_imm_j[2]));
DFFcell _33569_ (.C(clk), .D(_00006_), .Q(is_lui_auipc_jal));
DFFcell _33570_ (.C(clk), .D(_00365_), .Q(is_lb_lh_lw_lbu_lhu));
DFFcell _33571_ (.C(clk), .D(_00366_), .Q(is_slli_srli_srai));
DFFcell _33572_ (.C(clk), .D(_00367_), .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
DFFcell _33573_ (.C(clk), .D(_00368_), .Q(instr_lui));
DFFcell _33574_ (.C(clk), .D(_00369_), .Q(is_sb_sh_sw));
DFFcell _33575_ (.C(clk), .D(_00007_), .Q(is_slti_blt_slt));
DFFcell _33576_ (.C(clk), .D(_00008_), .Q(is_sltiu_bltu_sltu));
DFFcell _33577_ (.C(clk), .D(_00370_), .Q(is_beq_bne_blt_bge_bltu_bgeu));
DFFcell _33578_ (.C(clk), .D(_00005_), .Q(is_lbu_lhu_lw));
DFFcell _33579_ (.C(clk), .D(_00371_), .Q(is_lui_auipc_jal_jalr_addi_add_sub));
DFFcell _33580_ (.C(clk), .D(_00372_), .Q(is_alu_reg_imm));
DFFcell _33581_ (.C(clk), .D(_00373_), .Q(is_alu_reg_reg));
DFFcell _33582_ (.C(clk), .D(_00374_), .Q(is_compare));
DFFcell _33583_ (.C(clk), .D(_00375_), .Q(mem_do_prefetch));
DFFcell _33584_ (.C(clk), .D(_00376_), .Q(reg_pc[1]));
DFFcell _33585_ (.C(clk), .D(_00377_), .Q(reg_pc[2]));
DFFcell _33586_ (.C(clk), .D(_00378_), .Q(reg_pc[3]));
DFFcell _33587_ (.C(clk), .D(_00379_), .Q(reg_pc[4]));
DFFcell _33588_ (.C(clk), .D(_00380_), .Q(reg_pc[5]));
DFFcell _33589_ (.C(clk), .D(_00381_), .Q(reg_pc[6]));
DFFcell _33590_ (.C(clk), .D(_00382_), .Q(reg_pc[7]));
DFFcell _33591_ (.C(clk), .D(_00383_), .Q(reg_pc[8]));
DFFcell _33592_ (.C(clk), .D(_00384_), .Q(reg_pc[9]));
DFFcell _33593_ (.C(clk), .D(_00385_), .Q(reg_pc[10]));
DFFcell _33594_ (.C(clk), .D(_00386_), .Q(reg_pc[11]));
DFFcell _33595_ (.C(clk), .D(_00387_), .Q(reg_pc[12]));
DFFcell _33596_ (.C(clk), .D(_00388_), .Q(reg_pc[13]));
DFFcell _33597_ (.C(clk), .D(_00389_), .Q(reg_pc[14]));
DFFcell _33598_ (.C(clk), .D(_00390_), .Q(reg_pc[15]));
DFFcell _33599_ (.C(clk), .D(_00391_), .Q(reg_pc[16]));
DFFcell _33600_ (.C(clk), .D(_00392_), .Q(reg_pc[17]));
DFFcell _33601_ (.C(clk), .D(_00393_), .Q(reg_pc[18]));
DFFcell _33602_ (.C(clk), .D(_00394_), .Q(reg_pc[19]));
DFFcell _33603_ (.C(clk), .D(_00395_), .Q(reg_pc[20]));
DFFcell _33604_ (.C(clk), .D(_00396_), .Q(reg_pc[21]));
DFFcell _33605_ (.C(clk), .D(_00397_), .Q(reg_pc[22]));
DFFcell _33606_ (.C(clk), .D(_00398_), .Q(reg_pc[23]));
DFFcell _33607_ (.C(clk), .D(_00399_), .Q(reg_pc[24]));
DFFcell _33608_ (.C(clk), .D(_00400_), .Q(reg_pc[25]));
DFFcell _33609_ (.C(clk), .D(_00401_), .Q(reg_pc[26]));
DFFcell _33610_ (.C(clk), .D(_00402_), .Q(reg_pc[27]));
DFFcell _33611_ (.C(clk), .D(_00403_), .Q(reg_pc[28]));
DFFcell _33612_ (.C(clk), .D(_00404_), .Q(reg_pc[29]));
DFFcell _33613_ (.C(clk), .D(_00405_), .Q(reg_pc[30]));
DFFcell _33614_ (.C(clk), .D(_00406_), .Q(reg_pc[31]));
DFFcell _33615_ (.C(clk), .D(_00407_), .Q(reg_next_pc[1]));
DFFcell _33616_ (.C(clk), .D(_00408_), .Q(reg_next_pc[2]));
DFFcell _33617_ (.C(clk), .D(_00409_), .Q(reg_next_pc[3]));
DFFcell _33618_ (.C(clk), .D(_00410_), .Q(reg_next_pc[4]));
DFFcell _33619_ (.C(clk), .D(_00411_), .Q(reg_next_pc[5]));
DFFcell _33620_ (.C(clk), .D(_00412_), .Q(reg_next_pc[6]));
DFFcell _33621_ (.C(clk), .D(_00413_), .Q(reg_next_pc[7]));
DFFcell _33622_ (.C(clk), .D(_00414_), .Q(reg_next_pc[8]));
DFFcell _33623_ (.C(clk), .D(_00415_), .Q(reg_next_pc[9]));
DFFcell _33624_ (.C(clk), .D(_00416_), .Q(reg_next_pc[10]));
DFFcell _33625_ (.C(clk), .D(_00417_), .Q(reg_next_pc[11]));
DFFcell _33626_ (.C(clk), .D(_00418_), .Q(reg_next_pc[12]));
DFFcell _33627_ (.C(clk), .D(_00419_), .Q(reg_next_pc[13]));
DFFcell _33628_ (.C(clk), .D(_00420_), .Q(reg_next_pc[14]));
DFFcell _33629_ (.C(clk), .D(_00421_), .Q(reg_next_pc[15]));
DFFcell _33630_ (.C(clk), .D(_00422_), .Q(reg_next_pc[16]));
DFFcell _33631_ (.C(clk), .D(_00423_), .Q(reg_next_pc[17]));
DFFcell _33632_ (.C(clk), .D(_00424_), .Q(reg_next_pc[18]));
DFFcell _33633_ (.C(clk), .D(_00425_), .Q(reg_next_pc[19]));
DFFcell _33634_ (.C(clk), .D(_00426_), .Q(reg_next_pc[20]));
DFFcell _33635_ (.C(clk), .D(_00427_), .Q(reg_next_pc[21]));
DFFcell _33636_ (.C(clk), .D(_00428_), .Q(reg_next_pc[22]));
DFFcell _33637_ (.C(clk), .D(_00429_), .Q(reg_next_pc[23]));
DFFcell _33638_ (.C(clk), .D(_00430_), .Q(reg_next_pc[24]));
DFFcell _33639_ (.C(clk), .D(_00431_), .Q(reg_next_pc[25]));
DFFcell _33640_ (.C(clk), .D(_00432_), .Q(reg_next_pc[26]));
DFFcell _33641_ (.C(clk), .D(_00433_), .Q(reg_next_pc[27]));
DFFcell _33642_ (.C(clk), .D(_00434_), .Q(reg_next_pc[28]));
DFFcell _33643_ (.C(clk), .D(_00435_), .Q(reg_next_pc[29]));
DFFcell _33644_ (.C(clk), .D(_00436_), .Q(reg_next_pc[30]));
DFFcell _33645_ (.C(clk), .D(_00437_), .Q(reg_next_pc[31]));
DFFcell _33646_ (.C(clk), .D(_00438_), .Q(count_cycle[0]));
DFFcell _33647_ (.C(clk), .D(_00439_), .Q(count_cycle[1]));
DFFcell _33648_ (.C(clk), .D(_00440_), .Q(count_cycle[2]));
DFFcell _33649_ (.C(clk), .D(_00441_), .Q(count_cycle[3]));
DFFcell _33650_ (.C(clk), .D(_00442_), .Q(count_cycle[4]));
DFFcell _33651_ (.C(clk), .D(_00443_), .Q(count_cycle[5]));
DFFcell _33652_ (.C(clk), .D(_00444_), .Q(count_cycle[6]));
DFFcell _33653_ (.C(clk), .D(_00445_), .Q(count_cycle[7]));
DFFcell _33654_ (.C(clk), .D(_00446_), .Q(count_cycle[8]));
DFFcell _33655_ (.C(clk), .D(_00447_), .Q(count_cycle[9]));
DFFcell _33656_ (.C(clk), .D(_00448_), .Q(count_cycle[10]));
DFFcell _33657_ (.C(clk), .D(_00449_), .Q(count_cycle[11]));
DFFcell _33658_ (.C(clk), .D(_00450_), .Q(count_cycle[12]));
DFFcell _33659_ (.C(clk), .D(_00451_), .Q(count_cycle[13]));
DFFcell _33660_ (.C(clk), .D(_00452_), .Q(count_cycle[14]));
DFFcell _33661_ (.C(clk), .D(_00453_), .Q(count_cycle[15]));
DFFcell _33662_ (.C(clk), .D(_00454_), .Q(count_cycle[16]));
DFFcell _33663_ (.C(clk), .D(_00455_), .Q(count_cycle[17]));
DFFcell _33664_ (.C(clk), .D(_00456_), .Q(count_cycle[18]));
DFFcell _33665_ (.C(clk), .D(_00457_), .Q(count_cycle[19]));
DFFcell _33666_ (.C(clk), .D(_00458_), .Q(count_cycle[20]));
DFFcell _33667_ (.C(clk), .D(_00459_), .Q(count_cycle[21]));
DFFcell _33668_ (.C(clk), .D(_00460_), .Q(count_cycle[22]));
DFFcell _33669_ (.C(clk), .D(_00461_), .Q(count_cycle[23]));
DFFcell _33670_ (.C(clk), .D(_00462_), .Q(count_cycle[24]));
DFFcell _33671_ (.C(clk), .D(_00463_), .Q(count_cycle[25]));
DFFcell _33672_ (.C(clk), .D(_00464_), .Q(count_cycle[26]));
DFFcell _33673_ (.C(clk), .D(_00465_), .Q(count_cycle[27]));
DFFcell _33674_ (.C(clk), .D(_00466_), .Q(count_cycle[28]));
DFFcell _33675_ (.C(clk), .D(_00467_), .Q(count_cycle[29]));
DFFcell _33676_ (.C(clk), .D(_00468_), .Q(count_cycle[30]));
DFFcell _33677_ (.C(clk), .D(_00469_), .Q(count_cycle[31]));
DFFcell _33678_ (.C(clk), .D(_00470_), .Q(count_cycle[32]));
DFFcell _33679_ (.C(clk), .D(_00471_), .Q(count_cycle[33]));
DFFcell _33680_ (.C(clk), .D(_00472_), .Q(count_cycle[34]));
DFFcell _33681_ (.C(clk), .D(_00473_), .Q(count_cycle[35]));
DFFcell _33682_ (.C(clk), .D(_00474_), .Q(count_cycle[36]));
DFFcell _33683_ (.C(clk), .D(_00475_), .Q(count_cycle[37]));
DFFcell _33684_ (.C(clk), .D(_00476_), .Q(count_cycle[38]));
DFFcell _33685_ (.C(clk), .D(_00477_), .Q(count_cycle[39]));
DFFcell _33686_ (.C(clk), .D(_00478_), .Q(count_cycle[40]));
DFFcell _33687_ (.C(clk), .D(_00479_), .Q(count_cycle[41]));
DFFcell _33688_ (.C(clk), .D(_00480_), .Q(count_cycle[42]));
DFFcell _33689_ (.C(clk), .D(_00481_), .Q(count_cycle[43]));
DFFcell _33690_ (.C(clk), .D(_00482_), .Q(count_cycle[44]));
DFFcell _33691_ (.C(clk), .D(_00483_), .Q(count_cycle[45]));
DFFcell _33692_ (.C(clk), .D(_00484_), .Q(count_cycle[46]));
DFFcell _33693_ (.C(clk), .D(_00485_), .Q(count_cycle[47]));
DFFcell _33694_ (.C(clk), .D(_00486_), .Q(count_cycle[48]));
DFFcell _33695_ (.C(clk), .D(_00487_), .Q(count_cycle[49]));
DFFcell _33696_ (.C(clk), .D(_00488_), .Q(count_cycle[50]));
DFFcell _33697_ (.C(clk), .D(_00489_), .Q(count_cycle[51]));
DFFcell _33698_ (.C(clk), .D(_00490_), .Q(count_cycle[52]));
DFFcell _33699_ (.C(clk), .D(_00491_), .Q(count_cycle[53]));
DFFcell _33700_ (.C(clk), .D(_00492_), .Q(count_cycle[54]));
DFFcell _33701_ (.C(clk), .D(_00493_), .Q(count_cycle[55]));
DFFcell _33702_ (.C(clk), .D(_00494_), .Q(count_cycle[56]));
DFFcell _33703_ (.C(clk), .D(_00495_), .Q(count_cycle[57]));
DFFcell _33704_ (.C(clk), .D(_00496_), .Q(count_cycle[58]));
DFFcell _33705_ (.C(clk), .D(_00497_), .Q(count_cycle[59]));
DFFcell _33706_ (.C(clk), .D(_00498_), .Q(count_cycle[60]));
DFFcell _33707_ (.C(clk), .D(_00499_), .Q(count_cycle[61]));
DFFcell _33708_ (.C(clk), .D(_00500_), .Q(count_cycle[62]));
DFFcell _33709_ (.C(clk), .D(_00501_), .Q(count_cycle[63]));
DFFcell _33710_ (.C(clk), .D(_00502_), .Q(pcpi_rs1[31]));
DFFcell _33711_ (.C(clk), .D(_00009_[0]), .Q(reg_out[0]));
DFFcell _33712_ (.C(clk), .D(_00009_[1]), .Q(reg_out[1]));
DFFcell _33713_ (.C(clk), .D(_00009_[2]), .Q(reg_out[2]));
DFFcell _33714_ (.C(clk), .D(_00009_[3]), .Q(reg_out[3]));
DFFcell _33715_ (.C(clk), .D(_00009_[4]), .Q(reg_out[4]));
DFFcell _33716_ (.C(clk), .D(_00009_[5]), .Q(reg_out[5]));
DFFcell _33717_ (.C(clk), .D(_00009_[6]), .Q(reg_out[6]));
DFFcell _33718_ (.C(clk), .D(_00009_[7]), .Q(reg_out[7]));
DFFcell _33719_ (.C(clk), .D(_00009_[8]), .Q(reg_out[8]));
DFFcell _33720_ (.C(clk), .D(_00009_[9]), .Q(reg_out[9]));
DFFcell _33721_ (.C(clk), .D(_00009_[10]), .Q(reg_out[10]));
DFFcell _33722_ (.C(clk), .D(_00009_[11]), .Q(reg_out[11]));
DFFcell _33723_ (.C(clk), .D(_00009_[12]), .Q(reg_out[12]));
DFFcell _33724_ (.C(clk), .D(_00009_[13]), .Q(reg_out[13]));
DFFcell _33725_ (.C(clk), .D(_00009_[14]), .Q(reg_out[14]));
DFFcell _33726_ (.C(clk), .D(_00009_[15]), .Q(reg_out[15]));
DFFcell _33727_ (.C(clk), .D(_00009_[16]), .Q(reg_out[16]));
DFFcell _33728_ (.C(clk), .D(_00009_[17]), .Q(reg_out[17]));
DFFcell _33729_ (.C(clk), .D(_00009_[18]), .Q(reg_out[18]));
DFFcell _33730_ (.C(clk), .D(_00009_[19]), .Q(reg_out[19]));
DFFcell _33731_ (.C(clk), .D(_00009_[20]), .Q(reg_out[20]));
DFFcell _33732_ (.C(clk), .D(_00009_[21]), .Q(reg_out[21]));
DFFcell _33733_ (.C(clk), .D(_00009_[22]), .Q(reg_out[22]));
DFFcell _33734_ (.C(clk), .D(_00009_[23]), .Q(reg_out[23]));
DFFcell _33735_ (.C(clk), .D(_00009_[24]), .Q(reg_out[24]));
DFFcell _33736_ (.C(clk), .D(_00009_[25]), .Q(reg_out[25]));
DFFcell _33737_ (.C(clk), .D(_00009_[26]), .Q(reg_out[26]));
DFFcell _33738_ (.C(clk), .D(_00009_[27]), .Q(reg_out[27]));
DFFcell _33739_ (.C(clk), .D(_00009_[28]), .Q(reg_out[28]));
DFFcell _33740_ (.C(clk), .D(_00009_[29]), .Q(reg_out[29]));
DFFcell _33741_ (.C(clk), .D(_00009_[30]), .Q(reg_out[30]));
DFFcell _33742_ (.C(clk), .D(_00009_[31]), .Q(reg_out[31]));
DFFcell _33743_ (.C(clk), .D(_00010_[0]), .Q(reg_sh[0]));
DFFcell _33744_ (.C(clk), .D(_00010_[1]), .Q(reg_sh[1]));
DFFcell _33745_ (.C(clk), .D(_00010_[2]), .Q(reg_sh[2]));
DFFcell _33746_ (.C(clk), .D(_00010_[3]), .Q(reg_sh[3]));
DFFcell _33747_ (.C(clk), .D(_00010_[4]), .Q(reg_sh[4]));
DFFcell _33748_ (.C(clk), .D(_00503_), .Q(pcpi_rs2[0]));
DFFcell _33749_ (.C(clk), .D(_00504_), .Q(pcpi_rs2[1]));
DFFcell _33750_ (.C(clk), .D(_00505_), .Q(pcpi_rs2[2]));
DFFcell _33751_ (.C(clk), .D(_00506_), .Q(pcpi_rs2[3]));
DFFcell _33752_ (.C(clk), .D(_00507_), .Q(pcpi_rs2[4]));
DFFcell _33753_ (.C(clk), .D(_00508_), .Q(pcpi_rs2[5]));
DFFcell _33754_ (.C(clk), .D(_00509_), .Q(pcpi_rs2[6]));
DFFcell _33755_ (.C(clk), .D(_00510_), .Q(pcpi_rs2[7]));
DFFcell _33756_ (.C(clk), .D(_00511_), .Q(pcpi_rs2[8]));
DFFcell _33757_ (.C(clk), .D(_00512_), .Q(pcpi_rs2[9]));
DFFcell _33758_ (.C(clk), .D(_00513_), .Q(pcpi_rs2[10]));
DFFcell _33759_ (.C(clk), .D(_00514_), .Q(pcpi_rs2[11]));
DFFcell _33760_ (.C(clk), .D(_00515_), .Q(pcpi_rs2[12]));
DFFcell _33761_ (.C(clk), .D(_00516_), .Q(pcpi_rs2[13]));
DFFcell _33762_ (.C(clk), .D(_00517_), .Q(pcpi_rs2[14]));
DFFcell _33763_ (.C(clk), .D(_00518_), .Q(pcpi_rs2[15]));
DFFcell _33764_ (.C(clk), .D(_00519_), .Q(pcpi_rs2[16]));
DFFcell _33765_ (.C(clk), .D(_00520_), .Q(pcpi_rs2[17]));
DFFcell _33766_ (.C(clk), .D(_00521_), .Q(pcpi_rs2[18]));
DFFcell _33767_ (.C(clk), .D(_00522_), .Q(pcpi_rs2[19]));
DFFcell _33768_ (.C(clk), .D(_00523_), .Q(pcpi_rs2[20]));
DFFcell _33769_ (.C(clk), .D(_00524_), .Q(pcpi_rs2[21]));
DFFcell _33770_ (.C(clk), .D(_00525_), .Q(pcpi_rs2[22]));
DFFcell _33771_ (.C(clk), .D(_00526_), .Q(pcpi_rs2[23]));
DFFcell _33772_ (.C(clk), .D(_00527_), .Q(pcpi_rs2[24]));
DFFcell _33773_ (.C(clk), .D(_00528_), .Q(pcpi_rs2[25]));
DFFcell _33774_ (.C(clk), .D(_00529_), .Q(pcpi_rs2[26]));
DFFcell _33775_ (.C(clk), .D(_00530_), .Q(pcpi_rs2[27]));
DFFcell _33776_ (.C(clk), .D(_00531_), .Q(pcpi_rs2[28]));
DFFcell _33777_ (.C(clk), .D(_00532_), .Q(pcpi_rs2[29]));
DFFcell _33778_ (.C(clk), .D(_00533_), .Q(pcpi_rs2[30]));
DFFcell _33779_ (.C(clk), .D(_00534_), .Q(pcpi_rs2[31]));
DFFcell _33780_ (.C(clk), .D(_00535_), .Q(decoder_pseudo_trigger));
DFFcell _33781_ (.C(clk), .D(_00536_), .Q(mem_do_rinst));
DFFcell _33782_ (.C(clk), .D(_00537_), .Q(mem_do_rdata));
DFFcell _33783_ (.C(clk), .D(_00538_), .Q(mem_do_wdata));
DFFcell _33784_ (.C(clk), .D(_00004_), .Q(decoder_trigger));
DFFcell _33785_ (.C(clk), .D(decoder_trigger), .Q(decoder_trigger_q));
DFFcell _33786_ (.C(clk), .D(_00539_), .Q(mem_wordsize[0]));
DFFcell _33787_ (.C(clk), .D(_00540_), .Q(mem_wordsize[1]));
DFFcell _33788_ (.C(clk), .D(decoder_pseudo_trigger), .Q(decoder_pseudo_trigger_q));
DFFcell _33789_ (.C(clk), .D(_00000_[0]), .Q(dbg_rs1val[0]));
DFFcell _33790_ (.C(clk), .D(_00000_[1]), .Q(dbg_rs1val[1]));
DFFcell _33791_ (.C(clk), .D(_00000_[2]), .Q(dbg_rs1val[2]));
DFFcell _33792_ (.C(clk), .D(_00000_[3]), .Q(dbg_rs1val[3]));
DFFcell _33793_ (.C(clk), .D(_00000_[4]), .Q(dbg_rs1val[4]));
DFFcell _33794_ (.C(clk), .D(_00000_[5]), .Q(dbg_rs1val[5]));
DFFcell _33795_ (.C(clk), .D(_00000_[6]), .Q(dbg_rs1val[6]));
DFFcell _33796_ (.C(clk), .D(_00000_[7]), .Q(dbg_rs1val[7]));
DFFcell _33797_ (.C(clk), .D(_00000_[8]), .Q(dbg_rs1val[8]));
DFFcell _33798_ (.C(clk), .D(_00000_[9]), .Q(dbg_rs1val[9]));
DFFcell _33799_ (.C(clk), .D(_00000_[10]), .Q(dbg_rs1val[10]));
DFFcell _33800_ (.C(clk), .D(_00000_[11]), .Q(dbg_rs1val[11]));
DFFcell _33801_ (.C(clk), .D(_00000_[12]), .Q(dbg_rs1val[12]));
DFFcell _33802_ (.C(clk), .D(_00000_[13]), .Q(dbg_rs1val[13]));
DFFcell _33803_ (.C(clk), .D(_00000_[14]), .Q(dbg_rs1val[14]));
DFFcell _33804_ (.C(clk), .D(_00000_[15]), .Q(dbg_rs1val[15]));
DFFcell _33805_ (.C(clk), .D(_00000_[16]), .Q(dbg_rs1val[16]));
DFFcell _33806_ (.C(clk), .D(_00000_[17]), .Q(dbg_rs1val[17]));
DFFcell _33807_ (.C(clk), .D(_00000_[18]), .Q(dbg_rs1val[18]));
DFFcell _33808_ (.C(clk), .D(_00000_[19]), .Q(dbg_rs1val[19]));
DFFcell _33809_ (.C(clk), .D(_00000_[20]), .Q(dbg_rs1val[20]));
DFFcell _33810_ (.C(clk), .D(_00000_[21]), .Q(dbg_rs1val[21]));
DFFcell _33811_ (.C(clk), .D(_00000_[22]), .Q(dbg_rs1val[22]));
DFFcell _33812_ (.C(clk), .D(_00000_[23]), .Q(dbg_rs1val[23]));
DFFcell _33813_ (.C(clk), .D(_00000_[24]), .Q(dbg_rs1val[24]));
DFFcell _33814_ (.C(clk), .D(_00000_[25]), .Q(dbg_rs1val[25]));
DFFcell _33815_ (.C(clk), .D(_00000_[26]), .Q(dbg_rs1val[26]));
DFFcell _33816_ (.C(clk), .D(_00000_[27]), .Q(dbg_rs1val[27]));
DFFcell _33817_ (.C(clk), .D(_00000_[28]), .Q(dbg_rs1val[28]));
DFFcell _33818_ (.C(clk), .D(_00000_[29]), .Q(dbg_rs1val[29]));
DFFcell _33819_ (.C(clk), .D(_00000_[30]), .Q(dbg_rs1val[30]));
DFFcell _33820_ (.C(clk), .D(_00000_[31]), .Q(dbg_rs1val[31]));
DFFcell _33821_ (.C(clk), .D(_00002_[0]), .Q(dbg_rs2val[0]));
DFFcell _33822_ (.C(clk), .D(_00002_[1]), .Q(dbg_rs2val[1]));
DFFcell _33823_ (.C(clk), .D(_00002_[2]), .Q(dbg_rs2val[2]));
DFFcell _33824_ (.C(clk), .D(_00002_[3]), .Q(dbg_rs2val[3]));
DFFcell _33825_ (.C(clk), .D(_00002_[4]), .Q(dbg_rs2val[4]));
DFFcell _33826_ (.C(clk), .D(_00002_[5]), .Q(dbg_rs2val[5]));
DFFcell _33827_ (.C(clk), .D(_00002_[6]), .Q(dbg_rs2val[6]));
DFFcell _33828_ (.C(clk), .D(_00002_[7]), .Q(dbg_rs2val[7]));
DFFcell _33829_ (.C(clk), .D(_00002_[8]), .Q(dbg_rs2val[8]));
DFFcell _33830_ (.C(clk), .D(_00002_[9]), .Q(dbg_rs2val[9]));
DFFcell _33831_ (.C(clk), .D(_00002_[10]), .Q(dbg_rs2val[10]));
DFFcell _33832_ (.C(clk), .D(_00002_[11]), .Q(dbg_rs2val[11]));
DFFcell _33833_ (.C(clk), .D(_00002_[12]), .Q(dbg_rs2val[12]));
DFFcell _33834_ (.C(clk), .D(_00002_[13]), .Q(dbg_rs2val[13]));
DFFcell _33835_ (.C(clk), .D(_00002_[14]), .Q(dbg_rs2val[14]));
DFFcell _33836_ (.C(clk), .D(_00002_[15]), .Q(dbg_rs2val[15]));
DFFcell _33837_ (.C(clk), .D(_00002_[16]), .Q(dbg_rs2val[16]));
DFFcell _33838_ (.C(clk), .D(_00002_[17]), .Q(dbg_rs2val[17]));
DFFcell _33839_ (.C(clk), .D(_00002_[18]), .Q(dbg_rs2val[18]));
DFFcell _33840_ (.C(clk), .D(_00002_[19]), .Q(dbg_rs2val[19]));
DFFcell _33841_ (.C(clk), .D(_00002_[20]), .Q(dbg_rs2val[20]));
DFFcell _33842_ (.C(clk), .D(_00002_[21]), .Q(dbg_rs2val[21]));
DFFcell _33843_ (.C(clk), .D(_00002_[22]), .Q(dbg_rs2val[22]));
DFFcell _33844_ (.C(clk), .D(_00002_[23]), .Q(dbg_rs2val[23]));
DFFcell _33845_ (.C(clk), .D(_00002_[24]), .Q(dbg_rs2val[24]));
DFFcell _33846_ (.C(clk), .D(_00002_[25]), .Q(dbg_rs2val[25]));
DFFcell _33847_ (.C(clk), .D(_00002_[26]), .Q(dbg_rs2val[26]));
DFFcell _33848_ (.C(clk), .D(_00002_[27]), .Q(dbg_rs2val[27]));
DFFcell _33849_ (.C(clk), .D(_00002_[28]), .Q(dbg_rs2val[28]));
DFFcell _33850_ (.C(clk), .D(_00002_[29]), .Q(dbg_rs2val[29]));
DFFcell _33851_ (.C(clk), .D(_00002_[30]), .Q(dbg_rs2val[30]));
DFFcell _33852_ (.C(clk), .D(_00002_[31]), .Q(dbg_rs2val[31]));
DFFcell _33853_ (.C(clk), .D(_00001_), .Q(dbg_rs1val_valid));
DFFcell _33854_ (.C(clk), .D(_00003_), .Q(dbg_rs2val_valid));
DFFcell _33855_ (.C(clk), .D(_00541_), .Q(mem_valid));
DFFcell _33856_ (.C(clk), .D(_00542_), .Q(trap));
DFFcell _33857_ (.C(clk), .D(_00543_), .Q(latched_store));
DFFcell _33858_ (.C(clk), .D(_00544_), .Q(latched_stalu));
DFFcell _33859_ (.C(clk), .D(_00545_), .Q(latched_branch));
DFFcell _33860_ (.C(clk), .D(_00546_), .Q(cpuregs_22[0]));
DFFcell _33861_ (.C(clk), .D(_00547_), .Q(cpuregs_22[1]));
DFFcell _33862_ (.C(clk), .D(_00548_), .Q(cpuregs_22[2]));
DFFcell _33863_ (.C(clk), .D(_00549_), .Q(cpuregs_22[3]));
DFFcell _33864_ (.C(clk), .D(_00550_), .Q(cpuregs_22[4]));
DFFcell _33865_ (.C(clk), .D(_00551_), .Q(cpuregs_22[5]));
DFFcell _33866_ (.C(clk), .D(_00552_), .Q(cpuregs_22[6]));
DFFcell _33867_ (.C(clk), .D(_00553_), .Q(cpuregs_22[7]));
DFFcell _33868_ (.C(clk), .D(_00554_), .Q(cpuregs_22[8]));
DFFcell _33869_ (.C(clk), .D(_00555_), .Q(cpuregs_22[9]));
DFFcell _33870_ (.C(clk), .D(_00556_), .Q(cpuregs_22[10]));
DFFcell _33871_ (.C(clk), .D(_00557_), .Q(cpuregs_22[11]));
DFFcell _33872_ (.C(clk), .D(_00558_), .Q(cpuregs_22[12]));
DFFcell _33873_ (.C(clk), .D(_00559_), .Q(cpuregs_22[13]));
DFFcell _33874_ (.C(clk), .D(_00560_), .Q(cpuregs_22[14]));
DFFcell _33875_ (.C(clk), .D(_00561_), .Q(cpuregs_22[15]));
DFFcell _33876_ (.C(clk), .D(_00562_), .Q(cpuregs_22[16]));
DFFcell _33877_ (.C(clk), .D(_00563_), .Q(cpuregs_22[17]));
DFFcell _33878_ (.C(clk), .D(_00564_), .Q(cpuregs_22[18]));
DFFcell _33879_ (.C(clk), .D(_00565_), .Q(cpuregs_22[19]));
DFFcell _33880_ (.C(clk), .D(_00566_), .Q(cpuregs_22[20]));
DFFcell _33881_ (.C(clk), .D(_00567_), .Q(cpuregs_22[21]));
DFFcell _33882_ (.C(clk), .D(_00568_), .Q(cpuregs_22[22]));
DFFcell _33883_ (.C(clk), .D(_00569_), .Q(cpuregs_22[23]));
DFFcell _33884_ (.C(clk), .D(_00570_), .Q(cpuregs_22[24]));
DFFcell _33885_ (.C(clk), .D(_00571_), .Q(cpuregs_22[25]));
DFFcell _33886_ (.C(clk), .D(_00572_), .Q(cpuregs_22[26]));
DFFcell _33887_ (.C(clk), .D(_00573_), .Q(cpuregs_22[27]));
DFFcell _33888_ (.C(clk), .D(_00574_), .Q(cpuregs_22[28]));
DFFcell _33889_ (.C(clk), .D(_00575_), .Q(cpuregs_22[29]));
DFFcell _33890_ (.C(clk), .D(_00576_), .Q(cpuregs_22[30]));
DFFcell _33891_ (.C(clk), .D(_00577_), .Q(cpuregs_22[31]));
DFFcell _33892_ (.C(clk), .D(_00578_), .Q(cpuregs_21[0]));
DFFcell _33893_ (.C(clk), .D(_00579_), .Q(cpuregs_21[1]));
DFFcell _33894_ (.C(clk), .D(_00580_), .Q(cpuregs_21[2]));
DFFcell _33895_ (.C(clk), .D(_00581_), .Q(cpuregs_21[3]));
DFFcell _33896_ (.C(clk), .D(_00582_), .Q(cpuregs_21[4]));
DFFcell _33897_ (.C(clk), .D(_00583_), .Q(cpuregs_21[5]));
DFFcell _33898_ (.C(clk), .D(_00584_), .Q(cpuregs_21[6]));
DFFcell _33899_ (.C(clk), .D(_00585_), .Q(cpuregs_21[7]));
DFFcell _33900_ (.C(clk), .D(_00586_), .Q(cpuregs_21[8]));
DFFcell _33901_ (.C(clk), .D(_00587_), .Q(cpuregs_21[9]));
DFFcell _33902_ (.C(clk), .D(_00588_), .Q(cpuregs_21[10]));
DFFcell _33903_ (.C(clk), .D(_00589_), .Q(cpuregs_21[11]));
DFFcell _33904_ (.C(clk), .D(_00590_), .Q(cpuregs_21[12]));
DFFcell _33905_ (.C(clk), .D(_00591_), .Q(cpuregs_21[13]));
DFFcell _33906_ (.C(clk), .D(_00592_), .Q(cpuregs_21[14]));
DFFcell _33907_ (.C(clk), .D(_00593_), .Q(cpuregs_21[15]));
DFFcell _33908_ (.C(clk), .D(_00594_), .Q(cpuregs_21[16]));
DFFcell _33909_ (.C(clk), .D(_00595_), .Q(cpuregs_21[17]));
DFFcell _33910_ (.C(clk), .D(_00596_), .Q(cpuregs_21[18]));
DFFcell _33911_ (.C(clk), .D(_00597_), .Q(cpuregs_21[19]));
DFFcell _33912_ (.C(clk), .D(_00598_), .Q(cpuregs_21[20]));
DFFcell _33913_ (.C(clk), .D(_00599_), .Q(cpuregs_21[21]));
DFFcell _33914_ (.C(clk), .D(_00600_), .Q(cpuregs_21[22]));
DFFcell _33915_ (.C(clk), .D(_00601_), .Q(cpuregs_21[23]));
DFFcell _33916_ (.C(clk), .D(_00602_), .Q(cpuregs_21[24]));
DFFcell _33917_ (.C(clk), .D(_00603_), .Q(cpuregs_21[25]));
DFFcell _33918_ (.C(clk), .D(_00604_), .Q(cpuregs_21[26]));
DFFcell _33919_ (.C(clk), .D(_00605_), .Q(cpuregs_21[27]));
DFFcell _33920_ (.C(clk), .D(_00606_), .Q(cpuregs_21[28]));
DFFcell _33921_ (.C(clk), .D(_00607_), .Q(cpuregs_21[29]));
DFFcell _33922_ (.C(clk), .D(_00608_), .Q(cpuregs_21[30]));
DFFcell _33923_ (.C(clk), .D(_00609_), .Q(cpuregs_21[31]));
DFFcell _33924_ (.C(clk), .D(_00610_), .Q(latched_is_lu));
DFFcell _33925_ (.C(clk), .D(_00611_), .Q(latched_is_lh));
DFFcell _33926_ (.C(clk), .D(_00612_), .Q(latched_is_lb));
DFFcell _33927_ (.C(clk), .D(_00613_), .Q(q_insn_rs2[0]));
DFFcell _33928_ (.C(clk), .D(_00614_), .Q(q_insn_rs2[1]));
DFFcell _33929_ (.C(clk), .D(_00615_), .Q(q_insn_rs2[2]));
DFFcell _33930_ (.C(clk), .D(_00616_), .Q(q_insn_rs2[3]));
DFFcell _33931_ (.C(clk), .D(_00617_), .Q(q_insn_rs2[4]));
DFFcell _33932_ (.C(clk), .D(_00618_), .Q(latched_rd[0]));
DFFcell _33933_ (.C(clk), .D(_00619_), .Q(latched_rd[1]));
DFFcell _33934_ (.C(clk), .D(_00620_), .Q(latched_rd[2]));
DFFcell _33935_ (.C(clk), .D(_00621_), .Q(latched_rd[3]));
DFFcell _33936_ (.C(clk), .D(_00622_), .Q(latched_rd[4]));
DFFcell _33937_ (.C(clk), .D(alu_out[0]), .Q(alu_out_q[0]));
DFFcell _33938_ (.C(clk), .D(alu_out[1]), .Q(alu_out_q[1]));
DFFcell _33939_ (.C(clk), .D(alu_out[2]), .Q(alu_out_q[2]));
DFFcell _33940_ (.C(clk), .D(alu_out[3]), .Q(alu_out_q[3]));
DFFcell _33941_ (.C(clk), .D(alu_out[4]), .Q(alu_out_q[4]));
DFFcell _33942_ (.C(clk), .D(alu_out[5]), .Q(alu_out_q[5]));
DFFcell _33943_ (.C(clk), .D(alu_out[6]), .Q(alu_out_q[6]));
DFFcell _33944_ (.C(clk), .D(alu_out[7]), .Q(alu_out_q[7]));
DFFcell _33945_ (.C(clk), .D(alu_out[8]), .Q(alu_out_q[8]));
DFFcell _33946_ (.C(clk), .D(alu_out[9]), .Q(alu_out_q[9]));
DFFcell _33947_ (.C(clk), .D(alu_out[10]), .Q(alu_out_q[10]));
DFFcell _33948_ (.C(clk), .D(alu_out[11]), .Q(alu_out_q[11]));
DFFcell _33949_ (.C(clk), .D(alu_out[12]), .Q(alu_out_q[12]));
DFFcell _33950_ (.C(clk), .D(alu_out[13]), .Q(alu_out_q[13]));
DFFcell _33951_ (.C(clk), .D(alu_out[14]), .Q(alu_out_q[14]));
DFFcell _33952_ (.C(clk), .D(alu_out[15]), .Q(alu_out_q[15]));
DFFcell _33953_ (.C(clk), .D(alu_out[16]), .Q(alu_out_q[16]));
DFFcell _33954_ (.C(clk), .D(alu_out[17]), .Q(alu_out_q[17]));
DFFcell _33955_ (.C(clk), .D(alu_out[18]), .Q(alu_out_q[18]));
DFFcell _33956_ (.C(clk), .D(alu_out[19]), .Q(alu_out_q[19]));
DFFcell _33957_ (.C(clk), .D(alu_out[20]), .Q(alu_out_q[20]));
DFFcell _33958_ (.C(clk), .D(alu_out[21]), .Q(alu_out_q[21]));
DFFcell _33959_ (.C(clk), .D(alu_out[22]), .Q(alu_out_q[22]));
DFFcell _33960_ (.C(clk), .D(alu_out[23]), .Q(alu_out_q[23]));
DFFcell _33961_ (.C(clk), .D(alu_out[24]), .Q(alu_out_q[24]));
DFFcell _33962_ (.C(clk), .D(alu_out[25]), .Q(alu_out_q[25]));
DFFcell _33963_ (.C(clk), .D(alu_out[26]), .Q(alu_out_q[26]));
DFFcell _33964_ (.C(clk), .D(alu_out[27]), .Q(alu_out_q[27]));
DFFcell _33965_ (.C(clk), .D(alu_out[28]), .Q(alu_out_q[28]));
DFFcell _33966_ (.C(clk), .D(alu_out[29]), .Q(alu_out_q[29]));
DFFcell _33967_ (.C(clk), .D(alu_out[30]), .Q(alu_out_q[30]));
DFFcell _33968_ (.C(clk), .D(alu_out[31]), .Q(alu_out_q[31]));
DFFcell _33969_ (.C(clk), .D(_00623_), .Q(q_ascii_instr[0]));
DFFcell _33970_ (.C(clk), .D(_00624_), .Q(q_ascii_instr[1]));
DFFcell _33971_ (.C(clk), .D(_00625_), .Q(q_ascii_instr[2]));
DFFcell _33972_ (.C(clk), .D(_00626_), .Q(q_ascii_instr[3]));
DFFcell _33973_ (.C(clk), .D(_00627_), .Q(q_ascii_instr[4]));
DFFcell _33974_ (.C(clk), .D(_00628_), .Q(q_ascii_instr[8]));
DFFcell _33975_ (.C(clk), .D(_00629_), .Q(q_ascii_instr[9]));
DFFcell _33976_ (.C(clk), .D(_00630_), .Q(q_ascii_instr[10]));
DFFcell _33977_ (.C(clk), .D(_00631_), .Q(q_ascii_instr[11]));
DFFcell _33978_ (.C(clk), .D(_00632_), .Q(q_ascii_instr[12]));
DFFcell _33979_ (.C(clk), .D(_00633_), .Q(q_ascii_instr[14]));
DFFcell _33980_ (.C(clk), .D(_00634_), .Q(q_ascii_instr[16]));
DFFcell _33981_ (.C(clk), .D(_00635_), .Q(q_ascii_instr[17]));
DFFcell _33982_ (.C(clk), .D(_00636_), .Q(q_ascii_instr[18]));
DFFcell _33983_ (.C(clk), .D(_00637_), .Q(q_ascii_instr[19]));
DFFcell _33984_ (.C(clk), .D(_00638_), .Q(q_ascii_instr[20]));
DFFcell _33985_ (.C(clk), .D(_00639_), .Q(q_ascii_instr[22]));
DFFcell _33986_ (.C(clk), .D(_00640_), .Q(q_ascii_instr[24]));
DFFcell _33987_ (.C(clk), .D(_00641_), .Q(q_ascii_instr[25]));
DFFcell _33988_ (.C(clk), .D(_00642_), .Q(q_ascii_instr[26]));
DFFcell _33989_ (.C(clk), .D(_00643_), .Q(q_ascii_instr[27]));
DFFcell _33990_ (.C(clk), .D(_00644_), .Q(q_ascii_instr[28]));
DFFcell _33991_ (.C(clk), .D(_00645_), .Q(q_ascii_instr[30]));
DFFcell _33992_ (.C(clk), .D(_00646_), .Q(q_ascii_instr[32]));
DFFcell _33993_ (.C(clk), .D(_00647_), .Q(q_ascii_instr[33]));
DFFcell _33994_ (.C(clk), .D(_00648_), .Q(q_ascii_instr[35]));
DFFcell _33995_ (.C(clk), .D(_00649_), .Q(q_ascii_instr[36]));
DFFcell _33996_ (.C(clk), .D(_00650_), .Q(q_ascii_instr[38]));
DFFcell _33997_ (.C(clk), .D(_00651_), .Q(q_ascii_instr[41]));
DFFcell _33998_ (.C(clk), .D(_00652_), .Q(q_ascii_instr[43]));
DFFcell _33999_ (.C(clk), .D(_00653_), .Q(q_ascii_instr[52]));
DFFcell _34000_ (.C(clk), .D(_00654_), .Q(q_ascii_instr[54]));
DFFcell _34001_ (.C(clk), .D(_00655_), .Q(q_ascii_instr[62]));
DFFcell _34002_ (.C(clk), .D(_00656_), .Q(q_insn_imm[0]));
DFFcell _34003_ (.C(clk), .D(_00657_), .Q(q_insn_imm[1]));
DFFcell _34004_ (.C(clk), .D(_00658_), .Q(q_insn_imm[2]));
DFFcell _34005_ (.C(clk), .D(_00659_), .Q(q_insn_imm[3]));
DFFcell _34006_ (.C(clk), .D(_00660_), .Q(q_insn_imm[4]));
DFFcell _34007_ (.C(clk), .D(_00661_), .Q(q_insn_imm[5]));
DFFcell _34008_ (.C(clk), .D(_00662_), .Q(q_insn_imm[6]));
DFFcell _34009_ (.C(clk), .D(_00663_), .Q(q_insn_imm[7]));
DFFcell _34010_ (.C(clk), .D(_00664_), .Q(q_insn_imm[8]));
DFFcell _34011_ (.C(clk), .D(_00665_), .Q(q_insn_imm[9]));
DFFcell _34012_ (.C(clk), .D(_00666_), .Q(q_insn_imm[10]));
DFFcell _34013_ (.C(clk), .D(_00667_), .Q(q_insn_imm[11]));
DFFcell _34014_ (.C(clk), .D(_00668_), .Q(q_insn_imm[12]));
DFFcell _34015_ (.C(clk), .D(_00669_), .Q(q_insn_imm[13]));
DFFcell _34016_ (.C(clk), .D(_00670_), .Q(q_insn_imm[14]));
DFFcell _34017_ (.C(clk), .D(_00671_), .Q(q_insn_imm[15]));
DFFcell _34018_ (.C(clk), .D(_00672_), .Q(q_insn_imm[16]));
DFFcell _34019_ (.C(clk), .D(_00673_), .Q(q_insn_imm[17]));
DFFcell _34020_ (.C(clk), .D(_00674_), .Q(q_insn_imm[18]));
DFFcell _34021_ (.C(clk), .D(_00675_), .Q(q_insn_imm[19]));
DFFcell _34022_ (.C(clk), .D(_00676_), .Q(q_insn_imm[20]));
DFFcell _34023_ (.C(clk), .D(_00677_), .Q(q_insn_imm[21]));
DFFcell _34024_ (.C(clk), .D(_00678_), .Q(q_insn_imm[22]));
DFFcell _34025_ (.C(clk), .D(_00679_), .Q(q_insn_imm[23]));
DFFcell _34026_ (.C(clk), .D(_00680_), .Q(q_insn_imm[24]));
DFFcell _34027_ (.C(clk), .D(_00681_), .Q(q_insn_imm[25]));
DFFcell _34028_ (.C(clk), .D(_00682_), .Q(q_insn_imm[26]));
DFFcell _34029_ (.C(clk), .D(_00683_), .Q(q_insn_imm[27]));
DFFcell _34030_ (.C(clk), .D(_00684_), .Q(q_insn_imm[28]));
DFFcell _34031_ (.C(clk), .D(_00685_), .Q(q_insn_imm[29]));
DFFcell _34032_ (.C(clk), .D(_00686_), .Q(q_insn_imm[30]));
DFFcell _34033_ (.C(clk), .D(_00687_), .Q(q_insn_imm[31]));
DFFcell _34034_ (.C(clk), .D(_00688_), .Q(q_insn_rd[0]));
DFFcell _34035_ (.C(clk), .D(_00689_), .Q(q_insn_rd[1]));
DFFcell _34036_ (.C(clk), .D(_00690_), .Q(q_insn_rd[2]));
DFFcell _34037_ (.C(clk), .D(_00691_), .Q(q_insn_rd[3]));
DFFcell _34038_ (.C(clk), .D(_00692_), .Q(q_insn_rd[4]));
DFFcell _34039_ (.C(clk), .D(_00693_), .Q(q_insn_rs1[0]));
DFFcell _34040_ (.C(clk), .D(_00694_), .Q(q_insn_rs1[1]));
DFFcell _34041_ (.C(clk), .D(_00695_), .Q(q_insn_rs1[2]));
DFFcell _34042_ (.C(clk), .D(_00696_), .Q(q_insn_rs1[3]));
DFFcell _34043_ (.C(clk), .D(_00697_), .Q(q_insn_rs1[4]));
DFFcell _34044_ (.C(clk), .D(launch_next_insn), .Q(dbg_next));
DFFcell _34045_ (.C(clk), .D(_00698_), .Q(cached_insn_rd[0]));
DFFcell _34046_ (.C(clk), .D(_00699_), .Q(cached_insn_rd[1]));
DFFcell _34047_ (.C(clk), .D(_00700_), .Q(cached_insn_rd[2]));
DFFcell _34048_ (.C(clk), .D(_00701_), .Q(cached_insn_rd[3]));
DFFcell _34049_ (.C(clk), .D(_00702_), .Q(cached_insn_rd[4]));
DFFcell _34050_ (.C(clk), .D(_00703_), .Q(cached_insn_imm[0]));
DFFcell _34051_ (.C(clk), .D(_00704_), .Q(cached_insn_imm[1]));
DFFcell _34052_ (.C(clk), .D(_00705_), .Q(cached_insn_imm[2]));
DFFcell _34053_ (.C(clk), .D(_00706_), .Q(cached_insn_imm[3]));
DFFcell _34054_ (.C(clk), .D(_00707_), .Q(cached_insn_imm[4]));
DFFcell _34055_ (.C(clk), .D(_00708_), .Q(cached_insn_imm[5]));
DFFcell _34056_ (.C(clk), .D(_00709_), .Q(cached_insn_imm[6]));
DFFcell _34057_ (.C(clk), .D(_00710_), .Q(cached_insn_imm[7]));
DFFcell _34058_ (.C(clk), .D(_00711_), .Q(cached_insn_imm[8]));
DFFcell _34059_ (.C(clk), .D(_00712_), .Q(cached_insn_imm[9]));
DFFcell _34060_ (.C(clk), .D(_00713_), .Q(cached_insn_imm[10]));
DFFcell _34061_ (.C(clk), .D(_00714_), .Q(cached_insn_imm[11]));
DFFcell _34062_ (.C(clk), .D(_00715_), .Q(cached_insn_imm[12]));
DFFcell _34063_ (.C(clk), .D(_00716_), .Q(cached_insn_imm[13]));
DFFcell _34064_ (.C(clk), .D(_00717_), .Q(cached_insn_imm[14]));
DFFcell _34065_ (.C(clk), .D(_00718_), .Q(cached_insn_imm[15]));
DFFcell _34066_ (.C(clk), .D(_00719_), .Q(cached_insn_imm[16]));
DFFcell _34067_ (.C(clk), .D(_00720_), .Q(cached_insn_imm[17]));
DFFcell _34068_ (.C(clk), .D(_00721_), .Q(cached_insn_imm[18]));
DFFcell _34069_ (.C(clk), .D(_00722_), .Q(cached_insn_imm[19]));
DFFcell _34070_ (.C(clk), .D(_00723_), .Q(cached_insn_imm[20]));
DFFcell _34071_ (.C(clk), .D(_00724_), .Q(cached_insn_imm[21]));
DFFcell _34072_ (.C(clk), .D(_00725_), .Q(cached_insn_imm[22]));
DFFcell _34073_ (.C(clk), .D(_00726_), .Q(cached_insn_imm[23]));
DFFcell _34074_ (.C(clk), .D(_00727_), .Q(cached_insn_imm[24]));
DFFcell _34075_ (.C(clk), .D(_00728_), .Q(cached_insn_imm[25]));
DFFcell _34076_ (.C(clk), .D(_00729_), .Q(cached_insn_imm[26]));
DFFcell _34077_ (.C(clk), .D(_00730_), .Q(cached_insn_imm[27]));
DFFcell _34078_ (.C(clk), .D(_00731_), .Q(cached_insn_imm[28]));
DFFcell _34079_ (.C(clk), .D(_00732_), .Q(cached_insn_imm[29]));
DFFcell _34080_ (.C(clk), .D(_00733_), .Q(cached_insn_imm[30]));
DFFcell _34081_ (.C(clk), .D(_00734_), .Q(cached_insn_imm[31]));
DFFcell _34082_ (.C(clk), .D(_00735_), .Q(cached_insn_rs1[0]));
DFFcell _34083_ (.C(clk), .D(_00736_), .Q(cached_insn_rs1[1]));
DFFcell _34084_ (.C(clk), .D(_00737_), .Q(cached_insn_rs1[2]));
DFFcell _34085_ (.C(clk), .D(_00738_), .Q(cached_insn_rs1[3]));
DFFcell _34086_ (.C(clk), .D(_00739_), .Q(cached_insn_rs1[4]));
DFFcell _34087_ (.C(clk), .D(_00740_), .Q(cached_insn_rs2[0]));
DFFcell _34088_ (.C(clk), .D(_00741_), .Q(cached_insn_rs2[1]));
DFFcell _34089_ (.C(clk), .D(_00742_), .Q(cached_insn_rs2[2]));
DFFcell _34090_ (.C(clk), .D(_00743_), .Q(cached_insn_rs2[3]));
DFFcell _34091_ (.C(clk), .D(_00744_), .Q(cached_insn_rs2[4]));
DFFcell _34092_ (.C(clk), .D(_00745_), .Q(cached_ascii_instr[0]));
DFFcell _34093_ (.C(clk), .D(_00746_), .Q(cached_ascii_instr[1]));
DFFcell _34094_ (.C(clk), .D(_00747_), .Q(cached_ascii_instr[2]));
DFFcell _34095_ (.C(clk), .D(_00748_), .Q(cached_ascii_instr[3]));
DFFcell _34096_ (.C(clk), .D(_00749_), .Q(cached_ascii_instr[4]));
DFFcell _34097_ (.C(clk), .D(_00750_), .Q(cached_ascii_instr[8]));
DFFcell _34098_ (.C(clk), .D(_00751_), .Q(cached_ascii_instr[9]));
DFFcell _34099_ (.C(clk), .D(_00752_), .Q(cached_ascii_instr[10]));
DFFcell _34100_ (.C(clk), .D(_00753_), .Q(cached_ascii_instr[11]));
DFFcell _34101_ (.C(clk), .D(_00754_), .Q(cached_ascii_instr[12]));
DFFcell _34102_ (.C(clk), .D(_00755_), .Q(cached_ascii_instr[14]));
DFFcell _34103_ (.C(clk), .D(_00756_), .Q(cached_ascii_instr[16]));
DFFcell _34104_ (.C(clk), .D(_00757_), .Q(cached_ascii_instr[17]));
DFFcell _34105_ (.C(clk), .D(_00758_), .Q(cached_ascii_instr[18]));
DFFcell _34106_ (.C(clk), .D(_00759_), .Q(cached_ascii_instr[19]));
DFFcell _34107_ (.C(clk), .D(_00760_), .Q(cached_ascii_instr[20]));
DFFcell _34108_ (.C(clk), .D(_00761_), .Q(cached_ascii_instr[22]));
DFFcell _34109_ (.C(clk), .D(_00762_), .Q(cached_ascii_instr[24]));
DFFcell _34110_ (.C(clk), .D(_00763_), .Q(cached_ascii_instr[25]));
DFFcell _34111_ (.C(clk), .D(_00764_), .Q(cached_ascii_instr[26]));
DFFcell _34112_ (.C(clk), .D(_00765_), .Q(cached_ascii_instr[27]));
DFFcell _34113_ (.C(clk), .D(_00766_), .Q(cached_ascii_instr[28]));
DFFcell _34114_ (.C(clk), .D(_00767_), .Q(cached_ascii_instr[30]));
DFFcell _34115_ (.C(clk), .D(_00768_), .Q(cached_ascii_instr[32]));
DFFcell _34116_ (.C(clk), .D(_00769_), .Q(cached_ascii_instr[33]));
DFFcell _34117_ (.C(clk), .D(_00770_), .Q(cached_ascii_instr[35]));
DFFcell _34118_ (.C(clk), .D(_00771_), .Q(cached_ascii_instr[36]));
DFFcell _34119_ (.C(clk), .D(_00772_), .Q(cached_ascii_instr[38]));
DFFcell _34120_ (.C(clk), .D(_00773_), .Q(cached_ascii_instr[41]));
DFFcell _34121_ (.C(clk), .D(_00774_), .Q(cached_ascii_instr[43]));
DFFcell _34122_ (.C(clk), .D(_00775_), .Q(cached_ascii_instr[52]));
DFFcell _34123_ (.C(clk), .D(_00776_), .Q(cached_ascii_instr[54]));
DFFcell _34124_ (.C(clk), .D(_00777_), .Q(cached_ascii_instr[62]));
DFFcell _34125_ (.C(clk), .D(_00778_), .Q(mem_instr));
DFFcell _34126_ (.C(clk), .D(_00779_), .Q(mem_rdata_q[7]));
DFFcell _34127_ (.C(clk), .D(_00780_), .Q(mem_rdata_q[8]));
DFFcell _34128_ (.C(clk), .D(_00781_), .Q(mem_rdata_q[9]));
DFFcell _34129_ (.C(clk), .D(_00782_), .Q(mem_rdata_q[10]));
DFFcell _34130_ (.C(clk), .D(_00783_), .Q(mem_rdata_q[11]));
DFFcell _34131_ (.C(clk), .D(_00784_), .Q(mem_rdata_q[12]));
DFFcell _34132_ (.C(clk), .D(_00785_), .Q(mem_rdata_q[13]));
DFFcell _34133_ (.C(clk), .D(_00786_), .Q(mem_rdata_q[14]));
DFFcell _34134_ (.C(clk), .D(_00787_), .Q(mem_rdata_q[15]));
DFFcell _34135_ (.C(clk), .D(_00788_), .Q(mem_rdata_q[16]));
DFFcell _34136_ (.C(clk), .D(_00789_), .Q(mem_rdata_q[17]));
DFFcell _34137_ (.C(clk), .D(_00790_), .Q(mem_rdata_q[18]));
DFFcell _34138_ (.C(clk), .D(_00791_), .Q(mem_rdata_q[19]));
DFFcell _34139_ (.C(clk), .D(_00792_), .Q(mem_rdata_q[20]));
DFFcell _34140_ (.C(clk), .D(_00793_), .Q(mem_rdata_q[21]));
DFFcell _34141_ (.C(clk), .D(_00794_), .Q(mem_rdata_q[22]));
DFFcell _34142_ (.C(clk), .D(_00795_), .Q(mem_rdata_q[23]));
DFFcell _34143_ (.C(clk), .D(_00796_), .Q(mem_rdata_q[24]));
DFFcell _34144_ (.C(clk), .D(_00797_), .Q(mem_rdata_q[25]));
DFFcell _34145_ (.C(clk), .D(_00798_), .Q(mem_rdata_q[26]));
DFFcell _34146_ (.C(clk), .D(_00799_), .Q(mem_rdata_q[27]));
DFFcell _34147_ (.C(clk), .D(_00800_), .Q(mem_rdata_q[28]));
DFFcell _34148_ (.C(clk), .D(_00801_), .Q(mem_rdata_q[29]));
DFFcell _34149_ (.C(clk), .D(_00802_), .Q(mem_rdata_q[30]));
DFFcell _34150_ (.C(clk), .D(_00803_), .Q(mem_rdata_q[31]));
DFFcell _34151_ (.C(clk), .D(_00804_), .Q(mem_addr[2]));
DFFcell _34152_ (.C(clk), .D(_00805_), .Q(mem_addr[3]));
DFFcell _34153_ (.C(clk), .D(_00806_), .Q(mem_addr[4]));
DFFcell _34154_ (.C(clk), .D(_00807_), .Q(mem_addr[5]));
DFFcell _34155_ (.C(clk), .D(_00808_), .Q(mem_addr[6]));
DFFcell _34156_ (.C(clk), .D(_00809_), .Q(mem_addr[7]));
DFFcell _34157_ (.C(clk), .D(_00810_), .Q(mem_addr[8]));
DFFcell _34158_ (.C(clk), .D(_00811_), .Q(mem_addr[9]));
DFFcell _34159_ (.C(clk), .D(_00812_), .Q(mem_addr[10]));
DFFcell _34160_ (.C(clk), .D(_00813_), .Q(mem_addr[11]));
DFFcell _34161_ (.C(clk), .D(_00814_), .Q(mem_addr[12]));
DFFcell _34162_ (.C(clk), .D(_00815_), .Q(mem_addr[13]));
DFFcell _34163_ (.C(clk), .D(_00816_), .Q(mem_addr[14]));
DFFcell _34164_ (.C(clk), .D(_00817_), .Q(mem_addr[15]));
DFFcell _34165_ (.C(clk), .D(_00818_), .Q(mem_addr[16]));
DFFcell _34166_ (.C(clk), .D(_00819_), .Q(mem_addr[17]));
DFFcell _34167_ (.C(clk), .D(_00820_), .Q(mem_addr[18]));
DFFcell _34168_ (.C(clk), .D(_00821_), .Q(mem_addr[19]));
DFFcell _34169_ (.C(clk), .D(_00822_), .Q(mem_addr[20]));
DFFcell _34170_ (.C(clk), .D(_00823_), .Q(mem_addr[21]));
DFFcell _34171_ (.C(clk), .D(_00824_), .Q(mem_addr[22]));
DFFcell _34172_ (.C(clk), .D(_00825_), .Q(mem_addr[23]));
DFFcell _34173_ (.C(clk), .D(_00826_), .Q(mem_addr[24]));
DFFcell _34174_ (.C(clk), .D(_00827_), .Q(mem_addr[25]));
DFFcell _34175_ (.C(clk), .D(_00828_), .Q(mem_addr[26]));
DFFcell _34176_ (.C(clk), .D(_00829_), .Q(mem_addr[27]));
DFFcell _34177_ (.C(clk), .D(_00830_), .Q(mem_addr[28]));
DFFcell _34178_ (.C(clk), .D(_00831_), .Q(mem_addr[29]));
DFFcell _34179_ (.C(clk), .D(_00832_), .Q(mem_addr[30]));
DFFcell _34180_ (.C(clk), .D(_00833_), .Q(mem_addr[31]));
DFFcell _34181_ (.C(clk), .D(_00834_), .Q(mem_wdata[0]));
DFFcell _34182_ (.C(clk), .D(_00835_), .Q(mem_wdata[1]));
DFFcell _34183_ (.C(clk), .D(_00836_), .Q(mem_wdata[2]));
DFFcell _34184_ (.C(clk), .D(_00837_), .Q(mem_wdata[3]));
DFFcell _34185_ (.C(clk), .D(_00838_), .Q(mem_wdata[4]));
DFFcell _34186_ (.C(clk), .D(_00839_), .Q(mem_wdata[5]));
DFFcell _34187_ (.C(clk), .D(_00840_), .Q(mem_wdata[6]));
DFFcell _34188_ (.C(clk), .D(_00841_), .Q(mem_wdata[7]));
DFFcell _34189_ (.C(clk), .D(_00842_), .Q(mem_wdata[8]));
DFFcell _34190_ (.C(clk), .D(_00843_), .Q(mem_wdata[9]));
DFFcell _34191_ (.C(clk), .D(_00844_), .Q(mem_wdata[10]));
DFFcell _34192_ (.C(clk), .D(_00845_), .Q(mem_wdata[11]));
DFFcell _34193_ (.C(clk), .D(_00846_), .Q(mem_wdata[12]));
DFFcell _34194_ (.C(clk), .D(_00847_), .Q(mem_wdata[13]));
DFFcell _34195_ (.C(clk), .D(_00848_), .Q(mem_wdata[14]));
DFFcell _34196_ (.C(clk), .D(_00849_), .Q(mem_wdata[15]));
DFFcell _34197_ (.C(clk), .D(_00850_), .Q(mem_wdata[16]));
DFFcell _34198_ (.C(clk), .D(_00851_), .Q(mem_wdata[17]));
DFFcell _34199_ (.C(clk), .D(_00852_), .Q(mem_wdata[18]));
DFFcell _34200_ (.C(clk), .D(_00853_), .Q(mem_wdata[19]));
DFFcell _34201_ (.C(clk), .D(_00854_), .Q(mem_wdata[20]));
DFFcell _34202_ (.C(clk), .D(_00855_), .Q(mem_wdata[21]));
DFFcell _34203_ (.C(clk), .D(_00856_), .Q(mem_wdata[22]));
DFFcell _34204_ (.C(clk), .D(_00857_), .Q(mem_wdata[23]));
DFFcell _34205_ (.C(clk), .D(_00858_), .Q(mem_wdata[24]));
DFFcell _34206_ (.C(clk), .D(_00859_), .Q(mem_wdata[25]));
DFFcell _34207_ (.C(clk), .D(_00860_), .Q(mem_wdata[26]));
DFFcell _34208_ (.C(clk), .D(_00861_), .Q(mem_wdata[27]));
DFFcell _34209_ (.C(clk), .D(_00862_), .Q(mem_wdata[28]));
DFFcell _34210_ (.C(clk), .D(_00863_), .Q(mem_wdata[29]));
DFFcell _34211_ (.C(clk), .D(_00864_), .Q(mem_wdata[30]));
DFFcell _34212_ (.C(clk), .D(_00865_), .Q(mem_wdata[31]));
DFFcell _34213_ (.C(clk), .D(_00866_), .Q(mem_wstrb[0]));
DFFcell _34214_ (.C(clk), .D(_00867_), .Q(mem_wstrb[1]));
DFFcell _34215_ (.C(clk), .D(_00868_), .Q(mem_wstrb[2]));
DFFcell _34216_ (.C(clk), .D(_00869_), .Q(mem_wstrb[3]));
DFFcell _34217_ (.C(clk), .D(_00870_), .Q(mem_state[0]));
DFFcell _34218_ (.C(clk), .D(_00871_), .Q(mem_state[1]));
DFFcell _34219_ (.C(clk), .D(_00872_), .Q(mem_rdata_q[0]));
DFFcell _34220_ (.C(clk), .D(_00873_), .Q(mem_rdata_q[1]));
DFFcell _34221_ (.C(clk), .D(_00874_), .Q(mem_rdata_q[2]));
DFFcell _34222_ (.C(clk), .D(_00875_), .Q(mem_rdata_q[3]));
DFFcell _34223_ (.C(clk), .D(_00876_), .Q(mem_rdata_q[4]));
DFFcell _34224_ (.C(clk), .D(_00877_), .Q(mem_rdata_q[5]));
DFFcell _34225_ (.C(clk), .D(_00878_), .Q(mem_rdata_q[6]));
DFFcell _34226_ (.C(clk), .D(_00879_), .Q(reg_next_pc[0]));
DFFcell _34227_ (.C(clk), .D(_00880_), .Q(decoded_imm[31]));
DFFcell _34228_ (.C(clk), .D(_00881_), .Q(decoded_imm[30]));
DFFcell _34229_ (.C(clk), .D(_00882_), .Q(decoded_imm[29]));
DFFcell _34230_ (.C(clk), .D(_00883_), .Q(decoded_imm[28]));
DFFcell _34231_ (.C(clk), .D(_00884_), .Q(decoded_imm[27]));
DFFcell _34232_ (.C(clk), .D(_00885_), .Q(decoded_imm[26]));
DFFcell _34233_ (.C(clk), .D(_00886_), .Q(decoded_imm[25]));
DFFcell _34234_ (.C(clk), .D(_00887_), .Q(decoded_imm[24]));
DFFcell _34235_ (.C(clk), .D(_00888_), .Q(decoded_imm[23]));
DFFcell _34236_ (.C(clk), .D(_00889_), .Q(decoded_imm[22]));
DFFcell _34237_ (.C(clk), .D(_00890_), .Q(decoded_imm[21]));
DFFcell _34238_ (.C(clk), .D(_00891_), .Q(decoded_imm[20]));
DFFcell _34239_ (.C(clk), .D(_00892_), .Q(decoded_imm[19]));
DFFcell _34240_ (.C(clk), .D(_00893_), .Q(decoded_imm[18]));
DFFcell _34241_ (.C(clk), .D(_00894_), .Q(decoded_imm[17]));
DFFcell _34242_ (.C(clk), .D(_00895_), .Q(decoded_imm[16]));
DFFcell _34243_ (.C(clk), .D(_00896_), .Q(decoded_imm[15]));
DFFcell _34244_ (.C(clk), .D(_00897_), .Q(decoded_imm[14]));
DFFcell _34245_ (.C(clk), .D(_00898_), .Q(decoded_imm[13]));
DFFcell _34246_ (.C(clk), .D(_00899_), .Q(decoded_imm[12]));
DFFcell _34247_ (.C(clk), .D(_00900_), .Q(decoded_imm[11]));
DFFcell _34248_ (.C(clk), .D(_00901_), .Q(decoded_imm[10]));
DFFcell _34249_ (.C(clk), .D(_00902_), .Q(decoded_imm[9]));
DFFcell _34250_ (.C(clk), .D(_00903_), .Q(decoded_imm[8]));
DFFcell _34251_ (.C(clk), .D(_00904_), .Q(decoded_imm[7]));
DFFcell _34252_ (.C(clk), .D(_00905_), .Q(decoded_imm[6]));
DFFcell _34253_ (.C(clk), .D(_00906_), .Q(decoded_imm[5]));
DFFcell _34254_ (.C(clk), .D(_00907_), .Q(decoded_imm[4]));
DFFcell _34255_ (.C(clk), .D(_00908_), .Q(decoded_imm[3]));
DFFcell _34256_ (.C(clk), .D(_00909_), .Q(decoded_imm[2]));
DFFcell _34257_ (.C(clk), .D(_00910_), .Q(decoded_imm[1]));
DFFcell _34258_ (.C(clk), .D(_00911_), .Q(cpuregs_31[0]));
DFFcell _34259_ (.C(clk), .D(_00912_), .Q(cpuregs_31[1]));
DFFcell _34260_ (.C(clk), .D(_00913_), .Q(cpuregs_31[2]));
DFFcell _34261_ (.C(clk), .D(_00914_), .Q(cpuregs_31[3]));
DFFcell _34262_ (.C(clk), .D(_00915_), .Q(cpuregs_31[4]));
DFFcell _34263_ (.C(clk), .D(_00916_), .Q(cpuregs_31[5]));
DFFcell _34264_ (.C(clk), .D(_00917_), .Q(cpuregs_31[6]));
DFFcell _34265_ (.C(clk), .D(_00918_), .Q(cpuregs_31[7]));
DFFcell _34266_ (.C(clk), .D(_00919_), .Q(cpuregs_31[8]));
DFFcell _34267_ (.C(clk), .D(_00920_), .Q(cpuregs_31[9]));
DFFcell _34268_ (.C(clk), .D(_00921_), .Q(cpuregs_31[10]));
DFFcell _34269_ (.C(clk), .D(_00922_), .Q(cpuregs_31[11]));
DFFcell _34270_ (.C(clk), .D(_00923_), .Q(cpuregs_31[12]));
DFFcell _34271_ (.C(clk), .D(_00924_), .Q(cpuregs_31[13]));
DFFcell _34272_ (.C(clk), .D(_00925_), .Q(cpuregs_31[14]));
DFFcell _34273_ (.C(clk), .D(_00926_), .Q(cpuregs_31[15]));
DFFcell _34274_ (.C(clk), .D(_00927_), .Q(cpuregs_31[16]));
DFFcell _34275_ (.C(clk), .D(_00928_), .Q(cpuregs_31[17]));
DFFcell _34276_ (.C(clk), .D(_00929_), .Q(cpuregs_31[18]));
DFFcell _34277_ (.C(clk), .D(_00930_), .Q(cpuregs_31[19]));
DFFcell _34278_ (.C(clk), .D(_00931_), .Q(cpuregs_31[20]));
DFFcell _34279_ (.C(clk), .D(_00932_), .Q(cpuregs_31[21]));
DFFcell _34280_ (.C(clk), .D(_00933_), .Q(cpuregs_31[22]));
DFFcell _34281_ (.C(clk), .D(_00934_), .Q(cpuregs_31[23]));
DFFcell _34282_ (.C(clk), .D(_00935_), .Q(cpuregs_31[24]));
DFFcell _34283_ (.C(clk), .D(_00936_), .Q(cpuregs_31[25]));
DFFcell _34284_ (.C(clk), .D(_00937_), .Q(cpuregs_31[26]));
DFFcell _34285_ (.C(clk), .D(_00938_), .Q(cpuregs_31[27]));
DFFcell _34286_ (.C(clk), .D(_00939_), .Q(cpuregs_31[28]));
DFFcell _34287_ (.C(clk), .D(_00940_), .Q(cpuregs_31[29]));
DFFcell _34288_ (.C(clk), .D(_00941_), .Q(cpuregs_31[30]));
DFFcell _34289_ (.C(clk), .D(_00942_), .Q(cpuregs_31[31]));
DFFcell _34290_ (.C(clk), .D(_00943_), .Q(cpuregs_3[0]));
DFFcell _34291_ (.C(clk), .D(_00944_), .Q(cpuregs_3[1]));
DFFcell _34292_ (.C(clk), .D(_00945_), .Q(cpuregs_3[2]));
DFFcell _34293_ (.C(clk), .D(_00946_), .Q(cpuregs_3[3]));
DFFcell _34294_ (.C(clk), .D(_00947_), .Q(cpuregs_3[4]));
DFFcell _34295_ (.C(clk), .D(_00948_), .Q(cpuregs_3[5]));
DFFcell _34296_ (.C(clk), .D(_00949_), .Q(cpuregs_3[6]));
DFFcell _34297_ (.C(clk), .D(_00950_), .Q(cpuregs_3[7]));
DFFcell _34298_ (.C(clk), .D(_00951_), .Q(cpuregs_3[8]));
DFFcell _34299_ (.C(clk), .D(_00952_), .Q(cpuregs_3[9]));
DFFcell _34300_ (.C(clk), .D(_00953_), .Q(cpuregs_3[10]));
DFFcell _34301_ (.C(clk), .D(_00954_), .Q(cpuregs_3[11]));
DFFcell _34302_ (.C(clk), .D(_00955_), .Q(cpuregs_3[12]));
DFFcell _34303_ (.C(clk), .D(_00956_), .Q(cpuregs_3[13]));
DFFcell _34304_ (.C(clk), .D(_00957_), .Q(cpuregs_3[14]));
DFFcell _34305_ (.C(clk), .D(_00958_), .Q(cpuregs_3[15]));
DFFcell _34306_ (.C(clk), .D(_00959_), .Q(cpuregs_3[16]));
DFFcell _34307_ (.C(clk), .D(_00960_), .Q(cpuregs_3[17]));
DFFcell _34308_ (.C(clk), .D(_00961_), .Q(cpuregs_3[18]));
DFFcell _34309_ (.C(clk), .D(_00962_), .Q(cpuregs_3[19]));
DFFcell _34310_ (.C(clk), .D(_00963_), .Q(cpuregs_3[20]));
DFFcell _34311_ (.C(clk), .D(_00964_), .Q(cpuregs_3[21]));
DFFcell _34312_ (.C(clk), .D(_00965_), .Q(cpuregs_3[22]));
DFFcell _34313_ (.C(clk), .D(_00966_), .Q(cpuregs_3[23]));
DFFcell _34314_ (.C(clk), .D(_00967_), .Q(cpuregs_3[24]));
DFFcell _34315_ (.C(clk), .D(_00968_), .Q(cpuregs_3[25]));
DFFcell _34316_ (.C(clk), .D(_00969_), .Q(cpuregs_3[26]));
DFFcell _34317_ (.C(clk), .D(_00970_), .Q(cpuregs_3[27]));
DFFcell _34318_ (.C(clk), .D(_00971_), .Q(cpuregs_3[28]));
DFFcell _34319_ (.C(clk), .D(_00972_), .Q(cpuregs_3[29]));
DFFcell _34320_ (.C(clk), .D(_00973_), .Q(cpuregs_3[30]));
DFFcell _34321_ (.C(clk), .D(_00974_), .Q(cpuregs_3[31]));
DFFcell _34322_ (.C(clk), .D(_00975_), .Q(cpuregs_28[0]));
DFFcell _34323_ (.C(clk), .D(_00976_), .Q(cpuregs_28[1]));
DFFcell _34324_ (.C(clk), .D(_00977_), .Q(cpuregs_28[2]));
DFFcell _34325_ (.C(clk), .D(_00978_), .Q(cpuregs_28[3]));
DFFcell _34326_ (.C(clk), .D(_00979_), .Q(cpuregs_28[4]));
DFFcell _34327_ (.C(clk), .D(_00980_), .Q(cpuregs_28[5]));
DFFcell _34328_ (.C(clk), .D(_00981_), .Q(cpuregs_28[6]));
DFFcell _34329_ (.C(clk), .D(_00982_), .Q(cpuregs_28[7]));
DFFcell _34330_ (.C(clk), .D(_00983_), .Q(cpuregs_28[8]));
DFFcell _34331_ (.C(clk), .D(_00984_), .Q(cpuregs_28[9]));
DFFcell _34332_ (.C(clk), .D(_00985_), .Q(cpuregs_28[10]));
DFFcell _34333_ (.C(clk), .D(_00986_), .Q(cpuregs_28[11]));
DFFcell _34334_ (.C(clk), .D(_00987_), .Q(cpuregs_28[12]));
DFFcell _34335_ (.C(clk), .D(_00988_), .Q(cpuregs_28[13]));
DFFcell _34336_ (.C(clk), .D(_00989_), .Q(cpuregs_28[14]));
DFFcell _34337_ (.C(clk), .D(_00990_), .Q(cpuregs_28[15]));
DFFcell _34338_ (.C(clk), .D(_00991_), .Q(cpuregs_28[16]));
DFFcell _34339_ (.C(clk), .D(_00992_), .Q(cpuregs_28[17]));
DFFcell _34340_ (.C(clk), .D(_00993_), .Q(cpuregs_28[18]));
DFFcell _34341_ (.C(clk), .D(_00994_), .Q(cpuregs_28[19]));
DFFcell _34342_ (.C(clk), .D(_00995_), .Q(cpuregs_28[20]));
DFFcell _34343_ (.C(clk), .D(_00996_), .Q(cpuregs_28[21]));
DFFcell _34344_ (.C(clk), .D(_00997_), .Q(cpuregs_28[22]));
DFFcell _34345_ (.C(clk), .D(_00998_), .Q(cpuregs_28[23]));
DFFcell _34346_ (.C(clk), .D(_00999_), .Q(cpuregs_28[24]));
DFFcell _34347_ (.C(clk), .D(_01000_), .Q(cpuregs_28[25]));
DFFcell _34348_ (.C(clk), .D(_01001_), .Q(cpuregs_28[26]));
DFFcell _34349_ (.C(clk), .D(_01002_), .Q(cpuregs_28[27]));
DFFcell _34350_ (.C(clk), .D(_01003_), .Q(cpuregs_28[28]));
DFFcell _34351_ (.C(clk), .D(_01004_), .Q(cpuregs_28[29]));
DFFcell _34352_ (.C(clk), .D(_01005_), .Q(cpuregs_28[30]));
DFFcell _34353_ (.C(clk), .D(_01006_), .Q(cpuregs_28[31]));
DFFcell _34354_ (.C(clk), .D(_01007_), .Q(cpuregs_14[0]));
DFFcell _34355_ (.C(clk), .D(_01008_), .Q(cpuregs_14[1]));
DFFcell _34356_ (.C(clk), .D(_01009_), .Q(cpuregs_14[2]));
DFFcell _34357_ (.C(clk), .D(_01010_), .Q(cpuregs_14[3]));
DFFcell _34358_ (.C(clk), .D(_01011_), .Q(cpuregs_14[4]));
DFFcell _34359_ (.C(clk), .D(_01012_), .Q(cpuregs_14[5]));
DFFcell _34360_ (.C(clk), .D(_01013_), .Q(cpuregs_14[6]));
DFFcell _34361_ (.C(clk), .D(_01014_), .Q(cpuregs_14[7]));
DFFcell _34362_ (.C(clk), .D(_01015_), .Q(cpuregs_14[8]));
DFFcell _34363_ (.C(clk), .D(_01016_), .Q(cpuregs_14[9]));
DFFcell _34364_ (.C(clk), .D(_01017_), .Q(cpuregs_14[10]));
DFFcell _34365_ (.C(clk), .D(_01018_), .Q(cpuregs_14[11]));
DFFcell _34366_ (.C(clk), .D(_01019_), .Q(cpuregs_14[12]));
DFFcell _34367_ (.C(clk), .D(_01020_), .Q(cpuregs_14[13]));
DFFcell _34368_ (.C(clk), .D(_01021_), .Q(cpuregs_14[14]));
DFFcell _34369_ (.C(clk), .D(_01022_), .Q(cpuregs_14[15]));
DFFcell _34370_ (.C(clk), .D(_01023_), .Q(cpuregs_14[16]));
DFFcell _34371_ (.C(clk), .D(_01024_), .Q(cpuregs_14[17]));
DFFcell _34372_ (.C(clk), .D(_01025_), .Q(cpuregs_14[18]));
DFFcell _34373_ (.C(clk), .D(_01026_), .Q(cpuregs_14[19]));
DFFcell _34374_ (.C(clk), .D(_01027_), .Q(cpuregs_14[20]));
DFFcell _34375_ (.C(clk), .D(_01028_), .Q(cpuregs_14[21]));
DFFcell _34376_ (.C(clk), .D(_01029_), .Q(cpuregs_14[22]));
DFFcell _34377_ (.C(clk), .D(_01030_), .Q(cpuregs_14[23]));
DFFcell _34378_ (.C(clk), .D(_01031_), .Q(cpuregs_14[24]));
DFFcell _34379_ (.C(clk), .D(_01032_), .Q(cpuregs_14[25]));
DFFcell _34380_ (.C(clk), .D(_01033_), .Q(cpuregs_14[26]));
DFFcell _34381_ (.C(clk), .D(_01034_), .Q(cpuregs_14[27]));
DFFcell _34382_ (.C(clk), .D(_01035_), .Q(cpuregs_14[28]));
DFFcell _34383_ (.C(clk), .D(_01036_), .Q(cpuregs_14[29]));
DFFcell _34384_ (.C(clk), .D(_01037_), .Q(cpuregs_14[30]));
DFFcell _34385_ (.C(clk), .D(_01038_), .Q(cpuregs_14[31]));
DFFcell _34386_ (.C(clk), .D(_01039_), .Q(cpuregs_26[0]));
DFFcell _34387_ (.C(clk), .D(_01040_), .Q(cpuregs_26[1]));
DFFcell _34388_ (.C(clk), .D(_01041_), .Q(cpuregs_26[2]));
DFFcell _34389_ (.C(clk), .D(_01042_), .Q(cpuregs_26[3]));
DFFcell _34390_ (.C(clk), .D(_01043_), .Q(cpuregs_26[4]));
DFFcell _34391_ (.C(clk), .D(_01044_), .Q(cpuregs_26[5]));
DFFcell _34392_ (.C(clk), .D(_01045_), .Q(cpuregs_26[6]));
DFFcell _34393_ (.C(clk), .D(_01046_), .Q(cpuregs_26[7]));
DFFcell _34394_ (.C(clk), .D(_01047_), .Q(cpuregs_26[8]));
DFFcell _34395_ (.C(clk), .D(_01048_), .Q(cpuregs_26[9]));
DFFcell _34396_ (.C(clk), .D(_01049_), .Q(cpuregs_26[10]));
DFFcell _34397_ (.C(clk), .D(_01050_), .Q(cpuregs_26[11]));
DFFcell _34398_ (.C(clk), .D(_01051_), .Q(cpuregs_26[12]));
DFFcell _34399_ (.C(clk), .D(_01052_), .Q(cpuregs_26[13]));
DFFcell _34400_ (.C(clk), .D(_01053_), .Q(cpuregs_26[14]));
DFFcell _34401_ (.C(clk), .D(_01054_), .Q(cpuregs_26[15]));
DFFcell _34402_ (.C(clk), .D(_01055_), .Q(cpuregs_26[16]));
DFFcell _34403_ (.C(clk), .D(_01056_), .Q(cpuregs_26[17]));
DFFcell _34404_ (.C(clk), .D(_01057_), .Q(cpuregs_26[18]));
DFFcell _34405_ (.C(clk), .D(_01058_), .Q(cpuregs_26[19]));
DFFcell _34406_ (.C(clk), .D(_01059_), .Q(cpuregs_26[20]));
DFFcell _34407_ (.C(clk), .D(_01060_), .Q(cpuregs_26[21]));
DFFcell _34408_ (.C(clk), .D(_01061_), .Q(cpuregs_26[22]));
DFFcell _34409_ (.C(clk), .D(_01062_), .Q(cpuregs_26[23]));
DFFcell _34410_ (.C(clk), .D(_01063_), .Q(cpuregs_26[24]));
DFFcell _34411_ (.C(clk), .D(_01064_), .Q(cpuregs_26[25]));
DFFcell _34412_ (.C(clk), .D(_01065_), .Q(cpuregs_26[26]));
DFFcell _34413_ (.C(clk), .D(_01066_), .Q(cpuregs_26[27]));
DFFcell _34414_ (.C(clk), .D(_01067_), .Q(cpuregs_26[28]));
DFFcell _34415_ (.C(clk), .D(_01068_), .Q(cpuregs_26[29]));
DFFcell _34416_ (.C(clk), .D(_01069_), .Q(cpuregs_26[30]));
DFFcell _34417_ (.C(clk), .D(_01070_), .Q(cpuregs_26[31]));
DFFcell _34418_ (.C(clk), .D(_01071_), .Q(cpuregs_5[0]));
DFFcell _34419_ (.C(clk), .D(_01072_), .Q(cpuregs_5[1]));
DFFcell _34420_ (.C(clk), .D(_01073_), .Q(cpuregs_5[2]));
DFFcell _34421_ (.C(clk), .D(_01074_), .Q(cpuregs_5[3]));
DFFcell _34422_ (.C(clk), .D(_01075_), .Q(cpuregs_5[4]));
DFFcell _34423_ (.C(clk), .D(_01076_), .Q(cpuregs_5[5]));
DFFcell _34424_ (.C(clk), .D(_01077_), .Q(cpuregs_5[6]));
DFFcell _34425_ (.C(clk), .D(_01078_), .Q(cpuregs_5[7]));
DFFcell _34426_ (.C(clk), .D(_01079_), .Q(cpuregs_5[8]));
DFFcell _34427_ (.C(clk), .D(_01080_), .Q(cpuregs_5[9]));
DFFcell _34428_ (.C(clk), .D(_01081_), .Q(cpuregs_5[10]));
DFFcell _34429_ (.C(clk), .D(_01082_), .Q(cpuregs_5[11]));
DFFcell _34430_ (.C(clk), .D(_01083_), .Q(cpuregs_5[12]));
DFFcell _34431_ (.C(clk), .D(_01084_), .Q(cpuregs_5[13]));
DFFcell _34432_ (.C(clk), .D(_01085_), .Q(cpuregs_5[14]));
DFFcell _34433_ (.C(clk), .D(_01086_), .Q(cpuregs_5[15]));
DFFcell _34434_ (.C(clk), .D(_01087_), .Q(cpuregs_5[16]));
DFFcell _34435_ (.C(clk), .D(_01088_), .Q(cpuregs_5[17]));
DFFcell _34436_ (.C(clk), .D(_01089_), .Q(cpuregs_5[18]));
DFFcell _34437_ (.C(clk), .D(_01090_), .Q(cpuregs_5[19]));
DFFcell _34438_ (.C(clk), .D(_01091_), .Q(cpuregs_5[20]));
DFFcell _34439_ (.C(clk), .D(_01092_), .Q(cpuregs_5[21]));
DFFcell _34440_ (.C(clk), .D(_01093_), .Q(cpuregs_5[22]));
DFFcell _34441_ (.C(clk), .D(_01094_), .Q(cpuregs_5[23]));
DFFcell _34442_ (.C(clk), .D(_01095_), .Q(cpuregs_5[24]));
DFFcell _34443_ (.C(clk), .D(_01096_), .Q(cpuregs_5[25]));
DFFcell _34444_ (.C(clk), .D(_01097_), .Q(cpuregs_5[26]));
DFFcell _34445_ (.C(clk), .D(_01098_), .Q(cpuregs_5[27]));
DFFcell _34446_ (.C(clk), .D(_01099_), .Q(cpuregs_5[28]));
DFFcell _34447_ (.C(clk), .D(_01100_), .Q(cpuregs_5[29]));
DFFcell _34448_ (.C(clk), .D(_01101_), .Q(cpuregs_5[30]));
DFFcell _34449_ (.C(clk), .D(_01102_), .Q(cpuregs_5[31]));
DFFcell _34450_ (.C(clk), .D(_01103_), .Q(cpuregs_12[0]));
DFFcell _34451_ (.C(clk), .D(_01104_), .Q(cpuregs_12[1]));
DFFcell _34452_ (.C(clk), .D(_01105_), .Q(cpuregs_12[2]));
DFFcell _34453_ (.C(clk), .D(_01106_), .Q(cpuregs_12[3]));
DFFcell _34454_ (.C(clk), .D(_01107_), .Q(cpuregs_12[4]));
DFFcell _34455_ (.C(clk), .D(_01108_), .Q(cpuregs_12[5]));
DFFcell _34456_ (.C(clk), .D(_01109_), .Q(cpuregs_12[6]));
DFFcell _34457_ (.C(clk), .D(_01110_), .Q(cpuregs_12[7]));
DFFcell _34458_ (.C(clk), .D(_01111_), .Q(cpuregs_12[8]));
DFFcell _34459_ (.C(clk), .D(_01112_), .Q(cpuregs_12[9]));
DFFcell _34460_ (.C(clk), .D(_01113_), .Q(cpuregs_12[10]));
DFFcell _34461_ (.C(clk), .D(_01114_), .Q(cpuregs_12[11]));
DFFcell _34462_ (.C(clk), .D(_01115_), .Q(cpuregs_12[12]));
DFFcell _34463_ (.C(clk), .D(_01116_), .Q(cpuregs_12[13]));
DFFcell _34464_ (.C(clk), .D(_01117_), .Q(cpuregs_12[14]));
DFFcell _34465_ (.C(clk), .D(_01118_), .Q(cpuregs_12[15]));
DFFcell _34466_ (.C(clk), .D(_01119_), .Q(cpuregs_12[16]));
DFFcell _34467_ (.C(clk), .D(_01120_), .Q(cpuregs_12[17]));
DFFcell _34468_ (.C(clk), .D(_01121_), .Q(cpuregs_12[18]));
DFFcell _34469_ (.C(clk), .D(_01122_), .Q(cpuregs_12[19]));
DFFcell _34470_ (.C(clk), .D(_01123_), .Q(cpuregs_12[20]));
DFFcell _34471_ (.C(clk), .D(_01124_), .Q(cpuregs_12[21]));
DFFcell _34472_ (.C(clk), .D(_01125_), .Q(cpuregs_12[22]));
DFFcell _34473_ (.C(clk), .D(_01126_), .Q(cpuregs_12[23]));
DFFcell _34474_ (.C(clk), .D(_01127_), .Q(cpuregs_12[24]));
DFFcell _34475_ (.C(clk), .D(_01128_), .Q(cpuregs_12[25]));
DFFcell _34476_ (.C(clk), .D(_01129_), .Q(cpuregs_12[26]));
DFFcell _34477_ (.C(clk), .D(_01130_), .Q(cpuregs_12[27]));
DFFcell _34478_ (.C(clk), .D(_01131_), .Q(cpuregs_12[28]));
DFFcell _34479_ (.C(clk), .D(_01132_), .Q(cpuregs_12[29]));
DFFcell _34480_ (.C(clk), .D(_01133_), .Q(cpuregs_12[30]));
DFFcell _34481_ (.C(clk), .D(_01134_), .Q(cpuregs_12[31]));
DFFcell _34482_ (.C(clk), .D(_01135_), .Q(cpuregs_7[0]));
DFFcell _34483_ (.C(clk), .D(_01136_), .Q(cpuregs_7[1]));
DFFcell _34484_ (.C(clk), .D(_01137_), .Q(cpuregs_7[2]));
DFFcell _34485_ (.C(clk), .D(_01138_), .Q(cpuregs_7[3]));
DFFcell _34486_ (.C(clk), .D(_01139_), .Q(cpuregs_7[4]));
DFFcell _34487_ (.C(clk), .D(_01140_), .Q(cpuregs_7[5]));
DFFcell _34488_ (.C(clk), .D(_01141_), .Q(cpuregs_7[6]));
DFFcell _34489_ (.C(clk), .D(_01142_), .Q(cpuregs_7[7]));
DFFcell _34490_ (.C(clk), .D(_01143_), .Q(cpuregs_7[8]));
DFFcell _34491_ (.C(clk), .D(_01144_), .Q(cpuregs_7[9]));
DFFcell _34492_ (.C(clk), .D(_01145_), .Q(cpuregs_7[10]));
DFFcell _34493_ (.C(clk), .D(_01146_), .Q(cpuregs_7[11]));
DFFcell _34494_ (.C(clk), .D(_01147_), .Q(cpuregs_7[12]));
DFFcell _34495_ (.C(clk), .D(_01148_), .Q(cpuregs_7[13]));
DFFcell _34496_ (.C(clk), .D(_01149_), .Q(cpuregs_7[14]));
DFFcell _34497_ (.C(clk), .D(_01150_), .Q(cpuregs_7[15]));
DFFcell _34498_ (.C(clk), .D(_01151_), .Q(cpuregs_7[16]));
DFFcell _34499_ (.C(clk), .D(_01152_), .Q(cpuregs_7[17]));
DFFcell _34500_ (.C(clk), .D(_01153_), .Q(cpuregs_7[18]));
DFFcell _34501_ (.C(clk), .D(_01154_), .Q(cpuregs_7[19]));
DFFcell _34502_ (.C(clk), .D(_01155_), .Q(cpuregs_7[20]));
DFFcell _34503_ (.C(clk), .D(_01156_), .Q(cpuregs_7[21]));
DFFcell _34504_ (.C(clk), .D(_01157_), .Q(cpuregs_7[22]));
DFFcell _34505_ (.C(clk), .D(_01158_), .Q(cpuregs_7[23]));
DFFcell _34506_ (.C(clk), .D(_01159_), .Q(cpuregs_7[24]));
DFFcell _34507_ (.C(clk), .D(_01160_), .Q(cpuregs_7[25]));
DFFcell _34508_ (.C(clk), .D(_01161_), .Q(cpuregs_7[26]));
DFFcell _34509_ (.C(clk), .D(_01162_), .Q(cpuregs_7[27]));
DFFcell _34510_ (.C(clk), .D(_01163_), .Q(cpuregs_7[28]));
DFFcell _34511_ (.C(clk), .D(_01164_), .Q(cpuregs_7[29]));
DFFcell _34512_ (.C(clk), .D(_01165_), .Q(cpuregs_7[30]));
DFFcell _34513_ (.C(clk), .D(_01166_), .Q(cpuregs_7[31]));
DFFcell _34514_ (.C(clk), .D(_01167_), .Q(cpu_state[0]));
DFFcell _34515_ (.C(clk), .D(_01168_), .Q(cpu_state[1]));
DFFcell _34516_ (.C(clk), .D(_01169_), .Q(cpu_state[2]));
DFFcell _34517_ (.C(clk), .D(_01170_), .Q(cpu_state[3]));
DFFcell _34518_ (.C(clk), .D(_01171_), .Q(cpu_state[4]));
DFFcell _34519_ (.C(clk), .D(_01172_), .Q(cpu_state[5]));
DFFcell _34520_ (.C(clk), .D(_01173_), .Q(cpu_state[6]));
DFFcell _34521_ (.C(clk), .D(_01174_), .Q(cpu_state[7]));
DFFcell _34522_ (.C(clk), .D(_01175_), .Q(cpuregs_8[0]));
DFFcell _34523_ (.C(clk), .D(_01176_), .Q(cpuregs_8[1]));
DFFcell _34524_ (.C(clk), .D(_01177_), .Q(cpuregs_8[2]));
DFFcell _34525_ (.C(clk), .D(_01178_), .Q(cpuregs_8[3]));
DFFcell _34526_ (.C(clk), .D(_01179_), .Q(cpuregs_8[4]));
DFFcell _34527_ (.C(clk), .D(_01180_), .Q(cpuregs_8[5]));
DFFcell _34528_ (.C(clk), .D(_01181_), .Q(cpuregs_8[6]));
DFFcell _34529_ (.C(clk), .D(_01182_), .Q(cpuregs_8[7]));
DFFcell _34530_ (.C(clk), .D(_01183_), .Q(cpuregs_8[8]));
DFFcell _34531_ (.C(clk), .D(_01184_), .Q(cpuregs_8[9]));
DFFcell _34532_ (.C(clk), .D(_01185_), .Q(cpuregs_8[10]));
DFFcell _34533_ (.C(clk), .D(_01186_), .Q(cpuregs_8[11]));
DFFcell _34534_ (.C(clk), .D(_01187_), .Q(cpuregs_8[12]));
DFFcell _34535_ (.C(clk), .D(_01188_), .Q(cpuregs_8[13]));
DFFcell _34536_ (.C(clk), .D(_01189_), .Q(cpuregs_8[14]));
DFFcell _34537_ (.C(clk), .D(_01190_), .Q(cpuregs_8[15]));
DFFcell _34538_ (.C(clk), .D(_01191_), .Q(cpuregs_8[16]));
DFFcell _34539_ (.C(clk), .D(_01192_), .Q(cpuregs_8[17]));
DFFcell _34540_ (.C(clk), .D(_01193_), .Q(cpuregs_8[18]));
DFFcell _34541_ (.C(clk), .D(_01194_), .Q(cpuregs_8[19]));
DFFcell _34542_ (.C(clk), .D(_01195_), .Q(cpuregs_8[20]));
DFFcell _34543_ (.C(clk), .D(_01196_), .Q(cpuregs_8[21]));
DFFcell _34544_ (.C(clk), .D(_01197_), .Q(cpuregs_8[22]));
DFFcell _34545_ (.C(clk), .D(_01198_), .Q(cpuregs_8[23]));
DFFcell _34546_ (.C(clk), .D(_01199_), .Q(cpuregs_8[24]));
DFFcell _34547_ (.C(clk), .D(_01200_), .Q(cpuregs_8[25]));
DFFcell _34548_ (.C(clk), .D(_01201_), .Q(cpuregs_8[26]));
DFFcell _34549_ (.C(clk), .D(_01202_), .Q(cpuregs_8[27]));
DFFcell _34550_ (.C(clk), .D(_01203_), .Q(cpuregs_8[28]));
DFFcell _34551_ (.C(clk), .D(_01204_), .Q(cpuregs_8[29]));
DFFcell _34552_ (.C(clk), .D(_01205_), .Q(cpuregs_8[30]));
DFFcell _34553_ (.C(clk), .D(_01206_), .Q(cpuregs_8[31]));
DFFcell _34554_ (.C(clk), .D(_01207_), .Q(pcpi_rs1[0]));
DFFcell _34555_ (.C(clk), .D(_01208_), .Q(pcpi_rs1[1]));
DFFcell _34556_ (.C(clk), .D(_01209_), .Q(pcpi_rs1[2]));
DFFcell _34557_ (.C(clk), .D(_01210_), .Q(pcpi_rs1[3]));
DFFcell _34558_ (.C(clk), .D(_01211_), .Q(pcpi_rs1[4]));
DFFcell _34559_ (.C(clk), .D(_01212_), .Q(pcpi_rs1[5]));
DFFcell _34560_ (.C(clk), .D(_01213_), .Q(pcpi_rs1[6]));
DFFcell _34561_ (.C(clk), .D(_01214_), .Q(pcpi_rs1[7]));
DFFcell _34562_ (.C(clk), .D(_01215_), .Q(pcpi_rs1[8]));
DFFcell _34563_ (.C(clk), .D(_01216_), .Q(pcpi_rs1[9]));
DFFcell _34564_ (.C(clk), .D(_01217_), .Q(pcpi_rs1[10]));
DFFcell _34565_ (.C(clk), .D(_01218_), .Q(pcpi_rs1[11]));
DFFcell _34566_ (.C(clk), .D(_01219_), .Q(pcpi_rs1[12]));
DFFcell _34567_ (.C(clk), .D(_01220_), .Q(pcpi_rs1[13]));
DFFcell _34568_ (.C(clk), .D(_01221_), .Q(pcpi_rs1[14]));
DFFcell _34569_ (.C(clk), .D(_01222_), .Q(pcpi_rs1[15]));
DFFcell _34570_ (.C(clk), .D(_01223_), .Q(pcpi_rs1[16]));
DFFcell _34571_ (.C(clk), .D(_01224_), .Q(pcpi_rs1[17]));
DFFcell _34572_ (.C(clk), .D(_01225_), .Q(pcpi_rs1[18]));
DFFcell _34573_ (.C(clk), .D(_01226_), .Q(pcpi_rs1[19]));
DFFcell _34574_ (.C(clk), .D(_01227_), .Q(pcpi_rs1[20]));
DFFcell _34575_ (.C(clk), .D(_01228_), .Q(pcpi_rs1[21]));
DFFcell _34576_ (.C(clk), .D(_01229_), .Q(pcpi_rs1[22]));
DFFcell _34577_ (.C(clk), .D(_01230_), .Q(pcpi_rs1[23]));
DFFcell _34578_ (.C(clk), .D(_01231_), .Q(pcpi_rs1[24]));
DFFcell _34579_ (.C(clk), .D(_01232_), .Q(pcpi_rs1[25]));
DFFcell _34580_ (.C(clk), .D(_01233_), .Q(pcpi_rs1[26]));
DFFcell _34581_ (.C(clk), .D(_01234_), .Q(pcpi_rs1[27]));
DFFcell _34582_ (.C(clk), .D(_01235_), .Q(pcpi_rs1[28]));
DFFcell _34583_ (.C(clk), .D(_01236_), .Q(pcpi_rs1[29]));
DFFcell _34584_ (.C(clk), .D(_01237_), .Q(pcpi_rs1[30]));
DFFcell _34585_ (.C(clk), .D(_01238_), .Q(cpuregs_0[0]));
DFFcell _34586_ (.C(clk), .D(_01239_), .Q(cpuregs_0[1]));
DFFcell _34587_ (.C(clk), .D(_01240_), .Q(cpuregs_0[2]));
DFFcell _34588_ (.C(clk), .D(_01241_), .Q(cpuregs_0[3]));
DFFcell _34589_ (.C(clk), .D(_01242_), .Q(cpuregs_0[4]));
DFFcell _34590_ (.C(clk), .D(_01243_), .Q(cpuregs_0[5]));
DFFcell _34591_ (.C(clk), .D(_01244_), .Q(cpuregs_0[6]));
DFFcell _34592_ (.C(clk), .D(_01245_), .Q(cpuregs_0[7]));
DFFcell _34593_ (.C(clk), .D(_01246_), .Q(cpuregs_0[8]));
DFFcell _34594_ (.C(clk), .D(_01247_), .Q(cpuregs_0[9]));
DFFcell _34595_ (.C(clk), .D(_01248_), .Q(cpuregs_0[10]));
DFFcell _34596_ (.C(clk), .D(_01249_), .Q(cpuregs_0[11]));
DFFcell _34597_ (.C(clk), .D(_01250_), .Q(cpuregs_0[12]));
DFFcell _34598_ (.C(clk), .D(_01251_), .Q(cpuregs_0[13]));
DFFcell _34599_ (.C(clk), .D(_01252_), .Q(cpuregs_0[14]));
DFFcell _34600_ (.C(clk), .D(_01253_), .Q(cpuregs_0[15]));
DFFcell _34601_ (.C(clk), .D(_01254_), .Q(cpuregs_0[16]));
DFFcell _34602_ (.C(clk), .D(_01255_), .Q(cpuregs_0[17]));
DFFcell _34603_ (.C(clk), .D(_01256_), .Q(cpuregs_0[18]));
DFFcell _34604_ (.C(clk), .D(_01257_), .Q(cpuregs_0[19]));
DFFcell _34605_ (.C(clk), .D(_01258_), .Q(cpuregs_0[20]));
DFFcell _34606_ (.C(clk), .D(_01259_), .Q(cpuregs_0[21]));
DFFcell _34607_ (.C(clk), .D(_01260_), .Q(cpuregs_0[22]));
DFFcell _34608_ (.C(clk), .D(_01261_), .Q(cpuregs_0[23]));
DFFcell _34609_ (.C(clk), .D(_01262_), .Q(cpuregs_0[24]));
DFFcell _34610_ (.C(clk), .D(_01263_), .Q(cpuregs_0[25]));
DFFcell _34611_ (.C(clk), .D(_01264_), .Q(cpuregs_0[26]));
DFFcell _34612_ (.C(clk), .D(_01265_), .Q(cpuregs_0[27]));
DFFcell _34613_ (.C(clk), .D(_01266_), .Q(cpuregs_0[28]));
DFFcell _34614_ (.C(clk), .D(_01267_), .Q(cpuregs_0[29]));
DFFcell _34615_ (.C(clk), .D(_01268_), .Q(cpuregs_0[30]));
DFFcell _34616_ (.C(clk), .D(_01269_), .Q(cpuregs_0[31]));
DFFcell _34617_ (.C(clk), .D(_01270_), .Q(decoded_imm_j[6]));
DFFcell _34618_ (.C(clk), .D(_01271_), .Q(decoded_imm_j[7]));
DFFcell _34619_ (.C(clk), .D(_01272_), .Q(decoded_imm_j[10]));
DFFcell _34620_ (.C(clk), .D(_01273_), .Q(decoded_imm_j[4]));
DFFcell _34621_ (.C(clk), .D(_01274_), .Q(decoded_imm_j[31]));
DFFcell _34622_ (.C(clk), .D(_01275_), .Q(cpuregs_13[0]));
DFFcell _34623_ (.C(clk), .D(_01276_), .Q(cpuregs_13[1]));
DFFcell _34624_ (.C(clk), .D(_01277_), .Q(cpuregs_13[2]));
DFFcell _34625_ (.C(clk), .D(_01278_), .Q(cpuregs_13[3]));
DFFcell _34626_ (.C(clk), .D(_01279_), .Q(cpuregs_13[4]));
DFFcell _34627_ (.C(clk), .D(_01280_), .Q(cpuregs_13[5]));
DFFcell _34628_ (.C(clk), .D(_01281_), .Q(cpuregs_13[6]));
DFFcell _34629_ (.C(clk), .D(_01282_), .Q(cpuregs_13[7]));
DFFcell _34630_ (.C(clk), .D(_01283_), .Q(cpuregs_13[8]));
DFFcell _34631_ (.C(clk), .D(_01284_), .Q(cpuregs_13[9]));
DFFcell _34632_ (.C(clk), .D(_01285_), .Q(cpuregs_13[10]));
DFFcell _34633_ (.C(clk), .D(_01286_), .Q(cpuregs_13[11]));
DFFcell _34634_ (.C(clk), .D(_01287_), .Q(cpuregs_13[12]));
DFFcell _34635_ (.C(clk), .D(_01288_), .Q(cpuregs_13[13]));
DFFcell _34636_ (.C(clk), .D(_01289_), .Q(cpuregs_13[14]));
DFFcell _34637_ (.C(clk), .D(_01290_), .Q(cpuregs_13[15]));
DFFcell _34638_ (.C(clk), .D(_01291_), .Q(cpuregs_13[16]));
DFFcell _34639_ (.C(clk), .D(_01292_), .Q(cpuregs_13[17]));
DFFcell _34640_ (.C(clk), .D(_01293_), .Q(cpuregs_13[18]));
DFFcell _34641_ (.C(clk), .D(_01294_), .Q(cpuregs_13[19]));
DFFcell _34642_ (.C(clk), .D(_01295_), .Q(cpuregs_13[20]));
DFFcell _34643_ (.C(clk), .D(_01296_), .Q(cpuregs_13[21]));
DFFcell _34644_ (.C(clk), .D(_01297_), .Q(cpuregs_13[22]));
DFFcell _34645_ (.C(clk), .D(_01298_), .Q(cpuregs_13[23]));
DFFcell _34646_ (.C(clk), .D(_01299_), .Q(cpuregs_13[24]));
DFFcell _34647_ (.C(clk), .D(_01300_), .Q(cpuregs_13[25]));
DFFcell _34648_ (.C(clk), .D(_01301_), .Q(cpuregs_13[26]));
DFFcell _34649_ (.C(clk), .D(_01302_), .Q(cpuregs_13[27]));
DFFcell _34650_ (.C(clk), .D(_01303_), .Q(cpuregs_13[28]));
DFFcell _34651_ (.C(clk), .D(_01304_), .Q(cpuregs_13[29]));
DFFcell _34652_ (.C(clk), .D(_01305_), .Q(cpuregs_13[30]));
DFFcell _34653_ (.C(clk), .D(_01306_), .Q(cpuregs_13[31]));
DFFcell _34654_ (.C(clk), .D(_01307_), .Q(decoded_imm_j[12]));
DFFcell _34655_ (.C(clk), .D(_01308_), .Q(decoded_imm_j[13]));
DFFcell _34656_ (.C(clk), .D(_01309_), .Q(decoded_imm_j[14]));
DFFcell _34657_ (.C(clk), .D(_01310_), .Q(decoded_imm_j[18]));
DFFcell _34658_ (.C(clk), .D(_01311_), .Q(decoded_imm_j[19]));
DFFcell _34659_ (.C(clk), .D(_01312_), .Q(decoded_imm_j[15]));
DFFcell _34660_ (.C(clk), .D(_01313_), .Q(decoded_imm_j[16]));
DFFcell _34661_ (.C(clk), .D(_01314_), .Q(decoded_imm_j[17]));
DFFcell _34662_ (.C(clk), .D(_01315_), .Q(cpuregs_15[0]));
DFFcell _34663_ (.C(clk), .D(_01316_), .Q(cpuregs_15[1]));
DFFcell _34664_ (.C(clk), .D(_01317_), .Q(cpuregs_15[2]));
DFFcell _34665_ (.C(clk), .D(_01318_), .Q(cpuregs_15[3]));
DFFcell _34666_ (.C(clk), .D(_01319_), .Q(cpuregs_15[4]));
DFFcell _34667_ (.C(clk), .D(_01320_), .Q(cpuregs_15[5]));
DFFcell _34668_ (.C(clk), .D(_01321_), .Q(cpuregs_15[6]));
DFFcell _34669_ (.C(clk), .D(_01322_), .Q(cpuregs_15[7]));
DFFcell _34670_ (.C(clk), .D(_01323_), .Q(cpuregs_15[8]));
DFFcell _34671_ (.C(clk), .D(_01324_), .Q(cpuregs_15[9]));
DFFcell _34672_ (.C(clk), .D(_01325_), .Q(cpuregs_15[10]));
DFFcell _34673_ (.C(clk), .D(_01326_), .Q(cpuregs_15[11]));
DFFcell _34674_ (.C(clk), .D(_01327_), .Q(cpuregs_15[12]));
DFFcell _34675_ (.C(clk), .D(_01328_), .Q(cpuregs_15[13]));
DFFcell _34676_ (.C(clk), .D(_01329_), .Q(cpuregs_15[14]));
DFFcell _34677_ (.C(clk), .D(_01330_), .Q(cpuregs_15[15]));
DFFcell _34678_ (.C(clk), .D(_01331_), .Q(cpuregs_15[16]));
DFFcell _34679_ (.C(clk), .D(_01332_), .Q(cpuregs_15[17]));
DFFcell _34680_ (.C(clk), .D(_01333_), .Q(cpuregs_15[18]));
DFFcell _34681_ (.C(clk), .D(_01334_), .Q(cpuregs_15[19]));
DFFcell _34682_ (.C(clk), .D(_01335_), .Q(cpuregs_15[20]));
DFFcell _34683_ (.C(clk), .D(_01336_), .Q(cpuregs_15[21]));
DFFcell _34684_ (.C(clk), .D(_01337_), .Q(cpuregs_15[22]));
DFFcell _34685_ (.C(clk), .D(_01338_), .Q(cpuregs_15[23]));
DFFcell _34686_ (.C(clk), .D(_01339_), .Q(cpuregs_15[24]));
DFFcell _34687_ (.C(clk), .D(_01340_), .Q(cpuregs_15[25]));
DFFcell _34688_ (.C(clk), .D(_01341_), .Q(cpuregs_15[26]));
DFFcell _34689_ (.C(clk), .D(_01342_), .Q(cpuregs_15[27]));
DFFcell _34690_ (.C(clk), .D(_01343_), .Q(cpuregs_15[28]));
DFFcell _34691_ (.C(clk), .D(_01344_), .Q(cpuregs_15[29]));
DFFcell _34692_ (.C(clk), .D(_01345_), .Q(cpuregs_15[30]));
DFFcell _34693_ (.C(clk), .D(_01346_), .Q(cpuregs_15[31]));
DFFcell _34694_ (.C(clk), .D(_01347_), .Q(count_instr[0]));
DFFcell _34695_ (.C(clk), .D(_01348_), .Q(count_instr[1]));
DFFcell _34696_ (.C(clk), .D(_01349_), .Q(count_instr[2]));
DFFcell _34697_ (.C(clk), .D(_01350_), .Q(count_instr[3]));
DFFcell _34698_ (.C(clk), .D(_01351_), .Q(count_instr[4]));
DFFcell _34699_ (.C(clk), .D(_01352_), .Q(count_instr[5]));
DFFcell _34700_ (.C(clk), .D(_01353_), .Q(count_instr[6]));
DFFcell _34701_ (.C(clk), .D(_01354_), .Q(count_instr[7]));
DFFcell _34702_ (.C(clk), .D(_01355_), .Q(count_instr[8]));
DFFcell _34703_ (.C(clk), .D(_01356_), .Q(count_instr[9]));
DFFcell _34704_ (.C(clk), .D(_01357_), .Q(count_instr[10]));
DFFcell _34705_ (.C(clk), .D(_01358_), .Q(count_instr[11]));
DFFcell _34706_ (.C(clk), .D(_01359_), .Q(count_instr[12]));
DFFcell _34707_ (.C(clk), .D(_01360_), .Q(count_instr[13]));
DFFcell _34708_ (.C(clk), .D(_01361_), .Q(count_instr[14]));
DFFcell _34709_ (.C(clk), .D(_01362_), .Q(count_instr[15]));
DFFcell _34710_ (.C(clk), .D(_01363_), .Q(count_instr[16]));
DFFcell _34711_ (.C(clk), .D(_01364_), .Q(count_instr[17]));
DFFcell _34712_ (.C(clk), .D(_01365_), .Q(count_instr[18]));
DFFcell _34713_ (.C(clk), .D(_01366_), .Q(count_instr[19]));
DFFcell _34714_ (.C(clk), .D(_01367_), .Q(count_instr[20]));
DFFcell _34715_ (.C(clk), .D(_01368_), .Q(count_instr[21]));
DFFcell _34716_ (.C(clk), .D(_01369_), .Q(count_instr[22]));
DFFcell _34717_ (.C(clk), .D(_01370_), .Q(count_instr[23]));
DFFcell _34718_ (.C(clk), .D(_01371_), .Q(count_instr[24]));
DFFcell _34719_ (.C(clk), .D(_01372_), .Q(count_instr[25]));
DFFcell _34720_ (.C(clk), .D(_01373_), .Q(count_instr[26]));
DFFcell _34721_ (.C(clk), .D(_01374_), .Q(count_instr[27]));
DFFcell _34722_ (.C(clk), .D(_01375_), .Q(count_instr[28]));
DFFcell _34723_ (.C(clk), .D(_01376_), .Q(count_instr[29]));
DFFcell _34724_ (.C(clk), .D(_01377_), .Q(count_instr[30]));
DFFcell _34725_ (.C(clk), .D(_01378_), .Q(count_instr[31]));
DFFcell _34726_ (.C(clk), .D(_01379_), .Q(count_instr[32]));
DFFcell _34727_ (.C(clk), .D(_01380_), .Q(count_instr[33]));
DFFcell _34728_ (.C(clk), .D(_01381_), .Q(count_instr[34]));
DFFcell _34729_ (.C(clk), .D(_01382_), .Q(count_instr[35]));
DFFcell _34730_ (.C(clk), .D(_01383_), .Q(count_instr[36]));
DFFcell _34731_ (.C(clk), .D(_01384_), .Q(count_instr[37]));
DFFcell _34732_ (.C(clk), .D(_01385_), .Q(count_instr[38]));
DFFcell _34733_ (.C(clk), .D(_01386_), .Q(count_instr[39]));
DFFcell _34734_ (.C(clk), .D(_01387_), .Q(count_instr[40]));
DFFcell _34735_ (.C(clk), .D(_01388_), .Q(count_instr[41]));
DFFcell _34736_ (.C(clk), .D(_01389_), .Q(count_instr[42]));
DFFcell _34737_ (.C(clk), .D(_01390_), .Q(count_instr[43]));
DFFcell _34738_ (.C(clk), .D(_01391_), .Q(count_instr[44]));
DFFcell _34739_ (.C(clk), .D(_01392_), .Q(count_instr[45]));
DFFcell _34740_ (.C(clk), .D(_01393_), .Q(count_instr[46]));
DFFcell _34741_ (.C(clk), .D(_01394_), .Q(count_instr[47]));
DFFcell _34742_ (.C(clk), .D(_01395_), .Q(count_instr[48]));
DFFcell _34743_ (.C(clk), .D(_01396_), .Q(count_instr[49]));
DFFcell _34744_ (.C(clk), .D(_01397_), .Q(count_instr[50]));
DFFcell _34745_ (.C(clk), .D(_01398_), .Q(count_instr[51]));
DFFcell _34746_ (.C(clk), .D(_01399_), .Q(count_instr[52]));
DFFcell _34747_ (.C(clk), .D(_01400_), .Q(count_instr[53]));
DFFcell _34748_ (.C(clk), .D(_01401_), .Q(count_instr[54]));
DFFcell _34749_ (.C(clk), .D(_01402_), .Q(count_instr[55]));
DFFcell _34750_ (.C(clk), .D(_01403_), .Q(count_instr[56]));
DFFcell _34751_ (.C(clk), .D(_01404_), .Q(count_instr[57]));
DFFcell _34752_ (.C(clk), .D(_01405_), .Q(count_instr[58]));
DFFcell _34753_ (.C(clk), .D(_01406_), .Q(count_instr[59]));
DFFcell _34754_ (.C(clk), .D(_01407_), .Q(count_instr[60]));
DFFcell _34755_ (.C(clk), .D(_01408_), .Q(count_instr[61]));
DFFcell _34756_ (.C(clk), .D(_01409_), .Q(count_instr[62]));
DFFcell _34757_ (.C(clk), .D(_01410_), .Q(count_instr[63]));
DFFcell _34758_ (.C(clk), .D(_01411_), .Q(cpuregs_30[0]));
DFFcell _34759_ (.C(clk), .D(_01412_), .Q(cpuregs_30[1]));
DFFcell _34760_ (.C(clk), .D(_01413_), .Q(cpuregs_30[2]));
DFFcell _34761_ (.C(clk), .D(_01414_), .Q(cpuregs_30[3]));
DFFcell _34762_ (.C(clk), .D(_01415_), .Q(cpuregs_30[4]));
DFFcell _34763_ (.C(clk), .D(_01416_), .Q(cpuregs_30[5]));
DFFcell _34764_ (.C(clk), .D(_01417_), .Q(cpuregs_30[6]));
DFFcell _34765_ (.C(clk), .D(_01418_), .Q(cpuregs_30[7]));
DFFcell _34766_ (.C(clk), .D(_01419_), .Q(cpuregs_30[8]));
DFFcell _34767_ (.C(clk), .D(_01420_), .Q(cpuregs_30[9]));
DFFcell _34768_ (.C(clk), .D(_01421_), .Q(cpuregs_30[10]));
DFFcell _34769_ (.C(clk), .D(_01422_), .Q(cpuregs_30[11]));
DFFcell _34770_ (.C(clk), .D(_01423_), .Q(cpuregs_30[12]));
DFFcell _34771_ (.C(clk), .D(_01424_), .Q(cpuregs_30[13]));
DFFcell _34772_ (.C(clk), .D(_01425_), .Q(cpuregs_30[14]));
DFFcell _34773_ (.C(clk), .D(_01426_), .Q(cpuregs_30[15]));
DFFcell _34774_ (.C(clk), .D(_01427_), .Q(cpuregs_30[16]));
DFFcell _34775_ (.C(clk), .D(_01428_), .Q(cpuregs_30[17]));
DFFcell _34776_ (.C(clk), .D(_01429_), .Q(cpuregs_30[18]));
DFFcell _34777_ (.C(clk), .D(_01430_), .Q(cpuregs_30[19]));
DFFcell _34778_ (.C(clk), .D(_01431_), .Q(cpuregs_30[20]));
DFFcell _34779_ (.C(clk), .D(_01432_), .Q(cpuregs_30[21]));
DFFcell _34780_ (.C(clk), .D(_01433_), .Q(cpuregs_30[22]));
DFFcell _34781_ (.C(clk), .D(_01434_), .Q(cpuregs_30[23]));
DFFcell _34782_ (.C(clk), .D(_01435_), .Q(cpuregs_30[24]));
DFFcell _34783_ (.C(clk), .D(_01436_), .Q(cpuregs_30[25]));
DFFcell _34784_ (.C(clk), .D(_01437_), .Q(cpuregs_30[26]));
DFFcell _34785_ (.C(clk), .D(_01438_), .Q(cpuregs_30[27]));
DFFcell _34786_ (.C(clk), .D(_01439_), .Q(cpuregs_30[28]));
DFFcell _34787_ (.C(clk), .D(_01440_), .Q(cpuregs_30[29]));
DFFcell _34788_ (.C(clk), .D(_01441_), .Q(cpuregs_30[30]));
DFFcell _34789_ (.C(clk), .D(_01442_), .Q(cpuregs_30[31]));
DFFcell _34790_ (.C(clk), .D(_01443_), .Q(cpuregs_24[0]));
DFFcell _34791_ (.C(clk), .D(_01444_), .Q(cpuregs_24[1]));
DFFcell _34792_ (.C(clk), .D(_01445_), .Q(cpuregs_24[2]));
DFFcell _34793_ (.C(clk), .D(_01446_), .Q(cpuregs_24[3]));
DFFcell _34794_ (.C(clk), .D(_01447_), .Q(cpuregs_24[4]));
DFFcell _34795_ (.C(clk), .D(_01448_), .Q(cpuregs_24[5]));
DFFcell _34796_ (.C(clk), .D(_01449_), .Q(cpuregs_24[6]));
DFFcell _34797_ (.C(clk), .D(_01450_), .Q(cpuregs_24[7]));
DFFcell _34798_ (.C(clk), .D(_01451_), .Q(cpuregs_24[8]));
DFFcell _34799_ (.C(clk), .D(_01452_), .Q(cpuregs_24[9]));
DFFcell _34800_ (.C(clk), .D(_01453_), .Q(cpuregs_24[10]));
DFFcell _34801_ (.C(clk), .D(_01454_), .Q(cpuregs_24[11]));
DFFcell _34802_ (.C(clk), .D(_01455_), .Q(cpuregs_24[12]));
DFFcell _34803_ (.C(clk), .D(_01456_), .Q(cpuregs_24[13]));
DFFcell _34804_ (.C(clk), .D(_01457_), .Q(cpuregs_24[14]));
DFFcell _34805_ (.C(clk), .D(_01458_), .Q(cpuregs_24[15]));
DFFcell _34806_ (.C(clk), .D(_01459_), .Q(cpuregs_24[16]));
DFFcell _34807_ (.C(clk), .D(_01460_), .Q(cpuregs_24[17]));
DFFcell _34808_ (.C(clk), .D(_01461_), .Q(cpuregs_24[18]));
DFFcell _34809_ (.C(clk), .D(_01462_), .Q(cpuregs_24[19]));
DFFcell _34810_ (.C(clk), .D(_01463_), .Q(cpuregs_24[20]));
DFFcell _34811_ (.C(clk), .D(_01464_), .Q(cpuregs_24[21]));
DFFcell _34812_ (.C(clk), .D(_01465_), .Q(cpuregs_24[22]));
DFFcell _34813_ (.C(clk), .D(_01466_), .Q(cpuregs_24[23]));
DFFcell _34814_ (.C(clk), .D(_01467_), .Q(cpuregs_24[24]));
DFFcell _34815_ (.C(clk), .D(_01468_), .Q(cpuregs_24[25]));
DFFcell _34816_ (.C(clk), .D(_01469_), .Q(cpuregs_24[26]));
DFFcell _34817_ (.C(clk), .D(_01470_), .Q(cpuregs_24[27]));
DFFcell _34818_ (.C(clk), .D(_01471_), .Q(cpuregs_24[28]));
DFFcell _34819_ (.C(clk), .D(_01472_), .Q(cpuregs_24[29]));
DFFcell _34820_ (.C(clk), .D(_01473_), .Q(cpuregs_24[30]));
DFFcell _34821_ (.C(clk), .D(_01474_), .Q(cpuregs_24[31]));
DFFcell _34822_ (.C(clk), .D(_01475_), .Q(cpuregs_2[0]));
DFFcell _34823_ (.C(clk), .D(_01476_), .Q(cpuregs_2[1]));
DFFcell _34824_ (.C(clk), .D(_01477_), .Q(cpuregs_2[2]));
DFFcell _34825_ (.C(clk), .D(_01478_), .Q(cpuregs_2[3]));
DFFcell _34826_ (.C(clk), .D(_01479_), .Q(cpuregs_2[4]));
DFFcell _34827_ (.C(clk), .D(_01480_), .Q(cpuregs_2[5]));
DFFcell _34828_ (.C(clk), .D(_01481_), .Q(cpuregs_2[6]));
DFFcell _34829_ (.C(clk), .D(_01482_), .Q(cpuregs_2[7]));
DFFcell _34830_ (.C(clk), .D(_01483_), .Q(cpuregs_2[8]));
DFFcell _34831_ (.C(clk), .D(_01484_), .Q(cpuregs_2[9]));
DFFcell _34832_ (.C(clk), .D(_01485_), .Q(cpuregs_2[10]));
DFFcell _34833_ (.C(clk), .D(_01486_), .Q(cpuregs_2[11]));
DFFcell _34834_ (.C(clk), .D(_01487_), .Q(cpuregs_2[12]));
DFFcell _34835_ (.C(clk), .D(_01488_), .Q(cpuregs_2[13]));
DFFcell _34836_ (.C(clk), .D(_01489_), .Q(cpuregs_2[14]));
DFFcell _34837_ (.C(clk), .D(_01490_), .Q(cpuregs_2[15]));
DFFcell _34838_ (.C(clk), .D(_01491_), .Q(cpuregs_2[16]));
DFFcell _34839_ (.C(clk), .D(_01492_), .Q(cpuregs_2[17]));
DFFcell _34840_ (.C(clk), .D(_01493_), .Q(cpuregs_2[18]));
DFFcell _34841_ (.C(clk), .D(_01494_), .Q(cpuregs_2[19]));
DFFcell _34842_ (.C(clk), .D(_01495_), .Q(cpuregs_2[20]));
DFFcell _34843_ (.C(clk), .D(_01496_), .Q(cpuregs_2[21]));
DFFcell _34844_ (.C(clk), .D(_01497_), .Q(cpuregs_2[22]));
DFFcell _34845_ (.C(clk), .D(_01498_), .Q(cpuregs_2[23]));
DFFcell _34846_ (.C(clk), .D(_01499_), .Q(cpuregs_2[24]));
DFFcell _34847_ (.C(clk), .D(_01500_), .Q(cpuregs_2[25]));
DFFcell _34848_ (.C(clk), .D(_01501_), .Q(cpuregs_2[26]));
DFFcell _34849_ (.C(clk), .D(_01502_), .Q(cpuregs_2[27]));
DFFcell _34850_ (.C(clk), .D(_01503_), .Q(cpuregs_2[28]));
DFFcell _34851_ (.C(clk), .D(_01504_), .Q(cpuregs_2[29]));
DFFcell _34852_ (.C(clk), .D(_01505_), .Q(cpuregs_2[30]));
DFFcell _34853_ (.C(clk), .D(_01506_), .Q(cpuregs_2[31]));
DFFcell _34854_ (.C(clk), .D(_01507_), .Q(cpuregs_23[0]));
DFFcell _34855_ (.C(clk), .D(_01508_), .Q(cpuregs_23[1]));
DFFcell _34856_ (.C(clk), .D(_01509_), .Q(cpuregs_23[2]));
DFFcell _34857_ (.C(clk), .D(_01510_), .Q(cpuregs_23[3]));
DFFcell _34858_ (.C(clk), .D(_01511_), .Q(cpuregs_23[4]));
DFFcell _34859_ (.C(clk), .D(_01512_), .Q(cpuregs_23[5]));
DFFcell _34860_ (.C(clk), .D(_01513_), .Q(cpuregs_23[6]));
DFFcell _34861_ (.C(clk), .D(_01514_), .Q(cpuregs_23[7]));
DFFcell _34862_ (.C(clk), .D(_01515_), .Q(cpuregs_23[8]));
DFFcell _34863_ (.C(clk), .D(_01516_), .Q(cpuregs_23[9]));
DFFcell _34864_ (.C(clk), .D(_01517_), .Q(cpuregs_23[10]));
DFFcell _34865_ (.C(clk), .D(_01518_), .Q(cpuregs_23[11]));
DFFcell _34866_ (.C(clk), .D(_01519_), .Q(cpuregs_23[12]));
DFFcell _34867_ (.C(clk), .D(_01520_), .Q(cpuregs_23[13]));
DFFcell _34868_ (.C(clk), .D(_01521_), .Q(cpuregs_23[14]));
DFFcell _34869_ (.C(clk), .D(_01522_), .Q(cpuregs_23[15]));
DFFcell _34870_ (.C(clk), .D(_01523_), .Q(cpuregs_23[16]));
DFFcell _34871_ (.C(clk), .D(_01524_), .Q(cpuregs_23[17]));
DFFcell _34872_ (.C(clk), .D(_01525_), .Q(cpuregs_23[18]));
DFFcell _34873_ (.C(clk), .D(_01526_), .Q(cpuregs_23[19]));
DFFcell _34874_ (.C(clk), .D(_01527_), .Q(cpuregs_23[20]));
DFFcell _34875_ (.C(clk), .D(_01528_), .Q(cpuregs_23[21]));
DFFcell _34876_ (.C(clk), .D(_01529_), .Q(cpuregs_23[22]));
DFFcell _34877_ (.C(clk), .D(_01530_), .Q(cpuregs_23[23]));
DFFcell _34878_ (.C(clk), .D(_01531_), .Q(cpuregs_23[24]));
DFFcell _34879_ (.C(clk), .D(_01532_), .Q(cpuregs_23[25]));
DFFcell _34880_ (.C(clk), .D(_01533_), .Q(cpuregs_23[26]));
DFFcell _34881_ (.C(clk), .D(_01534_), .Q(cpuregs_23[27]));
DFFcell _34882_ (.C(clk), .D(_01535_), .Q(cpuregs_23[28]));
DFFcell _34883_ (.C(clk), .D(_01536_), .Q(cpuregs_23[29]));
DFFcell _34884_ (.C(clk), .D(_01537_), .Q(cpuregs_23[30]));
DFFcell _34885_ (.C(clk), .D(_01538_), .Q(cpuregs_23[31]));
DFFcell _34886_ (.C(clk), .D(_01539_), .Q(cpuregs_20[0]));
DFFcell _34887_ (.C(clk), .D(_01540_), .Q(cpuregs_20[1]));
DFFcell _34888_ (.C(clk), .D(_01541_), .Q(cpuregs_20[2]));
DFFcell _34889_ (.C(clk), .D(_01542_), .Q(cpuregs_20[3]));
DFFcell _34890_ (.C(clk), .D(_01543_), .Q(cpuregs_20[4]));
DFFcell _34891_ (.C(clk), .D(_01544_), .Q(cpuregs_20[5]));
DFFcell _34892_ (.C(clk), .D(_01545_), .Q(cpuregs_20[6]));
DFFcell _34893_ (.C(clk), .D(_01546_), .Q(cpuregs_20[7]));
DFFcell _34894_ (.C(clk), .D(_01547_), .Q(cpuregs_20[8]));
DFFcell _34895_ (.C(clk), .D(_01548_), .Q(cpuregs_20[9]));
DFFcell _34896_ (.C(clk), .D(_01549_), .Q(cpuregs_20[10]));
DFFcell _34897_ (.C(clk), .D(_01550_), .Q(cpuregs_20[11]));
DFFcell _34898_ (.C(clk), .D(_01551_), .Q(cpuregs_20[12]));
DFFcell _34899_ (.C(clk), .D(_01552_), .Q(cpuregs_20[13]));
DFFcell _34900_ (.C(clk), .D(_01553_), .Q(cpuregs_20[14]));
DFFcell _34901_ (.C(clk), .D(_01554_), .Q(cpuregs_20[15]));
DFFcell _34902_ (.C(clk), .D(_01555_), .Q(cpuregs_20[16]));
DFFcell _34903_ (.C(clk), .D(_01556_), .Q(cpuregs_20[17]));
DFFcell _34904_ (.C(clk), .D(_01557_), .Q(cpuregs_20[18]));
DFFcell _34905_ (.C(clk), .D(_01558_), .Q(cpuregs_20[19]));
DFFcell _34906_ (.C(clk), .D(_01559_), .Q(cpuregs_20[20]));
DFFcell _34907_ (.C(clk), .D(_01560_), .Q(cpuregs_20[21]));
DFFcell _34908_ (.C(clk), .D(_01561_), .Q(cpuregs_20[22]));
DFFcell _34909_ (.C(clk), .D(_01562_), .Q(cpuregs_20[23]));
DFFcell _34910_ (.C(clk), .D(_01563_), .Q(cpuregs_20[24]));
DFFcell _34911_ (.C(clk), .D(_01564_), .Q(cpuregs_20[25]));
DFFcell _34912_ (.C(clk), .D(_01565_), .Q(cpuregs_20[26]));
DFFcell _34913_ (.C(clk), .D(_01566_), .Q(cpuregs_20[27]));
DFFcell _34914_ (.C(clk), .D(_01567_), .Q(cpuregs_20[28]));
DFFcell _34915_ (.C(clk), .D(_01568_), .Q(cpuregs_20[29]));
DFFcell _34916_ (.C(clk), .D(_01569_), .Q(cpuregs_20[30]));
DFFcell _34917_ (.C(clk), .D(_01570_), .Q(cpuregs_20[31]));
DFFcell _34918_ (.C(clk), .D(_01571_), .Q(cpuregs_19[0]));
DFFcell _34919_ (.C(clk), .D(_01572_), .Q(cpuregs_19[1]));
DFFcell _34920_ (.C(clk), .D(_01573_), .Q(cpuregs_19[2]));
DFFcell _34921_ (.C(clk), .D(_01574_), .Q(cpuregs_19[3]));
DFFcell _34922_ (.C(clk), .D(_01575_), .Q(cpuregs_19[4]));
DFFcell _34923_ (.C(clk), .D(_01576_), .Q(cpuregs_19[5]));
DFFcell _34924_ (.C(clk), .D(_01577_), .Q(cpuregs_19[6]));
DFFcell _34925_ (.C(clk), .D(_01578_), .Q(cpuregs_19[7]));
DFFcell _34926_ (.C(clk), .D(_01579_), .Q(cpuregs_19[8]));
DFFcell _34927_ (.C(clk), .D(_01580_), .Q(cpuregs_19[9]));
DFFcell _34928_ (.C(clk), .D(_01581_), .Q(cpuregs_19[10]));
DFFcell _34929_ (.C(clk), .D(_01582_), .Q(cpuregs_19[11]));
DFFcell _34930_ (.C(clk), .D(_01583_), .Q(cpuregs_19[12]));
DFFcell _34931_ (.C(clk), .D(_01584_), .Q(cpuregs_19[13]));
DFFcell _34932_ (.C(clk), .D(_01585_), .Q(cpuregs_19[14]));
DFFcell _34933_ (.C(clk), .D(_01586_), .Q(cpuregs_19[15]));
DFFcell _34934_ (.C(clk), .D(_01587_), .Q(cpuregs_19[16]));
DFFcell _34935_ (.C(clk), .D(_01588_), .Q(cpuregs_19[17]));
DFFcell _34936_ (.C(clk), .D(_01589_), .Q(cpuregs_19[18]));
DFFcell _34937_ (.C(clk), .D(_01590_), .Q(cpuregs_19[19]));
DFFcell _34938_ (.C(clk), .D(_01591_), .Q(cpuregs_19[20]));
DFFcell _34939_ (.C(clk), .D(_01592_), .Q(cpuregs_19[21]));
DFFcell _34940_ (.C(clk), .D(_01593_), .Q(cpuregs_19[22]));
DFFcell _34941_ (.C(clk), .D(_01594_), .Q(cpuregs_19[23]));
DFFcell _34942_ (.C(clk), .D(_01595_), .Q(cpuregs_19[24]));
DFFcell _34943_ (.C(clk), .D(_01596_), .Q(cpuregs_19[25]));
DFFcell _34944_ (.C(clk), .D(_01597_), .Q(cpuregs_19[26]));
DFFcell _34945_ (.C(clk), .D(_01598_), .Q(cpuregs_19[27]));
DFFcell _34946_ (.C(clk), .D(_01599_), .Q(cpuregs_19[28]));
DFFcell _34947_ (.C(clk), .D(_01600_), .Q(cpuregs_19[29]));
DFFcell _34948_ (.C(clk), .D(_01601_), .Q(cpuregs_19[30]));
DFFcell _34949_ (.C(clk), .D(_01602_), .Q(cpuregs_19[31]));
DFFcell _34950_ (.C(clk), .D(_01603_), .Q(cpuregs_16[0]));
DFFcell _34951_ (.C(clk), .D(_01604_), .Q(cpuregs_16[1]));
DFFcell _34952_ (.C(clk), .D(_01605_), .Q(cpuregs_16[2]));
DFFcell _34953_ (.C(clk), .D(_01606_), .Q(cpuregs_16[3]));
DFFcell _34954_ (.C(clk), .D(_01607_), .Q(cpuregs_16[4]));
DFFcell _34955_ (.C(clk), .D(_01608_), .Q(cpuregs_16[5]));
DFFcell _34956_ (.C(clk), .D(_01609_), .Q(cpuregs_16[6]));
DFFcell _34957_ (.C(clk), .D(_01610_), .Q(cpuregs_16[7]));
DFFcell _34958_ (.C(clk), .D(_01611_), .Q(cpuregs_16[8]));
DFFcell _34959_ (.C(clk), .D(_01612_), .Q(cpuregs_16[9]));
DFFcell _34960_ (.C(clk), .D(_01613_), .Q(cpuregs_16[10]));
DFFcell _34961_ (.C(clk), .D(_01614_), .Q(cpuregs_16[11]));
DFFcell _34962_ (.C(clk), .D(_01615_), .Q(cpuregs_16[12]));
DFFcell _34963_ (.C(clk), .D(_01616_), .Q(cpuregs_16[13]));
DFFcell _34964_ (.C(clk), .D(_01617_), .Q(cpuregs_16[14]));
DFFcell _34965_ (.C(clk), .D(_01618_), .Q(cpuregs_16[15]));
DFFcell _34966_ (.C(clk), .D(_01619_), .Q(cpuregs_16[16]));
DFFcell _34967_ (.C(clk), .D(_01620_), .Q(cpuregs_16[17]));
DFFcell _34968_ (.C(clk), .D(_01621_), .Q(cpuregs_16[18]));
DFFcell _34969_ (.C(clk), .D(_01622_), .Q(cpuregs_16[19]));
DFFcell _34970_ (.C(clk), .D(_01623_), .Q(cpuregs_16[20]));
DFFcell _34971_ (.C(clk), .D(_01624_), .Q(cpuregs_16[21]));
DFFcell _34972_ (.C(clk), .D(_01625_), .Q(cpuregs_16[22]));
DFFcell _34973_ (.C(clk), .D(_01626_), .Q(cpuregs_16[23]));
DFFcell _34974_ (.C(clk), .D(_01627_), .Q(cpuregs_16[24]));
DFFcell _34975_ (.C(clk), .D(_01628_), .Q(cpuregs_16[25]));
DFFcell _34976_ (.C(clk), .D(_01629_), .Q(cpuregs_16[26]));
DFFcell _34977_ (.C(clk), .D(_01630_), .Q(cpuregs_16[27]));
DFFcell _34978_ (.C(clk), .D(_01631_), .Q(cpuregs_16[28]));
DFFcell _34979_ (.C(clk), .D(_01632_), .Q(cpuregs_16[29]));
DFFcell _34980_ (.C(clk), .D(_01633_), .Q(cpuregs_16[30]));
DFFcell _34981_ (.C(clk), .D(_01634_), .Q(cpuregs_16[31]));
DFFcell _34982_ (.C(clk), .D(_01635_), .Q(cpuregs_1[0]));
DFFcell _34983_ (.C(clk), .D(_01636_), .Q(cpuregs_1[1]));
DFFcell _34984_ (.C(clk), .D(_01637_), .Q(cpuregs_1[2]));
DFFcell _34985_ (.C(clk), .D(_01638_), .Q(cpuregs_1[3]));
DFFcell _34986_ (.C(clk), .D(_01639_), .Q(cpuregs_1[4]));
DFFcell _34987_ (.C(clk), .D(_01640_), .Q(cpuregs_1[5]));
DFFcell _34988_ (.C(clk), .D(_01641_), .Q(cpuregs_1[6]));
DFFcell _34989_ (.C(clk), .D(_01642_), .Q(cpuregs_1[7]));
DFFcell _34990_ (.C(clk), .D(_01643_), .Q(cpuregs_1[8]));
DFFcell _34991_ (.C(clk), .D(_01644_), .Q(cpuregs_1[9]));
DFFcell _34992_ (.C(clk), .D(_01645_), .Q(cpuregs_1[10]));
DFFcell _34993_ (.C(clk), .D(_01646_), .Q(cpuregs_1[11]));
DFFcell _34994_ (.C(clk), .D(_01647_), .Q(cpuregs_1[12]));
DFFcell _34995_ (.C(clk), .D(_01648_), .Q(cpuregs_1[13]));
DFFcell _34996_ (.C(clk), .D(_01649_), .Q(cpuregs_1[14]));
DFFcell _34997_ (.C(clk), .D(_01650_), .Q(cpuregs_1[15]));
DFFcell _34998_ (.C(clk), .D(_01651_), .Q(cpuregs_1[16]));
DFFcell _34999_ (.C(clk), .D(_01652_), .Q(cpuregs_1[17]));
DFFcell _35000_ (.C(clk), .D(_01653_), .Q(cpuregs_1[18]));
DFFcell _35001_ (.C(clk), .D(_01654_), .Q(cpuregs_1[19]));
DFFcell _35002_ (.C(clk), .D(_01655_), .Q(cpuregs_1[20]));
DFFcell _35003_ (.C(clk), .D(_01656_), .Q(cpuregs_1[21]));
DFFcell _35004_ (.C(clk), .D(_01657_), .Q(cpuregs_1[22]));
DFFcell _35005_ (.C(clk), .D(_01658_), .Q(cpuregs_1[23]));
DFFcell _35006_ (.C(clk), .D(_01659_), .Q(cpuregs_1[24]));
DFFcell _35007_ (.C(clk), .D(_01660_), .Q(cpuregs_1[25]));
DFFcell _35008_ (.C(clk), .D(_01661_), .Q(cpuregs_1[26]));
DFFcell _35009_ (.C(clk), .D(_01662_), .Q(cpuregs_1[27]));
DFFcell _35010_ (.C(clk), .D(_01663_), .Q(cpuregs_1[28]));
DFFcell _35011_ (.C(clk), .D(_01664_), .Q(cpuregs_1[29]));
DFFcell _35012_ (.C(clk), .D(_01665_), .Q(cpuregs_1[30]));
DFFcell _35013_ (.C(clk), .D(_01666_), .Q(cpuregs_1[31]));
DFFcell _35014_ (.C(clk), .D(_01667_), .Q(cpuregs_10[0]));
DFFcell _35015_ (.C(clk), .D(_01668_), .Q(cpuregs_10[1]));
DFFcell _35016_ (.C(clk), .D(_01669_), .Q(cpuregs_10[2]));
DFFcell _35017_ (.C(clk), .D(_01670_), .Q(cpuregs_10[3]));
DFFcell _35018_ (.C(clk), .D(_01671_), .Q(cpuregs_10[4]));
DFFcell _35019_ (.C(clk), .D(_01672_), .Q(cpuregs_10[5]));
DFFcell _35020_ (.C(clk), .D(_01673_), .Q(cpuregs_10[6]));
DFFcell _35021_ (.C(clk), .D(_01674_), .Q(cpuregs_10[7]));
DFFcell _35022_ (.C(clk), .D(_01675_), .Q(cpuregs_10[8]));
DFFcell _35023_ (.C(clk), .D(_01676_), .Q(cpuregs_10[9]));
DFFcell _35024_ (.C(clk), .D(_01677_), .Q(cpuregs_10[10]));
DFFcell _35025_ (.C(clk), .D(_01678_), .Q(cpuregs_10[11]));
DFFcell _35026_ (.C(clk), .D(_01679_), .Q(cpuregs_10[12]));
DFFcell _35027_ (.C(clk), .D(_01680_), .Q(cpuregs_10[13]));
DFFcell _35028_ (.C(clk), .D(_01681_), .Q(cpuregs_10[14]));
DFFcell _35029_ (.C(clk), .D(_01682_), .Q(cpuregs_10[15]));
DFFcell _35030_ (.C(clk), .D(_01683_), .Q(cpuregs_10[16]));
DFFcell _35031_ (.C(clk), .D(_01684_), .Q(cpuregs_10[17]));
DFFcell _35032_ (.C(clk), .D(_01685_), .Q(cpuregs_10[18]));
DFFcell _35033_ (.C(clk), .D(_01686_), .Q(cpuregs_10[19]));
DFFcell _35034_ (.C(clk), .D(_01687_), .Q(cpuregs_10[20]));
DFFcell _35035_ (.C(clk), .D(_01688_), .Q(cpuregs_10[21]));
DFFcell _35036_ (.C(clk), .D(_01689_), .Q(cpuregs_10[22]));
DFFcell _35037_ (.C(clk), .D(_01690_), .Q(cpuregs_10[23]));
DFFcell _35038_ (.C(clk), .D(_01691_), .Q(cpuregs_10[24]));
DFFcell _35039_ (.C(clk), .D(_01692_), .Q(cpuregs_10[25]));
DFFcell _35040_ (.C(clk), .D(_01693_), .Q(cpuregs_10[26]));
DFFcell _35041_ (.C(clk), .D(_01694_), .Q(cpuregs_10[27]));
DFFcell _35042_ (.C(clk), .D(_01695_), .Q(cpuregs_10[28]));
DFFcell _35043_ (.C(clk), .D(_01696_), .Q(cpuregs_10[29]));
DFFcell _35044_ (.C(clk), .D(_01697_), .Q(cpuregs_10[30]));
DFFcell _35045_ (.C(clk), .D(_01698_), .Q(cpuregs_10[31]));
assign eoi = 32'd0;
assign pcpi_insn = 32'hxxxxxxxx;
assign pcpi_valid = 1'h0;
assign trace_data = 36'hxxxxxxxxx;
assign trace_valid = 1'h0;
endmodule
