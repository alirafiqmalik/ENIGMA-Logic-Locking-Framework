module locked(inputA, inputB, out);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
wire _28_;
input [7:0] inputA;
wire [7:0] inputA;
input [7:0] inputB;
wire [7:0] inputB;
output [8:0] out;
wire [8:0] out;
NAND_g _29_ ( .A(inputA[7]), .B(inputB[7]), .Y(_00_) );
NOR_g _30_ ( .A(inputA[7]), .B(inputB[7]), .Y(_01_) );
NAND_g _31_ ( .A(inputA[6]), .B(inputB[6]), .Y(_02_) );
XOR_g _32_ ( .A(inputA[6]), .B(inputB[6]), .Y(_03_) );
NAND_g _33_ ( .A(inputA[5]), .B(inputB[5]), .Y(_04_) );
NAND_g _34_ ( .A(inputA[4]), .B(inputB[4]), .Y(_05_) );
NAND_g _35_ ( .A(inputA[3]), .B(inputB[3]), .Y(_06_) );
NAND_g _36_ ( .A(inputA[2]), .B(inputB[2]), .Y(_07_) );
NAND_g _37_ ( .A(inputA[1]), .B(inputB[1]), .Y(_08_) );
AND_g _38_ ( .A(inputA[0]), .B(inputB[0]), .Y(_09_) );
XOR_g _39_ ( .A(inputA[1]), .B(inputB[1]), .Y(_10_) );
NAND_g _40_ ( .A(_09_), .B(_10_), .Y(_11_) );
NAND_g _41_ ( .A(_08_), .B(_11_), .Y(_12_) );
XOR_g _42_ ( .A(inputA[2]), .B(inputB[2]), .Y(_13_) );
NAND_g _43_ ( .A(_12_), .B(_13_), .Y(_14_) );
NAND_g _44_ ( .A(_07_), .B(_14_), .Y(_15_) );
XOR_g _45_ ( .A(inputA[3]), .B(inputB[3]), .Y(_16_) );
NAND_g _46_ ( .A(_15_), .B(_16_), .Y(_17_) );
NAND_g _47_ ( .A(_06_), .B(_17_), .Y(_18_) );
XOR_g _48_ ( .A(inputA[4]), .B(inputB[4]), .Y(_19_) );
NAND_g _49_ ( .A(_18_), .B(_19_), .Y(_20_) );
NAND_g _50_ ( .A(_05_), .B(_20_), .Y(_21_) );
XOR_g _51_ ( .A(inputA[5]), .B(inputB[5]), .Y(_22_) );
NAND_g _52_ ( .A(_21_), .B(_22_), .Y(_23_) );
NAND_g _53_ ( .A(_04_), .B(_23_), .Y(_24_) );
NAND_g _54_ ( .A(_03_), .B(_24_), .Y(_25_) );
AND_g _55_ ( .A(_02_), .B(_25_), .Y(_26_) );
AND_g _56_ ( .A(_00_), .B(_26_), .Y(_27_) );
NOR_g _57_ ( .A(_01_), .B(_27_), .Y(out[8]) );
XOR_g _58_ ( .A(_09_), .B(_10_), .Y(out[1]) );
XOR_g _59_ ( .A(_12_), .B(_13_), .Y(out[2]) );
XOR_g _60_ ( .A(_15_), .B(_16_), .Y(out[3]) );
XOR_g _61_ ( .A(_18_), .B(_19_), .Y(out[4]) );
XOR_g _62_ ( .A(_21_), .B(_22_), .Y(out[5]) );
XOR_g _63_ ( .A(_03_), .B(_24_), .Y(out[6]) );
XOR_g _64_ ( .A(inputA[7]), .B(inputB[7]), .Y(_28_) );
XNOR_g _65_ ( .A(_26_), .B(_28_), .Y(out[7]) );
XOR_g _66_ ( .A(inputA[0]), .B(inputB[0]), .Y(out[0]) );
endmodule
