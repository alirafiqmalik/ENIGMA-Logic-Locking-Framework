module top(CLOCK_50, KEY_N, SW, vga_x, vga_y, vga_plot, vga_colour);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  input CLOCK_50;
  wire CLOCK_50;
  input [3:0] KEY_N;
  wire [3:0] KEY_N;
  input [9:0] SW;
  wire [9:0] SW;
  wire T2Done;
  wire [2:0] T2colour;
  wire T2plot;
  wire [7:0] T2x;
  wire [6:0] T2y;
  wire [2:0] T3colourcircle;
  wire [8:0] T3d;
  wire T3plot;
  wire [3:0] T3state;
  wire [7:0] T3x;
  wire [7:0] T3xp;
  wire [6:0] T3y;
  wire [6:0] T3yp;
  output [2:0] vga_colour;
  wire [2:0] vga_colour;
  output vga_plot;
  wire vga_plot;
  output [7:0] vga_x;
  wire [7:0] vga_x;
  output [6:0] vga_y;
  wire [6:0] vga_y;
  NOT_g _1038_ ( .A(T2Done), .Y(_0011_));
  NAND_g _1039_ ( .A(T3colourcircle[0]), .B(T2Done), .Y(_0012_));
  NAND_g _1040_ ( .A(T2colour[0]), .B(_0011_), .Y(_0013_));
  NAND_g _1041_ ( .A(_0012_), .B(_0013_), .Y(vga_colour[0]));
  NAND_g _1042_ ( .A(T2Done), .B(T3colourcircle[1]), .Y(_0014_));
  NAND_g _1043_ ( .A(_0011_), .B(T2colour[1]), .Y(_0015_));
  NAND_g _1044_ ( .A(_0014_), .B(_0015_), .Y(vga_colour[1]));
  NAND_g _1045_ ( .A(T2Done), .B(T3colourcircle[2]), .Y(_0016_));
  NAND_g _1046_ ( .A(_0011_), .B(T2colour[2]), .Y(_0017_));
  NAND_g _1047_ ( .A(_0016_), .B(_0017_), .Y(vga_colour[2]));
  NAND_g _1048_ ( .A(T2Done), .B(T3plot), .Y(_0018_));
  NAND_g _1049_ ( .A(_0011_), .B(T2plot), .Y(_0019_));
  NAND_g _1050_ ( .A(_0018_), .B(_0019_), .Y(vga_plot));
  NAND_g _1051_ ( .A(T2Done), .B(T3yp[0]), .Y(_0020_));
  NAND_g _1052_ ( .A(_0011_), .B(T2y[0]), .Y(_0021_));
  NAND_g _1053_ ( .A(_0020_), .B(_0021_), .Y(vga_y[0]));
  NAND_g _1054_ ( .A(T2Done), .B(T3yp[1]), .Y(_0022_));
  NAND_g _1055_ ( .A(_0011_), .B(T2y[1]), .Y(_0023_));
  NAND_g _1056_ ( .A(_0022_), .B(_0023_), .Y(vga_y[1]));
  NAND_g _1057_ ( .A(T2Done), .B(T3yp[2]), .Y(_0024_));
  NAND_g _1058_ ( .A(_0011_), .B(T2y[2]), .Y(_0025_));
  NAND_g _1059_ ( .A(_0024_), .B(_0025_), .Y(vga_y[2]));
  NAND_g _1060_ ( .A(T2Done), .B(T3yp[3]), .Y(_0026_));
  NAND_g _1061_ ( .A(_0011_), .B(T2y[3]), .Y(_0027_));
  NAND_g _1062_ ( .A(_0026_), .B(_0027_), .Y(vga_y[3]));
  NAND_g _1063_ ( .A(T2Done), .B(T3yp[4]), .Y(_0028_));
  NAND_g _1064_ ( .A(_0011_), .B(T2y[4]), .Y(_0029_));
  NAND_g _1065_ ( .A(_0028_), .B(_0029_), .Y(vga_y[4]));
  NAND_g _1066_ ( .A(T2Done), .B(T3yp[5]), .Y(_0030_));
  NAND_g _1067_ ( .A(_0011_), .B(T2y[5]), .Y(_0031_));
  NAND_g _1068_ ( .A(_0030_), .B(_0031_), .Y(vga_y[5]));
  NAND_g _1069_ ( .A(T2Done), .B(T3yp[6]), .Y(_0032_));
  NAND_g _1070_ ( .A(_0011_), .B(T2y[6]), .Y(_0033_));
  NAND_g _1071_ ( .A(_0032_), .B(_0033_), .Y(vga_y[6]));
  NAND_g _1072_ ( .A(T2Done), .B(T3xp[0]), .Y(_0034_));
  NAND_g _1073_ ( .A(_0011_), .B(T2x[0]), .Y(_0035_));
  NAND_g _1074_ ( .A(_0034_), .B(_0035_), .Y(vga_x[0]));
  NAND_g _1075_ ( .A(T2Done), .B(T3xp[1]), .Y(_0036_));
  NAND_g _1076_ ( .A(_0011_), .B(T2x[1]), .Y(_0037_));
  NAND_g _1077_ ( .A(_0036_), .B(_0037_), .Y(vga_x[1]));
  NAND_g _1078_ ( .A(T2Done), .B(T3xp[2]), .Y(_0038_));
  NAND_g _1079_ ( .A(_0011_), .B(T2x[2]), .Y(_0000_));
  NAND_g _1080_ ( .A(_0038_), .B(_0000_), .Y(vga_x[2]));
  NAND_g _1081_ ( .A(T2Done), .B(T3xp[3]), .Y(_0001_));
  NAND_g _1082_ ( .A(_0011_), .B(T2x[3]), .Y(_0002_));
  NAND_g _1083_ ( .A(_0001_), .B(_0002_), .Y(vga_x[3]));
  NAND_g _1084_ ( .A(T2Done), .B(T3xp[4]), .Y(_0003_));
  NAND_g _1085_ ( .A(_0011_), .B(T2x[4]), .Y(_0004_));
  NAND_g _1086_ ( .A(_0003_), .B(_0004_), .Y(vga_x[4]));
  NAND_g _1087_ ( .A(T2Done), .B(T3xp[5]), .Y(_0005_));
  NAND_g _1088_ ( .A(_0011_), .B(T2x[5]), .Y(_0006_));
  NAND_g _1089_ ( .A(_0005_), .B(_0006_), .Y(vga_x[5]));
  NAND_g _1090_ ( .A(T2Done), .B(T3xp[6]), .Y(_0007_));
  NAND_g _1091_ ( .A(_0011_), .B(T2x[6]), .Y(_0008_));
  NAND_g _1092_ ( .A(_0007_), .B(_0008_), .Y(vga_x[6]));
  NAND_g _1093_ ( .A(T2Done), .B(T3xp[7]), .Y(_0009_));
  NAND_g _1094_ ( .A(_0011_), .B(T2x[7]), .Y(_0010_));
  NAND_g _1095_ ( .A(_0009_), .B(_0010_), .Y(vga_x[7]));
  NOT_g _1096_ ( .A(T2y[0]), .Y(_0113_));
  NOT_g _1097_ ( .A(_0039_), .Y(T2plot));
  NOT_g _1098_ ( .A(T2x[7]), .Y(_0114_));
  NOT_g _1099_ ( .A(T2x[6]), .Y(_0115_));
  NOT_g _1100_ ( .A(KEY_N[3]), .Y(_0040_));
  AND_g _1101_ ( .A(T2x[1]), .B(T2x[0]), .Y(_0116_));
  AND_g _1102_ ( .A(T2x[2]), .B(_0116_), .Y(_0117_));
  AND_g _1103_ ( .A(T2x[3]), .B(_0117_), .Y(_0118_));
  AND_g _1104_ ( .A(T2x[4]), .B(_0118_), .Y(_0119_));
  NOR_g _1105_ ( .A(T2x[6]), .B(T2x[5]), .Y(_0120_));
  AND_g _1106_ ( .A(T2x[7]), .B(_0120_), .Y(_0121_));
  AND_g _1107_ ( .A(_0119_), .B(_0121_), .Y(_0122_));
  NAND_g _1108_ ( .A(_0119_), .B(_0121_), .Y(_0123_));
  AND_g _1109_ ( .A(T2y[1]), .B(T2y[0]), .Y(_0124_));
  AND_g _1110_ ( .A(T2y[2]), .B(_0124_), .Y(_0125_));
  AND_g _1111_ ( .A(T2y[6]), .B(T2y[5]), .Y(_0126_));
  NAND_g _1112_ ( .A(T2y[4]), .B(_0126_), .Y(_0127_));
  NOR_g _1113_ ( .A(T2y[3]), .B(_0127_), .Y(_0128_));
  AND_g _1114_ ( .A(_0125_), .B(_0128_), .Y(_0129_));
  NAND_g _1115_ ( .A(_0122_), .B(_0129_), .Y(_0130_));
  NAND_g _1116_ ( .A(T2plot), .B(_0130_), .Y(_0071_));
  NOR_g _1117_ ( .A(T2y[3]), .B(_0125_), .Y(_0131_));
  NOR_g _1118_ ( .A(_0127_), .B(_0131_), .Y(_0132_));
  NOR_g _1119_ ( .A(_0123_), .B(_0132_), .Y(_0133_));
  AND_g _1120_ ( .A(T2y[3]), .B(_0125_), .Y(_0134_));
  AND_g _1121_ ( .A(T2y[4]), .B(_0134_), .Y(_0135_));
  AND_g _1122_ ( .A(T2y[5]), .B(_0135_), .Y(_0136_));
  NOR_g _1123_ ( .A(T2x[5]), .B(_0119_), .Y(_0137_));
  NAND_g _1124_ ( .A(_0115_), .B(_0137_), .Y(_0138_));
  AND_g _1125_ ( .A(T2x[7]), .B(_0138_), .Y(_0139_));
  NAND_g _1126_ ( .A(T2x[7]), .B(_0138_), .Y(_0140_));
  NAND_g _1127_ ( .A(_0130_), .B(_0139_), .Y(_0141_));
  AND_g _1128_ ( .A(_0133_), .B(_0136_), .Y(_0142_));
  NOR_g _1129_ ( .A(T2y[6]), .B(_0142_), .Y(_0143_));
  NOR_g _1130_ ( .A(_0133_), .B(_0141_), .Y(_0144_));
  NOR_g _1131_ ( .A(_0143_), .B(_0144_), .Y(_0070_));
  NAND_g _1132_ ( .A(T2y[5]), .B(_0141_), .Y(_0145_));
  XOR_g _1133_ ( .A(T2y[5]), .B(_0135_), .Y(_0146_));
  NAND_g _1134_ ( .A(_0133_), .B(_0146_), .Y(_0147_));
  NAND_g _1135_ ( .A(_0145_), .B(_0147_), .Y(_0069_));
  NAND_g _1136_ ( .A(T2y[4]), .B(_0141_), .Y(_0148_));
  XOR_g _1137_ ( .A(T2y[4]), .B(_0134_), .Y(_0075_));
  NAND_g _1138_ ( .A(_0133_), .B(_0075_), .Y(_0076_));
  NAND_g _1139_ ( .A(_0148_), .B(_0076_), .Y(_0068_));
  NAND_g _1140_ ( .A(T2y[3]), .B(_0140_), .Y(_0077_));
  XOR_g _1141_ ( .A(T2y[3]), .B(_0125_), .Y(_0078_));
  NAND_g _1142_ ( .A(_0133_), .B(_0078_), .Y(_0079_));
  NAND_g _1143_ ( .A(_0077_), .B(_0079_), .Y(_0067_));
  NAND_g _1144_ ( .A(T2y[2]), .B(_0141_), .Y(_0080_));
  XOR_g _1145_ ( .A(T2y[2]), .B(_0124_), .Y(_0081_));
  NAND_g _1146_ ( .A(_0133_), .B(_0081_), .Y(_0082_));
  NAND_g _1147_ ( .A(_0080_), .B(_0082_), .Y(_0066_));
  NAND_g _1148_ ( .A(T2y[1]), .B(_0141_), .Y(_0083_));
  XOR_g _1149_ ( .A(T2y[1]), .B(T2y[0]), .Y(_0084_));
  NAND_g _1150_ ( .A(_0133_), .B(_0084_), .Y(_0085_));
  NAND_g _1151_ ( .A(_0083_), .B(_0085_), .Y(_0065_));
  NAND_g _1152_ ( .A(_0113_), .B(_0133_), .Y(_0086_));
  NAND_g _1153_ ( .A(T2y[0]), .B(_0141_), .Y(_0087_));
  NAND_g _1154_ ( .A(_0086_), .B(_0087_), .Y(_0064_));
  AND_g _1155_ ( .A(T2x[5]), .B(_0119_), .Y(_0088_));
  NOT_g _1156_ ( .A(_0088_), .Y(_0089_));
  NAND_g _1157_ ( .A(T2x[6]), .B(_0088_), .Y(_0090_));
  NAND_g _1158_ ( .A(_0114_), .B(_0090_), .Y(_0091_));
  AND_g _1159_ ( .A(_0141_), .B(_0091_), .Y(_0063_));
  NOR_g _1160_ ( .A(T2x[6]), .B(_0088_), .Y(_0092_));
  NOR_g _1161_ ( .A(_0091_), .B(_0092_), .Y(_0062_));
  NOR_g _1162_ ( .A(T2x[7]), .B(_0137_), .Y(_0093_));
  AND_g _1163_ ( .A(_0089_), .B(_0093_), .Y(_0061_));
  XOR_g _1164_ ( .A(T2x[4]), .B(_0118_), .Y(_0094_));
  NAND_g _1165_ ( .A(_0140_), .B(_0094_), .Y(_0095_));
  NAND_g _1166_ ( .A(_0130_), .B(_0095_), .Y(_0060_));
  XOR_g _1167_ ( .A(T2x[3]), .B(_0117_), .Y(_0096_));
  NAND_g _1168_ ( .A(_0140_), .B(_0096_), .Y(_0097_));
  NAND_g _1169_ ( .A(_0130_), .B(_0097_), .Y(_0059_));
  XOR_g _1170_ ( .A(T2x[2]), .B(_0116_), .Y(_0098_));
  NAND_g _1171_ ( .A(_0140_), .B(_0098_), .Y(_0099_));
  NAND_g _1172_ ( .A(_0130_), .B(_0099_), .Y(_0058_));
  XOR_g _1173_ ( .A(T2x[1]), .B(T2x[0]), .Y(_0100_));
  NAND_g _1174_ ( .A(_0140_), .B(_0100_), .Y(_0101_));
  NAND_g _1175_ ( .A(_0130_), .B(_0101_), .Y(_0057_));
  NAND_g _1176_ ( .A(T2x[0]), .B(_0130_), .Y(_0102_));
  AND_g _1177_ ( .A(_0141_), .B(_0102_), .Y(_0056_));
  AND_g _1178_ ( .A(KEY_N[3]), .B(_0140_), .Y(_0103_));
  NAND_g _1179_ ( .A(SW[9]), .B(T2y[0]), .Y(_0104_));
  AND_g _1180_ ( .A(_0103_), .B(_0104_), .Y(_0105_));
  NOR_g _1181_ ( .A(T2colour[0]), .B(_0103_), .Y(_0106_));
  NOR_g _1182_ ( .A(_0105_), .B(_0106_), .Y(_0072_));
  NAND_g _1183_ ( .A(SW[9]), .B(T2y[1]), .Y(_0107_));
  AND_g _1184_ ( .A(_0103_), .B(_0107_), .Y(_0108_));
  NOR_g _1185_ ( .A(T2colour[1]), .B(_0103_), .Y(_0109_));
  NOR_g _1186_ ( .A(_0108_), .B(_0109_), .Y(_0073_));
  NAND_g _1187_ ( .A(T2y[2]), .B(SW[9]), .Y(_0110_));
  AND_g _1188_ ( .A(_0103_), .B(_0110_), .Y(_0111_));
  NOR_g _1189_ ( .A(T2colour[2]), .B(_0103_), .Y(_0112_));
  NOR_g _1190_ ( .A(_0111_), .B(_0112_), .Y(_0074_));
  NOT_g _1191_ ( .A(KEY_N[3]), .Y(_0041_));
  NOT_g _1192_ ( .A(KEY_N[3]), .Y(_0042_));
  NOT_g _1193_ ( .A(KEY_N[3]), .Y(_0043_));
  NOT_g _1194_ ( .A(KEY_N[3]), .Y(_0044_));
  NOT_g _1195_ ( .A(KEY_N[3]), .Y(_0045_));
  NOT_g _1196_ ( .A(KEY_N[3]), .Y(_0046_));
  NOT_g _1197_ ( .A(KEY_N[3]), .Y(_0047_));
  NOT_g _1198_ ( .A(KEY_N[3]), .Y(_0048_));
  NOT_g _1199_ ( .A(KEY_N[3]), .Y(_0049_));
  NOT_g _1200_ ( .A(KEY_N[3]), .Y(_0050_));
  NOT_g _1201_ ( .A(KEY_N[3]), .Y(_0051_));
  NOT_g _1202_ ( .A(KEY_N[3]), .Y(_0052_));
  NOT_g _1203_ ( .A(KEY_N[3]), .Y(_0053_));
  NOT_g _1204_ ( .A(KEY_N[3]), .Y(_0054_));
  NOT_g _1205_ ( .A(KEY_N[3]), .Y(_0055_));
  BUF_g _1206_ ( .A(_0039_), .Y(T2Done));
  DFFRcell _1207_ ( .C(CLOCK_50), .D(_0056_), .Q(T2x[0]), .R(_0040_));
  DFFRcell _1208_ ( .C(CLOCK_50), .D(_0057_), .Q(T2x[1]), .R(_0041_));
  DFFRcell _1209_ ( .C(CLOCK_50), .D(_0058_), .Q(T2x[2]), .R(_0042_));
  DFFRcell _1210_ ( .C(CLOCK_50), .D(_0059_), .Q(T2x[3]), .R(_0043_));
  DFFRcell _1211_ ( .C(CLOCK_50), .D(_0060_), .Q(T2x[4]), .R(_0044_));
  DFFRcell _1212_ ( .C(CLOCK_50), .D(_0061_), .Q(T2x[5]), .R(_0045_));
  DFFRcell _1213_ ( .C(CLOCK_50), .D(_0062_), .Q(T2x[6]), .R(_0046_));
  DFFRcell _1214_ ( .C(CLOCK_50), .D(_0063_), .Q(T2x[7]), .R(_0047_));
  DFFRcell _1215_ ( .C(CLOCK_50), .D(_0064_), .Q(T2y[0]), .R(_0048_));
  DFFRcell _1216_ ( .C(CLOCK_50), .D(_0065_), .Q(T2y[1]), .R(_0049_));
  DFFRcell _1217_ ( .C(CLOCK_50), .D(_0066_), .Q(T2y[2]), .R(_0050_));
  DFFRcell _1218_ ( .C(CLOCK_50), .D(_0067_), .Q(T2y[3]), .R(_0051_));
  DFFRcell _1219_ ( .C(CLOCK_50), .D(_0068_), .Q(T2y[4]), .R(_0052_));
  DFFRcell _1220_ ( .C(CLOCK_50), .D(_0069_), .Q(T2y[5]), .R(_0053_));
  DFFRcell _1221_ ( .C(CLOCK_50), .D(_0070_), .Q(T2y[6]), .R(_0054_));
  DFFRcell _1222_ ( .C(CLOCK_50), .D(_0071_), .Q(_0039_), .R(_0055_));
  DFFcell _1223_ ( .C(CLOCK_50), .D(_0072_), .Q(T2colour[0]));
  DFFcell _1224_ ( .C(CLOCK_50), .D(_0073_), .Q(T2colour[1]));
  DFFcell _1225_ ( .C(CLOCK_50), .D(_0074_), .Q(T2colour[2]));
  NOT_g _1226_ ( .A(T3state[3]), .Y(_0210_));
  NOT_g _1227_ ( .A(T3state[2]), .Y(_0211_));
  NOT_g _1228_ ( .A(T3state[0]), .Y(_0212_));
  NOT_g _1229_ ( .A(KEY_N[3]), .Y(_0149_));
  NOT_g _1230_ ( .A(T3y[0]), .Y(_0213_));
  NOT_g _1231_ ( .A(T3y[1]), .Y(_0214_));
  NOT_g _1232_ ( .A(T3y[2]), .Y(_0215_));
  NOT_g _1233_ ( .A(T3y[3]), .Y(_0216_));
  NOT_g _1234_ ( .A(T3y[4]), .Y(_0217_));
  NOT_g _1235_ ( .A(T3y[5]), .Y(_0218_));
  NOT_g _1236_ ( .A(T3y[6]), .Y(_0219_));
  NOT_g _1237_ ( .A(T3d[1]), .Y(_0220_));
  NOT_g _1238_ ( .A(T3x[0]), .Y(_0221_));
  NOT_g _1239_ ( .A(T3x[1]), .Y(_0222_));
  NOT_g _1240_ ( .A(T3x[2]), .Y(_0223_));
  NOT_g _1241_ ( .A(T3x[3]), .Y(_0224_));
  NOT_g _1242_ ( .A(T3x[4]), .Y(_0225_));
  NOT_g _1243_ ( .A(T3x[5]), .Y(_0226_));
  NOT_g _1244_ ( .A(T3x[6]), .Y(_0227_));
  NOT_g _1245_ ( .A(SW[3]), .Y(_0228_));
  NOT_g _1246_ ( .A(SW[4]), .Y(_0229_));
  NOT_g _1247_ ( .A(1'h1), .Y(_0230_));
  NOT_g _1248_ ( .A(1'h1), .Y(_0231_));
  NOT_g _1249_ ( .A(1'h0), .Y(_0232_));
  NOT_g _1250_ ( .A(1'h1), .Y(_0233_));
  NOT_g _1251_ ( .A(1'h1), .Y(_0234_));
  NOT_g _1252_ ( .A(1'h1), .Y(_0235_));
  NOR_g _1253_ ( .A(T3state[1]), .B(T3state[0]), .Y(_0236_));
  AND_g _1254_ ( .A(_0211_), .B(_0236_), .Y(_0237_));
  NAND_g _1255_ ( .A(_0211_), .B(_0236_), .Y(_0238_));
  AND_g _1256_ ( .A(T3state[3]), .B(_0238_), .Y(_0239_));
  NAND_g _1257_ ( .A(T3state[3]), .B(_0238_), .Y(_0240_));
  AND_g _1258_ ( .A(T2Done), .B(_0240_), .Y(_0241_));
  NAND_g _1259_ ( .A(T2Done), .B(_0240_), .Y(_0242_));
  NOR_g _1260_ ( .A(T3y[0]), .B(T3y[1]), .Y(_0243_));
  NAND_g _1261_ ( .A(_0215_), .B(_0243_), .Y(_0244_));
  NOT_g _1262_ ( .A(_0244_), .Y(_0245_));
  NOR_g _1263_ ( .A(T3y[3]), .B(_0244_), .Y(_0246_));
  AND_g _1264_ ( .A(_0217_), .B(_0246_), .Y(_0247_));
  NAND_g _1265_ ( .A(_0218_), .B(_0247_), .Y(_0248_));
  NOT_g _1266_ ( .A(_0248_), .Y(_0249_));
  NOR_g _1267_ ( .A(T3y[6]), .B(_0248_), .Y(_0250_));
  AND_g _1268_ ( .A(_0210_), .B(T3state[2]), .Y(_0251_));
  AND_g _1269_ ( .A(T3state[0]), .B(_0251_), .Y(_0252_));
  NOT_g _1270_ ( .A(_0252_), .Y(_0253_));
  NAND_g _1271_ ( .A(T3state[1]), .B(_0252_), .Y(_0254_));
  NOR_g _1272_ ( .A(_0250_), .B(_0254_), .Y(_0255_));
  NOR_g _1273_ ( .A(_0242_), .B(_0255_), .Y(_0256_));
  NOR_g _1274_ ( .A(T3state[3]), .B(T2Done), .Y(_0257_));
  NOR_g _1275_ ( .A(_0256_), .B(_0257_), .Y(_0156_));
  NAND_g _1276_ ( .A(_0236_), .B(_0251_), .Y(_0258_));
  NOR_g _1277_ ( .A(T3state[3]), .B(T3state[2]), .Y(_0259_));
  AND_g _1278_ ( .A(T3state[0]), .B(_0259_), .Y(_0260_));
  NAND_g _1279_ ( .A(T3state[1]), .B(_0260_), .Y(_0261_));
  NAND_g _1280_ ( .A(_0258_), .B(_0261_), .Y(_0262_));
  AND_g _1281_ ( .A(T3state[1]), .B(_0212_), .Y(_0263_));
  XOR_g _1282_ ( .A(T3state[1]), .B(T3state[0]), .Y(_0264_));
  AND_g _1283_ ( .A(_0251_), .B(_0264_), .Y(_0265_));
  NOR_g _1284_ ( .A(_0262_), .B(_0265_), .Y(_0266_));
  NAND_g _1285_ ( .A(_0211_), .B(_0242_), .Y(_0267_));
  NAND_g _1286_ ( .A(_0241_), .B(_0266_), .Y(_0268_));
  AND_g _1287_ ( .A(_0267_), .B(_0268_), .Y(_0155_));
  NAND_g _1288_ ( .A(T3state[1]), .B(_0242_), .Y(_0269_));
  AND_g _1289_ ( .A(T2Done), .B(_0264_), .Y(_0270_));
  NAND_g _1290_ ( .A(_0210_), .B(_0270_), .Y(_0271_));
  NAND_g _1291_ ( .A(_0269_), .B(_0271_), .Y(_0154_));
  NAND_g _1292_ ( .A(T3y[6]), .B(_0227_), .Y(_0272_));
  NAND_g _1293_ ( .A(_0218_), .B(T3x[5]), .Y(_0273_));
  NAND_g _1294_ ( .A(T3y[3]), .B(_0224_), .Y(_0274_));
  NAND_g _1295_ ( .A(_0215_), .B(T3x[2]), .Y(_0275_));
  NAND_g _1296_ ( .A(_0214_), .B(T3x[1]), .Y(_0276_));
  NAND_g _1297_ ( .A(_0213_), .B(T3x[0]), .Y(_0277_));
  NAND_g _1298_ ( .A(_0276_), .B(_0277_), .Y(_0278_));
  NAND_g _1299_ ( .A(T3y[1]), .B(_0222_), .Y(_0279_));
  NAND_g _1300_ ( .A(T3y[2]), .B(_0223_), .Y(_0280_));
  AND_g _1301_ ( .A(_0279_), .B(_0280_), .Y(_0281_));
  NAND_g _1302_ ( .A(_0278_), .B(_0281_), .Y(_0282_));
  NAND_g _1303_ ( .A(_0275_), .B(_0282_), .Y(_0283_));
  NAND_g _1304_ ( .A(_0274_), .B(_0283_), .Y(_0284_));
  NAND_g _1305_ ( .A(_0217_), .B(T3x[4]), .Y(_0285_));
  NAND_g _1306_ ( .A(_0216_), .B(T3x[3]), .Y(_0286_));
  AND_g _1307_ ( .A(_0285_), .B(_0286_), .Y(_0287_));
  NAND_g _1308_ ( .A(_0284_), .B(_0287_), .Y(_0288_));
  NAND_g _1309_ ( .A(T3y[5]), .B(_0226_), .Y(_0289_));
  NAND_g _1310_ ( .A(T3y[4]), .B(_0225_), .Y(_0290_));
  AND_g _1311_ ( .A(_0289_), .B(_0290_), .Y(_0291_));
  NAND_g _1312_ ( .A(_0288_), .B(_0291_), .Y(_0292_));
  NAND_g _1313_ ( .A(_0273_), .B(_0292_), .Y(_0293_));
  NAND_g _1314_ ( .A(_0272_), .B(_0293_), .Y(_0294_));
  AND_g _1315_ ( .A(T3state[3]), .B(_0237_), .Y(_0295_));
  NAND_g _1316_ ( .A(T3state[3]), .B(_0237_), .Y(_0296_));
  NOR_g _1317_ ( .A(T3x[7]), .B(_0296_), .Y(_0297_));
  NAND_g _1318_ ( .A(_0219_), .B(T3x[6]), .Y(_0298_));
  AND_g _1319_ ( .A(_0297_), .B(_0298_), .Y(_0299_));
  NAND_g _1320_ ( .A(_0294_), .B(_0299_), .Y(_0300_));
  AND_g _1321_ ( .A(_0236_), .B(_0259_), .Y(_0301_));
  NOT_g _1322_ ( .A(_0301_), .Y(T3plot));
  NOR_g _1323_ ( .A(KEY_N[0]), .B(T3plot), .Y(_0302_));
  NAND_g _1324_ ( .A(_0251_), .B(_0263_), .Y(_0303_));
  NAND_g _1325_ ( .A(_0259_), .B(_0263_), .Y(_0304_));
  NAND_g _1326_ ( .A(_0258_), .B(_0304_), .Y(_0305_));
  NOR_g _1327_ ( .A(_0302_), .B(_0305_), .Y(_0306_));
  AND_g _1328_ ( .A(_0303_), .B(_0306_), .Y(_0307_));
  NAND_g _1329_ ( .A(_0300_), .B(_0307_), .Y(_0308_));
  NAND_g _1330_ ( .A(_0241_), .B(_0308_), .Y(_0309_));
  NAND_g _1331_ ( .A(T3state[0]), .B(_0242_), .Y(_0310_));
  NAND_g _1332_ ( .A(_0309_), .B(_0310_), .Y(_0153_));
  NOR_g _1333_ ( .A(T3d[4]), .B(T3d[5]), .Y(_0311_));
  NOR_g _1334_ ( .A(T3d[6]), .B(T3d[7]), .Y(_0312_));
  AND_g _1335_ ( .A(_0311_), .B(_0312_), .Y(_0313_));
  NOR_g _1336_ ( .A(T3d[2]), .B(T3d[3]), .Y(_0314_));
  NOR_g _1337_ ( .A(T3d[0]), .B(T3d[1]), .Y(_0315_));
  AND_g _1338_ ( .A(_0314_), .B(_0315_), .Y(_0316_));
  NAND_g _1339_ ( .A(_0313_), .B(_0316_), .Y(_0317_));
  NAND_g _1340_ ( .A(T3d[8]), .B(_0317_), .Y(_0318_));
  NOT_g _1341_ ( .A(_0318_), .Y(_0319_));
  AND_g _1342_ ( .A(_0237_), .B(_0318_), .Y(_0320_));
  NOR_g _1343_ ( .A(_0301_), .B(_0320_), .Y(_0321_));
  NAND_g _1344_ ( .A(T3y[0]), .B(_0321_), .Y(_0322_));
  AND_g _1345_ ( .A(SW[5]), .B(SW[6]), .Y(_0323_));
  AND_g _1346_ ( .A(SW[7]), .B(SW[8]), .Y(_0324_));
  NAND_g _1347_ ( .A(_0323_), .B(_0324_), .Y(_0325_));
  AND_g _1348_ ( .A(_0228_), .B(_0325_), .Y(_0326_));
  NOR_g _1349_ ( .A(T3plot), .B(_0326_), .Y(_0327_));
  AND_g _1350_ ( .A(_0295_), .B(_0318_), .Y(_0328_));
  AND_g _1351_ ( .A(_0213_), .B(_0328_), .Y(_0329_));
  NOR_g _1352_ ( .A(_0327_), .B(_0329_), .Y(_0330_));
  NAND_g _1353_ ( .A(_0322_), .B(_0330_), .Y(_0157_));
  NAND_g _1354_ ( .A(T3y[1]), .B(_0321_), .Y(_0331_));
  XNOR_g _1355_ ( .A(T3y[0]), .B(T3y[1]), .Y(_0332_));
  NAND_g _1356_ ( .A(_0328_), .B(_0332_), .Y(_0333_));
  NAND_g _1357_ ( .A(_0229_), .B(_0325_), .Y(_0334_));
  NAND_g _1358_ ( .A(_0301_), .B(_0334_), .Y(_0335_));
  NOT_g _1359_ ( .A(_0335_), .Y(_0336_));
  AND_g _1360_ ( .A(_0333_), .B(_0335_), .Y(_0337_));
  NAND_g _1361_ ( .A(_0331_), .B(_0337_), .Y(_0158_));
  NAND_g _1362_ ( .A(_0243_), .B(_0320_), .Y(_0338_));
  AND_g _1363_ ( .A(T3y[2]), .B(T3plot), .Y(_0339_));
  NAND_g _1364_ ( .A(_0338_), .B(_0339_), .Y(_0340_));
  AND_g _1365_ ( .A(SW[5]), .B(_0301_), .Y(_0341_));
  AND_g _1366_ ( .A(_0325_), .B(_0341_), .Y(_0342_));
  NAND_g _1367_ ( .A(_0325_), .B(_0341_), .Y(_0343_));
  NAND_g _1368_ ( .A(_0245_), .B(_0328_), .Y(_0344_));
  AND_g _1369_ ( .A(_0343_), .B(_0344_), .Y(_0345_));
  NAND_g _1370_ ( .A(_0340_), .B(_0345_), .Y(_0159_));
  NAND_g _1371_ ( .A(_0245_), .B(_0320_), .Y(_0346_));
  AND_g _1372_ ( .A(T3y[3]), .B(T3plot), .Y(_0347_));
  NAND_g _1373_ ( .A(_0346_), .B(_0347_), .Y(_0348_));
  NAND_g _1374_ ( .A(SW[6]), .B(_0301_), .Y(_0349_));
  NAND_g _1375_ ( .A(_0246_), .B(_0328_), .Y(_0350_));
  AND_g _1376_ ( .A(_0349_), .B(_0350_), .Y(_0351_));
  NAND_g _1377_ ( .A(_0348_), .B(_0351_), .Y(_0160_));
  NAND_g _1378_ ( .A(_0246_), .B(_0320_), .Y(_0352_));
  AND_g _1379_ ( .A(T3y[4]), .B(T3plot), .Y(_0353_));
  NAND_g _1380_ ( .A(_0352_), .B(_0353_), .Y(_0354_));
  AND_g _1381_ ( .A(SW[7]), .B(_0301_), .Y(_0355_));
  NAND_g _1382_ ( .A(SW[7]), .B(_0301_), .Y(_0356_));
  NAND_g _1383_ ( .A(_0247_), .B(_0328_), .Y(_0357_));
  AND_g _1384_ ( .A(_0356_), .B(_0357_), .Y(_0358_));
  NAND_g _1385_ ( .A(_0354_), .B(_0358_), .Y(_0161_));
  NAND_g _1386_ ( .A(SW[8]), .B(_0301_), .Y(_0359_));
  NAND_g _1387_ ( .A(T3y[5]), .B(_0321_), .Y(_0360_));
  XNOR_g _1388_ ( .A(_0218_), .B(_0247_), .Y(_0361_));
  NAND_g _1389_ ( .A(_0328_), .B(_0361_), .Y(_0362_));
  AND_g _1390_ ( .A(_0359_), .B(_0362_), .Y(_0363_));
  NAND_g _1391_ ( .A(_0360_), .B(_0363_), .Y(_0162_));
  NAND_g _1392_ ( .A(_0250_), .B(_0328_), .Y(_0364_));
  NAND_g _1393_ ( .A(_0249_), .B(_0320_), .Y(_0365_));
  AND_g _1394_ ( .A(T3y[6]), .B(T3plot), .Y(_0366_));
  NAND_g _1395_ ( .A(_0365_), .B(_0366_), .Y(_0367_));
  NAND_g _1396_ ( .A(_0364_), .B(_0367_), .Y(_0163_));
  NAND_g _1397_ ( .A(SW[0]), .B(_0301_), .Y(_0368_));
  NAND_g _1398_ ( .A(T3colourcircle[0]), .B(T3plot), .Y(_0369_));
  NAND_g _1399_ ( .A(_0368_), .B(_0369_), .Y(_0164_));
  NAND_g _1400_ ( .A(SW[1]), .B(_0301_), .Y(_0370_));
  NAND_g _1401_ ( .A(T3colourcircle[1]), .B(T3plot), .Y(_0371_));
  NAND_g _1402_ ( .A(_0370_), .B(_0371_), .Y(_0165_));
  NAND_g _1403_ ( .A(SW[2]), .B(_0301_), .Y(_0372_));
  NAND_g _1404_ ( .A(T3colourcircle[2]), .B(T3plot), .Y(_0373_));
  NAND_g _1405_ ( .A(_0372_), .B(_0373_), .Y(_0166_));
  NAND_g _1406_ ( .A(_0296_), .B(_0303_), .Y(_0374_));
  NOT_g _1407_ ( .A(_0374_), .Y(_0375_));
  NAND_g _1408_ ( .A(_0253_), .B(_0375_), .Y(_0376_));
  AND_g _1409_ ( .A(T3y[0]), .B(1'h1), .Y(_0377_));
  NAND_g _1410_ ( .A(T3y[0]), .B(1'h1), .Y(_0378_));
  XOR_g _1411_ ( .A(T3y[0]), .B(1'h1), .Y(_0379_));
  NAND_g _1412_ ( .A(_0376_), .B(_0379_), .Y(_0380_));
  AND_g _1413_ ( .A(_0259_), .B(_0264_), .Y(_0381_));
  NAND_g _1414_ ( .A(_0259_), .B(_0264_), .Y(_0382_));
  NOR_g _1415_ ( .A(_0260_), .B(_0305_), .Y(_0383_));
  NAND_g _1416_ ( .A(T3x[0]), .B(_0230_), .Y(_0384_));
  XNOR_g _1417_ ( .A(T3x[0]), .B(1'h1), .Y(_0385_));
  NOR_g _1418_ ( .A(_0383_), .B(_0385_), .Y(_0386_));
  NAND_g _1419_ ( .A(T3xp[0]), .B(_0239_), .Y(_0387_));
  NAND_g _1420_ ( .A(1'h1), .B(_0301_), .Y(_0388_));
  NAND_g _1421_ ( .A(_0387_), .B(_0388_), .Y(_0389_));
  NOR_g _1422_ ( .A(_0386_), .B(_0389_), .Y(_0390_));
  NAND_g _1423_ ( .A(_0380_), .B(_0390_), .Y(_0167_));
  NAND_g _1424_ ( .A(T3y[1]), .B(1'h1), .Y(_0391_));
  XOR_g _1425_ ( .A(T3y[1]), .B(1'h1), .Y(_0392_));
  XNOR_g _1426_ ( .A(T3y[1]), .B(1'h1), .Y(_0393_));
  NAND_g _1427_ ( .A(T3y[0]), .B(_0230_), .Y(_0394_));
  NAND_g _1428_ ( .A(_0393_), .B(_0394_), .Y(_0395_));
  XNOR_g _1429_ ( .A(_0392_), .B(_0394_), .Y(_0396_));
  NAND_g _1430_ ( .A(_0374_), .B(_0396_), .Y(_0397_));
  NAND_g _1431_ ( .A(T3xp[1]), .B(_0239_), .Y(_0398_));
  NAND_g _1432_ ( .A(1'h1), .B(_0301_), .Y(_0399_));
  AND_g _1433_ ( .A(_0398_), .B(_0399_), .Y(_0400_));
  NAND_g _1434_ ( .A(T3x[1]), .B(1'h1), .Y(_0401_));
  XOR_g _1435_ ( .A(T3x[1]), .B(1'h1), .Y(_0402_));
  XNOR_g _1436_ ( .A(T3x[1]), .B(1'h1), .Y(_0403_));
  NAND_g _1437_ ( .A(_0384_), .B(_0403_), .Y(_0404_));
  XNOR_g _1438_ ( .A(_0384_), .B(_0402_), .Y(_0405_));
  NAND_g _1439_ ( .A(_0305_), .B(_0405_), .Y(_0406_));
  AND_g _1440_ ( .A(T3x[0]), .B(1'h1), .Y(_0407_));
  NAND_g _1441_ ( .A(T3x[0]), .B(1'h1), .Y(_0408_));
  NAND_g _1442_ ( .A(_0403_), .B(_0408_), .Y(_0409_));
  NAND_g _1443_ ( .A(_0402_), .B(_0407_), .Y(_0410_));
  AND_g _1444_ ( .A(_0260_), .B(_0409_), .Y(_0411_));
  NAND_g _1445_ ( .A(_0410_), .B(_0411_), .Y(_0412_));
  NAND_g _1446_ ( .A(_0378_), .B(_0393_), .Y(_0413_));
  NAND_g _1447_ ( .A(_0377_), .B(_0392_), .Y(_0414_));
  AND_g _1448_ ( .A(_0252_), .B(_0413_), .Y(_0415_));
  NAND_g _1449_ ( .A(_0414_), .B(_0415_), .Y(_0416_));
  AND_g _1450_ ( .A(_0406_), .B(_0412_), .Y(_0417_));
  AND_g _1451_ ( .A(_0400_), .B(_0416_), .Y(_0418_));
  AND_g _1452_ ( .A(_0397_), .B(_0418_), .Y(_0419_));
  NAND_g _1453_ ( .A(_0417_), .B(_0419_), .Y(_0168_));
  NAND_g _1454_ ( .A(T3y[2]), .B(1'h1), .Y(_0420_));
  XOR_g _1455_ ( .A(T3y[2]), .B(1'h1), .Y(_0421_));
  XNOR_g _1456_ ( .A(T3y[2]), .B(1'h1), .Y(_0422_));
  NAND_g _1457_ ( .A(_0391_), .B(_0414_), .Y(_0423_));
  NAND_g _1458_ ( .A(_0421_), .B(_0423_), .Y(_0424_));
  XNOR_g _1459_ ( .A(_0422_), .B(_0423_), .Y(_0425_));
  NAND_g _1460_ ( .A(_0252_), .B(_0425_), .Y(_0426_));
  NAND_g _1461_ ( .A(T3xp[2]), .B(_0239_), .Y(_0427_));
  NAND_g _1462_ ( .A(1'h1), .B(_0301_), .Y(_0428_));
  AND_g _1463_ ( .A(_0427_), .B(_0428_), .Y(_0429_));
  AND_g _1464_ ( .A(_0426_), .B(_0429_), .Y(_0430_));
  NAND_g _1465_ ( .A(_0214_), .B(1'h1), .Y(_0431_));
  NAND_g _1466_ ( .A(_0395_), .B(_0431_), .Y(_0432_));
  NAND_g _1467_ ( .A(_0422_), .B(_0432_), .Y(_0433_));
  XNOR_g _1468_ ( .A(_0421_), .B(_0432_), .Y(_0434_));
  NAND_g _1469_ ( .A(_0374_), .B(_0434_), .Y(_0435_));
  NAND_g _1470_ ( .A(T3x[2]), .B(1'h1), .Y(_0436_));
  XOR_g _1471_ ( .A(T3x[2]), .B(1'h1), .Y(_0437_));
  XNOR_g _1472_ ( .A(T3x[2]), .B(1'h1), .Y(_0438_));
  AND_g _1473_ ( .A(_0401_), .B(_0410_), .Y(_0439_));
  NAND_g _1474_ ( .A(_0401_), .B(_0410_), .Y(_0440_));
  NAND_g _1475_ ( .A(_0437_), .B(_0440_), .Y(_0441_));
  NAND_g _1476_ ( .A(_0438_), .B(_0439_), .Y(_0442_));
  AND_g _1477_ ( .A(_0260_), .B(_0442_), .Y(_0443_));
  NAND_g _1478_ ( .A(_0441_), .B(_0443_), .Y(_0444_));
  NAND_g _1479_ ( .A(_0222_), .B(1'h1), .Y(_0445_));
  AND_g _1480_ ( .A(_0404_), .B(_0445_), .Y(_0446_));
  NAND_g _1481_ ( .A(_0404_), .B(_0445_), .Y(_0447_));
  NAND_g _1482_ ( .A(_0437_), .B(_0446_), .Y(_0448_));
  NAND_g _1483_ ( .A(_0438_), .B(_0447_), .Y(_0449_));
  AND_g _1484_ ( .A(_0305_), .B(_0449_), .Y(_0450_));
  NAND_g _1485_ ( .A(_0448_), .B(_0450_), .Y(_0451_));
  AND_g _1486_ ( .A(_0435_), .B(_0451_), .Y(_0452_));
  AND_g _1487_ ( .A(_0430_), .B(_0444_), .Y(_0453_));
  NAND_g _1488_ ( .A(_0452_), .B(_0453_), .Y(_0169_));
  NAND_g _1489_ ( .A(T3xp[3]), .B(_0239_), .Y(_0454_));
  NAND_g _1490_ ( .A(1'h1), .B(_0301_), .Y(_0455_));
  AND_g _1491_ ( .A(_0454_), .B(_0455_), .Y(_0456_));
  NAND_g _1492_ ( .A(_0216_), .B(_0231_), .Y(_0457_));
  NAND_g _1493_ ( .A(T3y[3]), .B(1'h1), .Y(_0458_));
  XOR_g _1494_ ( .A(T3y[3]), .B(1'h1), .Y(_0459_));
  AND_g _1495_ ( .A(_0420_), .B(_0424_), .Y(_0460_));
  XNOR_g _1496_ ( .A(_0459_), .B(_0460_), .Y(_0461_));
  NAND_g _1497_ ( .A(_0252_), .B(_0461_), .Y(_0462_));
  NAND_g _1498_ ( .A(_0224_), .B(_0231_), .Y(_0463_));
  NAND_g _1499_ ( .A(T3x[3]), .B(1'h1), .Y(_0464_));
  XNOR_g _1500_ ( .A(T3x[3]), .B(1'h1), .Y(_0465_));
  NAND_g _1501_ ( .A(_0223_), .B(1'h1), .Y(_0466_));
  NAND_g _1502_ ( .A(_0449_), .B(_0466_), .Y(_0467_));
  XOR_g _1503_ ( .A(_0465_), .B(_0467_), .Y(_0468_));
  NAND_g _1504_ ( .A(_0305_), .B(_0468_), .Y(_0469_));
  NAND_g _1505_ ( .A(_0215_), .B(1'h1), .Y(_0470_));
  AND_g _1506_ ( .A(_0433_), .B(_0470_), .Y(_0471_));
  XOR_g _1507_ ( .A(_0459_), .B(_0471_), .Y(_0472_));
  NAND_g _1508_ ( .A(_0374_), .B(_0472_), .Y(_0473_));
  AND_g _1509_ ( .A(_0436_), .B(_0441_), .Y(_0474_));
  XOR_g _1510_ ( .A(_0465_), .B(_0474_), .Y(_0475_));
  NAND_g _1511_ ( .A(_0260_), .B(_0475_), .Y(_0476_));
  AND_g _1512_ ( .A(_0456_), .B(_0473_), .Y(_0477_));
  AND_g _1513_ ( .A(_0462_), .B(_0469_), .Y(_0478_));
  AND_g _1514_ ( .A(_0476_), .B(_0478_), .Y(_0479_));
  NAND_g _1515_ ( .A(_0477_), .B(_0479_), .Y(_0170_));
  NAND_g _1516_ ( .A(T3y[4]), .B(1'h0), .Y(_0480_));
  XOR_g _1517_ ( .A(T3y[4]), .B(1'h0), .Y(_0481_));
  XNOR_g _1518_ ( .A(T3y[4]), .B(1'h0), .Y(_0482_));
  NAND_g _1519_ ( .A(_0458_), .B(_0460_), .Y(_0483_));
  AND_g _1520_ ( .A(_0457_), .B(_0483_), .Y(_0484_));
  NAND_g _1521_ ( .A(_0481_), .B(_0484_), .Y(_0485_));
  XNOR_g _1522_ ( .A(_0482_), .B(_0484_), .Y(_0486_));
  NAND_g _1523_ ( .A(_0252_), .B(_0486_), .Y(_0487_));
  NAND_g _1524_ ( .A(T3x[4]), .B(1'h0), .Y(_0488_));
  XOR_g _1525_ ( .A(T3x[4]), .B(1'h0), .Y(_0489_));
  XNOR_g _1526_ ( .A(T3x[4]), .B(1'h0), .Y(_0490_));
  NAND_g _1527_ ( .A(_0464_), .B(_0474_), .Y(_0491_));
  AND_g _1528_ ( .A(_0463_), .B(_0491_), .Y(_0492_));
  NOR_g _1529_ ( .A(_0489_), .B(_0492_), .Y(_0493_));
  NAND_g _1530_ ( .A(_0489_), .B(_0492_), .Y(_0494_));
  NAND_g _1531_ ( .A(_0260_), .B(_0494_), .Y(_0495_));
  NOR_g _1532_ ( .A(_0493_), .B(_0495_), .Y(_0496_));
  NAND_g _1533_ ( .A(T3xp[4]), .B(_0239_), .Y(_0497_));
  NAND_g _1534_ ( .A(1'h0), .B(_0301_), .Y(_0498_));
  NAND_g _1535_ ( .A(_0497_), .B(_0498_), .Y(_0499_));
  NOR_g _1536_ ( .A(_0496_), .B(_0499_), .Y(_0500_));
  AND_g _1537_ ( .A(_0487_), .B(_0500_), .Y(_0501_));
  NAND_g _1538_ ( .A(T3x[3]), .B(_0231_), .Y(_0502_));
  NAND_g _1539_ ( .A(_0224_), .B(1'h1), .Y(_0503_));
  NAND_g _1540_ ( .A(_0467_), .B(_0502_), .Y(_0504_));
  NAND_g _1541_ ( .A(_0503_), .B(_0504_), .Y(_0505_));
  AND_g _1542_ ( .A(_0503_), .B(_0504_), .Y(_0506_));
  NAND_g _1543_ ( .A(_0489_), .B(_0506_), .Y(_0507_));
  NAND_g _1544_ ( .A(_0490_), .B(_0505_), .Y(_0508_));
  AND_g _1545_ ( .A(_0305_), .B(_0508_), .Y(_0509_));
  NAND_g _1546_ ( .A(_0507_), .B(_0509_), .Y(_0510_));
  NAND_g _1547_ ( .A(T3y[3]), .B(_0231_), .Y(_0511_));
  NAND_g _1548_ ( .A(_0216_), .B(1'h1), .Y(_0512_));
  NAND_g _1549_ ( .A(_0471_), .B(_0512_), .Y(_0513_));
  AND_g _1550_ ( .A(_0511_), .B(_0513_), .Y(_0514_));
  NAND_g _1551_ ( .A(_0482_), .B(_0514_), .Y(_0515_));
  XNOR_g _1552_ ( .A(_0481_), .B(_0514_), .Y(_0516_));
  NAND_g _1553_ ( .A(_0374_), .B(_0516_), .Y(_0517_));
  AND_g _1554_ ( .A(_0510_), .B(_0517_), .Y(_0518_));
  NAND_g _1555_ ( .A(_0501_), .B(_0518_), .Y(_0171_));
  NAND_g _1556_ ( .A(_0226_), .B(_0232_), .Y(_0519_));
  NAND_g _1557_ ( .A(T3x[5]), .B(1'h0), .Y(_0520_));
  XOR_g _1558_ ( .A(T3x[5]), .B(1'h0), .Y(_0521_));
  NAND_g _1559_ ( .A(_0225_), .B(1'h0), .Y(_0522_));
  NAND_g _1560_ ( .A(_0508_), .B(_0522_), .Y(_0523_));
  AND_g _1561_ ( .A(_0488_), .B(_0494_), .Y(_0524_));
  NAND_g _1562_ ( .A(_0218_), .B(_0232_), .Y(_0525_));
  NAND_g _1563_ ( .A(T3y[5]), .B(1'h0), .Y(_0526_));
  XOR_g _1564_ ( .A(T3y[5]), .B(1'h0), .Y(_0527_));
  AND_g _1565_ ( .A(_0480_), .B(_0485_), .Y(_0528_));
  XNOR_g _1566_ ( .A(_0527_), .B(_0528_), .Y(_0529_));
  NAND_g _1567_ ( .A(_0252_), .B(_0529_), .Y(_0530_));
  NAND_g _1568_ ( .A(T3xp[5]), .B(_0239_), .Y(_0531_));
  NAND_g _1569_ ( .A(1'h0), .B(_0301_), .Y(_0532_));
  AND_g _1570_ ( .A(_0531_), .B(_0532_), .Y(_0533_));
  NAND_g _1571_ ( .A(_0217_), .B(1'h0), .Y(_0534_));
  AND_g _1572_ ( .A(_0515_), .B(_0534_), .Y(_0535_));
  XOR_g _1573_ ( .A(_0527_), .B(_0535_), .Y(_0536_));
  NAND_g _1574_ ( .A(_0374_), .B(_0536_), .Y(_0537_));
  AND_g _1575_ ( .A(_0530_), .B(_0537_), .Y(_0538_));
  XNOR_g _1576_ ( .A(_0521_), .B(_0524_), .Y(_0539_));
  NAND_g _1577_ ( .A(_0260_), .B(_0539_), .Y(_0540_));
  XNOR_g _1578_ ( .A(_0521_), .B(_0523_), .Y(_0541_));
  NAND_g _1579_ ( .A(_0305_), .B(_0541_), .Y(_0542_));
  AND_g _1580_ ( .A(_0533_), .B(_0542_), .Y(_0543_));
  AND_g _1581_ ( .A(_0540_), .B(_0543_), .Y(_0544_));
  NAND_g _1582_ ( .A(_0538_), .B(_0544_), .Y(_0172_));
  NAND_g _1583_ ( .A(T3x[6]), .B(1'h1), .Y(_0545_));
  XOR_g _1584_ ( .A(T3x[6]), .B(1'h1), .Y(_0546_));
  XNOR_g _1585_ ( .A(T3x[6]), .B(1'h1), .Y(_0547_));
  NAND_g _1586_ ( .A(_0520_), .B(_0524_), .Y(_0548_));
  AND_g _1587_ ( .A(_0519_), .B(_0548_), .Y(_0549_));
  NAND_g _1588_ ( .A(_0546_), .B(_0549_), .Y(_0550_));
  XNOR_g _1589_ ( .A(_0547_), .B(_0549_), .Y(_0551_));
  NAND_g _1590_ ( .A(_0260_), .B(_0551_), .Y(_0552_));
  NAND_g _1591_ ( .A(1'h1), .B(_0301_), .Y(_0553_));
  NAND_g _1592_ ( .A(T3xp[6]), .B(_0239_), .Y(_0554_));
  AND_g _1593_ ( .A(_0553_), .B(_0554_), .Y(_0555_));
  NAND_g _1594_ ( .A(T3y[6]), .B(1'h1), .Y(_0556_));
  XOR_g _1595_ ( .A(T3y[6]), .B(1'h1), .Y(_0557_));
  XNOR_g _1596_ ( .A(T3y[6]), .B(1'h1), .Y(_0558_));
  NAND_g _1597_ ( .A(_0526_), .B(_0528_), .Y(_0559_));
  AND_g _1598_ ( .A(_0525_), .B(_0559_), .Y(_0560_));
  NAND_g _1599_ ( .A(_0557_), .B(_0560_), .Y(_0561_));
  XNOR_g _1600_ ( .A(_0558_), .B(_0560_), .Y(_0562_));
  NAND_g _1601_ ( .A(_0252_), .B(_0562_), .Y(_0563_));
  AND_g _1602_ ( .A(_0555_), .B(_0563_), .Y(_0564_));
  AND_g _1603_ ( .A(_0552_), .B(_0564_), .Y(_0565_));
  NAND_g _1604_ ( .A(_0218_), .B(1'h0), .Y(_0566_));
  NAND_g _1605_ ( .A(T3y[5]), .B(_0232_), .Y(_0567_));
  NAND_g _1606_ ( .A(_0535_), .B(_0566_), .Y(_0568_));
  AND_g _1607_ ( .A(_0567_), .B(_0568_), .Y(_0569_));
  NAND_g _1608_ ( .A(_0558_), .B(_0569_), .Y(_0570_));
  XNOR_g _1609_ ( .A(_0557_), .B(_0569_), .Y(_0571_));
  NAND_g _1610_ ( .A(_0374_), .B(_0571_), .Y(_0572_));
  NAND_g _1611_ ( .A(_0226_), .B(1'h0), .Y(_0573_));
  NAND_g _1612_ ( .A(T3x[5]), .B(_0232_), .Y(_0574_));
  NAND_g _1613_ ( .A(_0523_), .B(_0574_), .Y(_0575_));
  AND_g _1614_ ( .A(_0573_), .B(_0575_), .Y(_0576_));
  NAND_g _1615_ ( .A(_0573_), .B(_0575_), .Y(_0577_));
  NAND_g _1616_ ( .A(_0547_), .B(_0577_), .Y(_0578_));
  NAND_g _1617_ ( .A(_0546_), .B(_0576_), .Y(_0579_));
  AND_g _1618_ ( .A(_0305_), .B(_0579_), .Y(_0580_));
  NAND_g _1619_ ( .A(_0578_), .B(_0580_), .Y(_0581_));
  AND_g _1620_ ( .A(_0572_), .B(_0581_), .Y(_0582_));
  NAND_g _1621_ ( .A(_0565_), .B(_0582_), .Y(_0173_));
  AND_g _1622_ ( .A(_0556_), .B(_0561_), .Y(_0583_));
  XNOR_g _1623_ ( .A(1'h0), .B(_0583_), .Y(_0584_));
  NAND_g _1624_ ( .A(_0252_), .B(_0584_), .Y(_0585_));
  NAND_g _1625_ ( .A(T3xp[7]), .B(_0239_), .Y(_0586_));
  NAND_g _1626_ ( .A(1'h0), .B(_0301_), .Y(_0587_));
  AND_g _1627_ ( .A(_0586_), .B(_0587_), .Y(_0588_));
  XOR_g _1628_ ( .A(T3x[7]), .B(1'h0), .Y(_0589_));
  AND_g _1629_ ( .A(_0545_), .B(_0550_), .Y(_0590_));
  XNOR_g _1630_ ( .A(_0589_), .B(_0590_), .Y(_0591_));
  NAND_g _1631_ ( .A(_0260_), .B(_0591_), .Y(_0592_));
  NAND_g _1632_ ( .A(_0227_), .B(1'h1), .Y(_0593_));
  NAND_g _1633_ ( .A(_0578_), .B(_0593_), .Y(_0594_));
  XNOR_g _1634_ ( .A(_0589_), .B(_0594_), .Y(_0595_));
  NAND_g _1635_ ( .A(_0305_), .B(_0595_), .Y(_0596_));
  NAND_g _1636_ ( .A(_0219_), .B(1'h1), .Y(_0597_));
  NAND_g _1637_ ( .A(_0570_), .B(_0597_), .Y(_0598_));
  XNOR_g _1638_ ( .A(1'h0), .B(_0598_), .Y(_0599_));
  NAND_g _1639_ ( .A(_0374_), .B(_0599_), .Y(_0600_));
  AND_g _1640_ ( .A(_0588_), .B(_0596_), .Y(_0601_));
  AND_g _1641_ ( .A(_0585_), .B(_0592_), .Y(_0602_));
  AND_g _1642_ ( .A(_0600_), .B(_0602_), .Y(_0603_));
  NAND_g _1643_ ( .A(_0601_), .B(_0603_), .Y(_0174_));
  NOR_g _1644_ ( .A(T3d[0]), .B(_0301_), .Y(_0604_));
  NOT_g _1645_ ( .A(_0604_), .Y(_0175_));
  NAND_g _1646_ ( .A(_0301_), .B(_0326_), .Y(_0605_));
  AND_g _1647_ ( .A(T3d[1]), .B(_0238_), .Y(_0606_));
  AND_g _1648_ ( .A(_0220_), .B(_0295_), .Y(_0607_));
  NOR_g _1649_ ( .A(_0606_), .B(_0607_), .Y(_0608_));
  NAND_g _1650_ ( .A(_0605_), .B(_0608_), .Y(_0176_));
  NAND_g _1651_ ( .A(T3y[0]), .B(T3x[0]), .Y(_0609_));
  XNOR_g _1652_ ( .A(T3y[0]), .B(T3x[0]), .Y(_0610_));
  AND_g _1653_ ( .A(T3d[2]), .B(_0610_), .Y(_0611_));
  XOR_g _1654_ ( .A(T3d[2]), .B(_0610_), .Y(_0612_));
  AND_g _1655_ ( .A(T3d[2]), .B(_0221_), .Y(_0613_));
  XOR_g _1656_ ( .A(T3d[2]), .B(T3x[0]), .Y(_0614_));
  NAND_g _1657_ ( .A(_0319_), .B(_0614_), .Y(_0615_));
  NAND_g _1658_ ( .A(_0318_), .B(_0612_), .Y(_0616_));
  NAND_g _1659_ ( .A(_0615_), .B(_0616_), .Y(_0617_));
  AND_g _1660_ ( .A(_0615_), .B(_0616_), .Y(_0618_));
  NAND_g _1661_ ( .A(_0607_), .B(_0617_), .Y(_0619_));
  AND_g _1662_ ( .A(T3d[1]), .B(_0295_), .Y(_0620_));
  NAND_g _1663_ ( .A(_0618_), .B(_0620_), .Y(_0621_));
  NAND_g _1664_ ( .A(T3d[2]), .B(_0238_), .Y(_0622_));
  AND_g _1665_ ( .A(_0335_), .B(_0622_), .Y(_0623_));
  AND_g _1666_ ( .A(_0621_), .B(_0623_), .Y(_0624_));
  NAND_g _1667_ ( .A(_0619_), .B(_0624_), .Y(_0177_));
  AND_g _1668_ ( .A(T3d[1]), .B(_0612_), .Y(_0625_));
  NAND_g _1669_ ( .A(T3d[1]), .B(_0612_), .Y(_0626_));
  AND_g _1670_ ( .A(T3x[0]), .B(T3x[1]), .Y(_0627_));
  XOR_g _1671_ ( .A(T3x[0]), .B(T3x[1]), .Y(_0628_));
  NAND_g _1672_ ( .A(_0214_), .B(_0628_), .Y(_0629_));
  XNOR_g _1673_ ( .A(T3y[1]), .B(_0628_), .Y(_0630_));
  NAND_g _1674_ ( .A(_0609_), .B(_0630_), .Y(_0631_));
  XOR_g _1675_ ( .A(_0609_), .B(_0630_), .Y(_0632_));
  NAND_g _1676_ ( .A(T3d[3]), .B(_0632_), .Y(_0633_));
  XOR_g _1677_ ( .A(T3d[3]), .B(_0632_), .Y(_0634_));
  NAND_g _1678_ ( .A(_0611_), .B(_0634_), .Y(_0635_));
  XNOR_g _1679_ ( .A(_0611_), .B(_0634_), .Y(_0636_));
  NAND_g _1680_ ( .A(_0626_), .B(_0636_), .Y(_0637_));
  NAND_g _1681_ ( .A(_0625_), .B(_0634_), .Y(_0638_));
  NAND_g _1682_ ( .A(_0220_), .B(_0614_), .Y(_0639_));
  NAND_g _1683_ ( .A(T3d[3]), .B(_0628_), .Y(_0640_));
  XOR_g _1684_ ( .A(T3d[3]), .B(_0628_), .Y(_0641_));
  NAND_g _1685_ ( .A(_0613_), .B(_0641_), .Y(_0642_));
  XOR_g _1686_ ( .A(_0613_), .B(_0641_), .Y(_0643_));
  AND_g _1687_ ( .A(_0639_), .B(_0643_), .Y(_0644_));
  XOR_g _1688_ ( .A(_0639_), .B(_0643_), .Y(_0645_));
  NOR_g _1689_ ( .A(_0318_), .B(_0645_), .Y(_0646_));
  NOR_g _1690_ ( .A(_0296_), .B(_0646_), .Y(_0647_));
  AND_g _1691_ ( .A(_0318_), .B(_0638_), .Y(_0648_));
  NAND_g _1692_ ( .A(_0637_), .B(_0648_), .Y(_0649_));
  NAND_g _1693_ ( .A(_0647_), .B(_0649_), .Y(_0650_));
  AND_g _1694_ ( .A(T3d[3]), .B(_0238_), .Y(_0651_));
  AND_g _1695_ ( .A(_0335_), .B(_0343_), .Y(_0652_));
  AND_g _1696_ ( .A(SW[4]), .B(_0342_), .Y(_0653_));
  NOR_g _1697_ ( .A(_0652_), .B(_0653_), .Y(_0654_));
  NOR_g _1698_ ( .A(_0651_), .B(_0654_), .Y(_0655_));
  NAND_g _1699_ ( .A(_0650_), .B(_0655_), .Y(_0178_));
  NAND_g _1700_ ( .A(_0633_), .B(_0635_), .Y(_0656_));
  NAND_g _1701_ ( .A(_0629_), .B(_0631_), .Y(_0657_));
  AND_g _1702_ ( .A(T3x[2]), .B(_0627_), .Y(_0658_));
  XNOR_g _1703_ ( .A(_0223_), .B(_0627_), .Y(_0659_));
  NAND_g _1704_ ( .A(_0215_), .B(_0659_), .Y(_0660_));
  XNOR_g _1705_ ( .A(T3y[2]), .B(_0659_), .Y(_0661_));
  NAND_g _1706_ ( .A(_0657_), .B(_0661_), .Y(_0662_));
  XOR_g _1707_ ( .A(_0657_), .B(_0661_), .Y(_0663_));
  NAND_g _1708_ ( .A(T3d[4]), .B(_0663_), .Y(_0664_));
  XOR_g _1709_ ( .A(T3d[4]), .B(_0663_), .Y(_0665_));
  NAND_g _1710_ ( .A(_0656_), .B(_0665_), .Y(_0666_));
  XOR_g _1711_ ( .A(_0656_), .B(_0665_), .Y(_0667_));
  AND_g _1712_ ( .A(_0637_), .B(_0667_), .Y(_0668_));
  XOR_g _1713_ ( .A(_0637_), .B(_0667_), .Y(_0669_));
  NAND_g _1714_ ( .A(_0318_), .B(_0669_), .Y(_0670_));
  NAND_g _1715_ ( .A(_0640_), .B(_0642_), .Y(_0671_));
  NAND_g _1716_ ( .A(T3d[4]), .B(_0659_), .Y(_0672_));
  XOR_g _1717_ ( .A(T3d[4]), .B(_0659_), .Y(_0673_));
  NAND_g _1718_ ( .A(_0671_), .B(_0673_), .Y(_0674_));
  XOR_g _1719_ ( .A(_0671_), .B(_0673_), .Y(_0675_));
  AND_g _1720_ ( .A(_0644_), .B(_0675_), .Y(_0676_));
  NOT_g _1721_ ( .A(_0676_), .Y(_0677_));
  NOR_g _1722_ ( .A(_0644_), .B(_0675_), .Y(_0678_));
  NOR_g _1723_ ( .A(_0318_), .B(_0678_), .Y(_0679_));
  NAND_g _1724_ ( .A(_0677_), .B(_0679_), .Y(_0680_));
  NAND_g _1725_ ( .A(_0670_), .B(_0680_), .Y(_0681_));
  NAND_g _1726_ ( .A(_0295_), .B(_0681_), .Y(_0682_));
  NAND_g _1727_ ( .A(T3d[4]), .B(_0238_), .Y(_0683_));
  AND_g _1728_ ( .A(_0349_), .B(_0652_), .Y(_0684_));
  XNOR_g _1729_ ( .A(_0349_), .B(_0652_), .Y(_0685_));
  AND_g _1730_ ( .A(_0683_), .B(_0685_), .Y(_0686_));
  NAND_g _1731_ ( .A(_0682_), .B(_0686_), .Y(_0179_));
  NAND_g _1732_ ( .A(_0664_), .B(_0666_), .Y(_0687_));
  NAND_g _1733_ ( .A(_0660_), .B(_0662_), .Y(_0688_));
  AND_g _1734_ ( .A(T3x[3]), .B(_0658_), .Y(_0689_));
  XNOR_g _1735_ ( .A(_0224_), .B(_0658_), .Y(_0690_));
  XNOR_g _1736_ ( .A(T3x[3]), .B(_0658_), .Y(_0691_));
  NAND_g _1737_ ( .A(_0216_), .B(_0690_), .Y(_0692_));
  NAND_g _1738_ ( .A(T3y[3]), .B(_0691_), .Y(_0693_));
  XNOR_g _1739_ ( .A(_0216_), .B(_0690_), .Y(_0694_));
  XNOR_g _1740_ ( .A(_0688_), .B(_0694_), .Y(_0695_));
  NAND_g _1741_ ( .A(T3d[5]), .B(_0695_), .Y(_0696_));
  XOR_g _1742_ ( .A(T3d[5]), .B(_0695_), .Y(_0697_));
  NAND_g _1743_ ( .A(_0687_), .B(_0697_), .Y(_0698_));
  XOR_g _1744_ ( .A(_0687_), .B(_0697_), .Y(_0699_));
  AND_g _1745_ ( .A(_0668_), .B(_0699_), .Y(_0700_));
  XOR_g _1746_ ( .A(_0668_), .B(_0699_), .Y(_0701_));
  NAND_g _1747_ ( .A(_0318_), .B(_0701_), .Y(_0702_));
  NAND_g _1748_ ( .A(_0672_), .B(_0674_), .Y(_0703_));
  NAND_g _1749_ ( .A(T3d[5]), .B(_0690_), .Y(_0704_));
  XNOR_g _1750_ ( .A(T3d[5]), .B(_0691_), .Y(_0705_));
  NAND_g _1751_ ( .A(_0703_), .B(_0705_), .Y(_0706_));
  XOR_g _1752_ ( .A(_0703_), .B(_0705_), .Y(_0707_));
  AND_g _1753_ ( .A(_0676_), .B(_0707_), .Y(_0708_));
  XNOR_g _1754_ ( .A(_0677_), .B(_0707_), .Y(_0709_));
  NAND_g _1755_ ( .A(_0319_), .B(_0709_), .Y(_0710_));
  NAND_g _1756_ ( .A(_0702_), .B(_0710_), .Y(_0711_));
  NAND_g _1757_ ( .A(_0295_), .B(_0711_), .Y(_0712_));
  NAND_g _1758_ ( .A(T3d[5]), .B(_0238_), .Y(_0713_));
  AND_g _1759_ ( .A(_0356_), .B(_0684_), .Y(_0714_));
  XNOR_g _1760_ ( .A(_0356_), .B(_0684_), .Y(_0715_));
  AND_g _1761_ ( .A(_0713_), .B(_0715_), .Y(_0716_));
  NAND_g _1762_ ( .A(_0712_), .B(_0716_), .Y(_0180_));
  NAND_g _1763_ ( .A(_0696_), .B(_0698_), .Y(_0717_));
  AND_g _1764_ ( .A(T3x[4]), .B(_0689_), .Y(_0718_));
  XNOR_g _1765_ ( .A(_0225_), .B(_0689_), .Y(_0719_));
  NAND_g _1766_ ( .A(_0217_), .B(_0719_), .Y(_0720_));
  XNOR_g _1767_ ( .A(T3y[4]), .B(_0719_), .Y(_0721_));
  NAND_g _1768_ ( .A(_0688_), .B(_0693_), .Y(_0722_));
  NAND_g _1769_ ( .A(_0692_), .B(_0722_), .Y(_0723_));
  NAND_g _1770_ ( .A(_0721_), .B(_0723_), .Y(_0724_));
  XOR_g _1771_ ( .A(_0721_), .B(_0723_), .Y(_0725_));
  NAND_g _1772_ ( .A(T3d[6]), .B(_0725_), .Y(_0726_));
  XOR_g _1773_ ( .A(T3d[6]), .B(_0725_), .Y(_0727_));
  NAND_g _1774_ ( .A(_0717_), .B(_0727_), .Y(_0728_));
  XOR_g _1775_ ( .A(_0717_), .B(_0727_), .Y(_0729_));
  AND_g _1776_ ( .A(_0700_), .B(_0729_), .Y(_0730_));
  XOR_g _1777_ ( .A(_0700_), .B(_0729_), .Y(_0731_));
  NAND_g _1778_ ( .A(_0318_), .B(_0731_), .Y(_0732_));
  NAND_g _1779_ ( .A(_0704_), .B(_0706_), .Y(_0733_));
  NAND_g _1780_ ( .A(T3d[6]), .B(_0719_), .Y(_0734_));
  XOR_g _1781_ ( .A(T3d[6]), .B(_0719_), .Y(_0735_));
  NAND_g _1782_ ( .A(_0733_), .B(_0735_), .Y(_0736_));
  XOR_g _1783_ ( .A(_0733_), .B(_0735_), .Y(_0737_));
  AND_g _1784_ ( .A(_0708_), .B(_0737_), .Y(_0738_));
  NOT_g _1785_ ( .A(_0738_), .Y(_0739_));
  NOR_g _1786_ ( .A(_0708_), .B(_0737_), .Y(_0740_));
  NOR_g _1787_ ( .A(_0318_), .B(_0740_), .Y(_0741_));
  NAND_g _1788_ ( .A(_0739_), .B(_0741_), .Y(_0742_));
  NAND_g _1789_ ( .A(_0732_), .B(_0742_), .Y(_0743_));
  NAND_g _1790_ ( .A(_0295_), .B(_0743_), .Y(_0744_));
  NAND_g _1791_ ( .A(T3d[6]), .B(_0238_), .Y(_0745_));
  AND_g _1792_ ( .A(_0359_), .B(_0714_), .Y(_0746_));
  XNOR_g _1793_ ( .A(_0359_), .B(_0714_), .Y(_0747_));
  AND_g _1794_ ( .A(_0745_), .B(_0747_), .Y(_0748_));
  NAND_g _1795_ ( .A(_0744_), .B(_0748_), .Y(_0181_));
  NAND_g _1796_ ( .A(_0726_), .B(_0728_), .Y(_0749_));
  NAND_g _1797_ ( .A(_0720_), .B(_0724_), .Y(_0750_));
  AND_g _1798_ ( .A(T3x[5]), .B(_0718_), .Y(_0751_));
  XNOR_g _1799_ ( .A(_0226_), .B(_0718_), .Y(_0752_));
  XNOR_g _1800_ ( .A(T3x[5]), .B(_0718_), .Y(_0753_));
  NAND_g _1801_ ( .A(_0218_), .B(_0752_), .Y(_0754_));
  NAND_g _1802_ ( .A(T3y[5]), .B(_0753_), .Y(_0755_));
  XNOR_g _1803_ ( .A(_0218_), .B(_0752_), .Y(_0756_));
  XNOR_g _1804_ ( .A(_0750_), .B(_0756_), .Y(_0757_));
  NAND_g _1805_ ( .A(T3d[7]), .B(_0757_), .Y(_0758_));
  XOR_g _1806_ ( .A(T3d[7]), .B(_0757_), .Y(_0759_));
  NAND_g _1807_ ( .A(_0749_), .B(_0759_), .Y(_0760_));
  XOR_g _1808_ ( .A(_0749_), .B(_0759_), .Y(_0761_));
  AND_g _1809_ ( .A(_0730_), .B(_0761_), .Y(_0762_));
  XOR_g _1810_ ( .A(_0730_), .B(_0761_), .Y(_0763_));
  NAND_g _1811_ ( .A(_0318_), .B(_0763_), .Y(_0764_));
  NAND_g _1812_ ( .A(_0734_), .B(_0736_), .Y(_0765_));
  NAND_g _1813_ ( .A(T3d[7]), .B(_0752_), .Y(_0766_));
  XNOR_g _1814_ ( .A(T3d[7]), .B(_0753_), .Y(_0767_));
  NAND_g _1815_ ( .A(_0765_), .B(_0767_), .Y(_0768_));
  XOR_g _1816_ ( .A(_0765_), .B(_0767_), .Y(_0769_));
  NOR_g _1817_ ( .A(_0738_), .B(_0769_), .Y(_0770_));
  NAND_g _1818_ ( .A(_0738_), .B(_0769_), .Y(_0771_));
  NOR_g _1819_ ( .A(_0318_), .B(_0770_), .Y(_0772_));
  NAND_g _1820_ ( .A(_0771_), .B(_0772_), .Y(_0773_));
  NAND_g _1821_ ( .A(_0764_), .B(_0773_), .Y(_0774_));
  NAND_g _1822_ ( .A(_0295_), .B(_0774_), .Y(_0775_));
  NAND_g _1823_ ( .A(T3d[7]), .B(_0238_), .Y(_0776_));
  AND_g _1824_ ( .A(_0746_), .B(_0776_), .Y(_0777_));
  NAND_g _1825_ ( .A(_0775_), .B(_0777_), .Y(_0182_));
  NAND_g _1826_ ( .A(_0758_), .B(_0760_), .Y(_0778_));
  NAND_g _1827_ ( .A(_0750_), .B(_0755_), .Y(_0779_));
  AND_g _1828_ ( .A(_0754_), .B(_0779_), .Y(_0780_));
  AND_g _1829_ ( .A(T3x[6]), .B(_0751_), .Y(_0781_));
  XNOR_g _1830_ ( .A(_0227_), .B(_0751_), .Y(_0782_));
  XNOR_g _1831_ ( .A(T3d[8]), .B(_0782_), .Y(_0783_));
  XNOR_g _1832_ ( .A(_0219_), .B(_0783_), .Y(_0784_));
  XNOR_g _1833_ ( .A(_0780_), .B(_0784_), .Y(_0785_));
  XNOR_g _1834_ ( .A(_0778_), .B(_0785_), .Y(_0786_));
  XNOR_g _1835_ ( .A(_0762_), .B(_0786_), .Y(_0787_));
  NAND_g _1836_ ( .A(_0318_), .B(_0787_), .Y(_0788_));
  NAND_g _1837_ ( .A(_0766_), .B(_0768_), .Y(_0789_));
  XNOR_g _1838_ ( .A(_0783_), .B(_0789_), .Y(_0790_));
  XNOR_g _1839_ ( .A(_0771_), .B(_0790_), .Y(_0791_));
  NAND_g _1840_ ( .A(_0319_), .B(_0791_), .Y(_0792_));
  NAND_g _1841_ ( .A(_0788_), .B(_0792_), .Y(_0793_));
  NAND_g _1842_ ( .A(_0295_), .B(_0793_), .Y(_0794_));
  NAND_g _1843_ ( .A(T3d[8]), .B(_0238_), .Y(_0795_));
  AND_g _1844_ ( .A(_0746_), .B(_0795_), .Y(_0796_));
  NAND_g _1845_ ( .A(_0794_), .B(_0796_), .Y(_0183_));
  NAND_g _1846_ ( .A(T3x[0]), .B(_0238_), .Y(_0797_));
  NAND_g _1847_ ( .A(_0221_), .B(_0295_), .Y(_0798_));
  NAND_g _1848_ ( .A(_0797_), .B(_0798_), .Y(_0184_));
  NAND_g _1849_ ( .A(T3x[1]), .B(_0238_), .Y(_0799_));
  NAND_g _1850_ ( .A(_0295_), .B(_0628_), .Y(_0800_));
  NAND_g _1851_ ( .A(_0799_), .B(_0800_), .Y(_0185_));
  NAND_g _1852_ ( .A(T3x[2]), .B(_0238_), .Y(_0801_));
  NAND_g _1853_ ( .A(_0295_), .B(_0659_), .Y(_0802_));
  NAND_g _1854_ ( .A(_0801_), .B(_0802_), .Y(_0186_));
  NAND_g _1855_ ( .A(T3x[3]), .B(_0238_), .Y(_0803_));
  NAND_g _1856_ ( .A(_0295_), .B(_0690_), .Y(_0804_));
  NAND_g _1857_ ( .A(_0803_), .B(_0804_), .Y(_0187_));
  NAND_g _1858_ ( .A(T3x[4]), .B(_0238_), .Y(_0805_));
  NAND_g _1859_ ( .A(_0295_), .B(_0719_), .Y(_0806_));
  NAND_g _1860_ ( .A(_0805_), .B(_0806_), .Y(_0188_));
  NAND_g _1861_ ( .A(T3x[5]), .B(_0238_), .Y(_0807_));
  NAND_g _1862_ ( .A(_0295_), .B(_0752_), .Y(_0808_));
  NAND_g _1863_ ( .A(_0807_), .B(_0808_), .Y(_0189_));
  NAND_g _1864_ ( .A(T3x[6]), .B(_0238_), .Y(_0809_));
  NAND_g _1865_ ( .A(_0295_), .B(_0782_), .Y(_0810_));
  NAND_g _1866_ ( .A(_0809_), .B(_0810_), .Y(_0190_));
  NAND_g _1867_ ( .A(_0297_), .B(_0781_), .Y(_0811_));
  NAND_g _1868_ ( .A(_0237_), .B(_0781_), .Y(_0812_));
  AND_g _1869_ ( .A(T3x[7]), .B(T3plot), .Y(_0813_));
  NAND_g _1870_ ( .A(_0812_), .B(_0813_), .Y(_0814_));
  NAND_g _1871_ ( .A(_0811_), .B(_0814_), .Y(_0191_));
  AND_g _1872_ ( .A(T3y[0]), .B(1'h1), .Y(_0815_));
  NAND_g _1873_ ( .A(T3y[0]), .B(_0233_), .Y(_0816_));
  XNOR_g _1874_ ( .A(T3y[0]), .B(1'h1), .Y(_0817_));
  NOR_g _1875_ ( .A(_0383_), .B(_0817_), .Y(_0818_));
  AND_g _1876_ ( .A(T3yp[0]), .B(_0239_), .Y(_0819_));
  NOR_g _1877_ ( .A(_0818_), .B(_0819_), .Y(_0820_));
  AND_g _1878_ ( .A(T3x[0]), .B(1'h1), .Y(_0821_));
  XOR_g _1879_ ( .A(T3x[0]), .B(1'h1), .Y(_0822_));
  AND_g _1880_ ( .A(_0376_), .B(_0822_), .Y(_0823_));
  NOR_g _1881_ ( .A(1'h1), .B(_0327_), .Y(_0824_));
  AND_g _1882_ ( .A(1'h1), .B(_0605_), .Y(_0825_));
  NOR_g _1883_ ( .A(_0824_), .B(_0825_), .Y(_0826_));
  NOR_g _1884_ ( .A(_0823_), .B(_0826_), .Y(_0827_));
  NAND_g _1885_ ( .A(_0820_), .B(_0827_), .Y(_0192_));
  AND_g _1886_ ( .A(1'h1), .B(_0327_), .Y(_0828_));
  NAND_g _1887_ ( .A(1'h1), .B(_0336_), .Y(_0829_));
  XNOR_g _1888_ ( .A(1'h1), .B(_0335_), .Y(_0830_));
  NAND_g _1889_ ( .A(_0828_), .B(_0830_), .Y(_0831_));
  XOR_g _1890_ ( .A(_0828_), .B(_0830_), .Y(_0832_));
  NAND_g _1891_ ( .A(_0301_), .B(_0832_), .Y(_0833_));
  NAND_g _1892_ ( .A(T3yp[1]), .B(_0239_), .Y(_0834_));
  NAND_g _1893_ ( .A(T3y[1]), .B(1'h1), .Y(_0835_));
  XOR_g _1894_ ( .A(T3y[1]), .B(1'h1), .Y(_0836_));
  XNOR_g _1895_ ( .A(T3y[1]), .B(1'h1), .Y(_0837_));
  NAND_g _1896_ ( .A(_0815_), .B(_0836_), .Y(_0838_));
  XNOR_g _1897_ ( .A(_0815_), .B(_0837_), .Y(_0839_));
  NAND_g _1898_ ( .A(_0381_), .B(_0839_), .Y(_0840_));
  NAND_g _1899_ ( .A(T3x[1]), .B(1'h1), .Y(_0841_));
  XOR_g _1900_ ( .A(T3x[1]), .B(1'h1), .Y(_0842_));
  XNOR_g _1901_ ( .A(T3x[1]), .B(1'h1), .Y(_0843_));
  NAND_g _1902_ ( .A(_0821_), .B(_0842_), .Y(_0844_));
  XNOR_g _1903_ ( .A(_0821_), .B(_0843_), .Y(_0845_));
  NAND_g _1904_ ( .A(_0265_), .B(_0845_), .Y(_0846_));
  NAND_g _1905_ ( .A(_0816_), .B(_0837_), .Y(_0847_));
  XNOR_g _1906_ ( .A(_0816_), .B(_0836_), .Y(_0848_));
  NAND_g _1907_ ( .A(_0262_), .B(_0848_), .Y(_0849_));
  NAND_g _1908_ ( .A(_0254_), .B(_0296_), .Y(_0850_));
  NAND_g _1909_ ( .A(T3x[0]), .B(_0233_), .Y(_0851_));
  NAND_g _1910_ ( .A(_0843_), .B(_0851_), .Y(_0852_));
  XNOR_g _1911_ ( .A(_0842_), .B(_0851_), .Y(_0853_));
  NAND_g _1912_ ( .A(_0850_), .B(_0853_), .Y(_0854_));
  AND_g _1913_ ( .A(_0834_), .B(_0849_), .Y(_0855_));
  AND_g _1914_ ( .A(_0846_), .B(_0854_), .Y(_0856_));
  AND_g _1915_ ( .A(_0855_), .B(_0856_), .Y(_0857_));
  AND_g _1916_ ( .A(_0840_), .B(_0857_), .Y(_0858_));
  NAND_g _1917_ ( .A(_0833_), .B(_0858_), .Y(_0193_));
  NAND_g _1918_ ( .A(_0829_), .B(_0831_), .Y(_0859_));
  NAND_g _1919_ ( .A(1'h0), .B(_0342_), .Y(_0860_));
  XNOR_g _1920_ ( .A(1'h0), .B(_0343_), .Y(_0861_));
  NAND_g _1921_ ( .A(_0859_), .B(_0861_), .Y(_0862_));
  XOR_g _1922_ ( .A(_0859_), .B(_0861_), .Y(_0863_));
  NAND_g _1923_ ( .A(_0301_), .B(_0863_), .Y(_0864_));
  NAND_g _1924_ ( .A(T3x[2]), .B(1'h0), .Y(_0865_));
  XOR_g _1925_ ( .A(T3x[2]), .B(1'h0), .Y(_0866_));
  XNOR_g _1926_ ( .A(T3x[2]), .B(1'h0), .Y(_0867_));
  AND_g _1927_ ( .A(_0841_), .B(_0844_), .Y(_0868_));
  NAND_g _1928_ ( .A(_0841_), .B(_0844_), .Y(_0869_));
  NAND_g _1929_ ( .A(_0866_), .B(_0869_), .Y(_0870_));
  NAND_g _1930_ ( .A(_0867_), .B(_0868_), .Y(_0871_));
  AND_g _1931_ ( .A(_0265_), .B(_0871_), .Y(_0872_));
  NAND_g _1932_ ( .A(_0870_), .B(_0872_), .Y(_0873_));
  NAND_g _1933_ ( .A(T3yp[2]), .B(_0239_), .Y(_0874_));
  AND_g _1934_ ( .A(_0873_), .B(_0874_), .Y(_0875_));
  NAND_g _1935_ ( .A(_0222_), .B(1'h1), .Y(_0876_));
  NAND_g _1936_ ( .A(_0852_), .B(_0876_), .Y(_0877_));
  NAND_g _1937_ ( .A(_0867_), .B(_0877_), .Y(_0878_));
  XNOR_g _1938_ ( .A(_0866_), .B(_0877_), .Y(_0879_));
  NAND_g _1939_ ( .A(_0850_), .B(_0879_), .Y(_0880_));
  NAND_g _1940_ ( .A(T3y[2]), .B(1'h0), .Y(_0881_));
  XOR_g _1941_ ( .A(T3y[2]), .B(1'h0), .Y(_0882_));
  XNOR_g _1942_ ( .A(T3y[2]), .B(1'h0), .Y(_0883_));
  NAND_g _1943_ ( .A(_0214_), .B(1'h1), .Y(_0884_));
  NAND_g _1944_ ( .A(_0847_), .B(_0884_), .Y(_0885_));
  NAND_g _1945_ ( .A(_0883_), .B(_0885_), .Y(_0886_));
  XNOR_g _1946_ ( .A(_0882_), .B(_0885_), .Y(_0887_));
  NAND_g _1947_ ( .A(_0262_), .B(_0887_), .Y(_0888_));
  AND_g _1948_ ( .A(_0835_), .B(_0838_), .Y(_0889_));
  NAND_g _1949_ ( .A(_0835_), .B(_0838_), .Y(_0890_));
  NAND_g _1950_ ( .A(_0883_), .B(_0889_), .Y(_0891_));
  NAND_g _1951_ ( .A(_0882_), .B(_0890_), .Y(_0892_));
  AND_g _1952_ ( .A(_0381_), .B(_0892_), .Y(_0893_));
  NAND_g _1953_ ( .A(_0891_), .B(_0893_), .Y(_0894_));
  AND_g _1954_ ( .A(_0888_), .B(_0894_), .Y(_0895_));
  AND_g _1955_ ( .A(_0880_), .B(_0895_), .Y(_0896_));
  AND_g _1956_ ( .A(_0875_), .B(_0896_), .Y(_0897_));
  NAND_g _1957_ ( .A(_0864_), .B(_0897_), .Y(_0194_));
  NAND_g _1958_ ( .A(_0860_), .B(_0862_), .Y(_0898_));
  NOR_g _1959_ ( .A(_0234_), .B(_0349_), .Y(_0899_));
  AND_g _1960_ ( .A(_0234_), .B(_0349_), .Y(_0900_));
  XNOR_g _1961_ ( .A(_0234_), .B(_0349_), .Y(_0901_));
  XNOR_g _1962_ ( .A(_0898_), .B(_0901_), .Y(_0902_));
  NAND_g _1963_ ( .A(_0301_), .B(_0902_), .Y(_0903_));
  NAND_g _1964_ ( .A(_0224_), .B(_0234_), .Y(_0904_));
  NAND_g _1965_ ( .A(T3x[3]), .B(1'h1), .Y(_0905_));
  XOR_g _1966_ ( .A(T3x[3]), .B(1'h1), .Y(_0906_));
  NAND_g _1967_ ( .A(_0223_), .B(1'h0), .Y(_0907_));
  NAND_g _1968_ ( .A(_0878_), .B(_0907_), .Y(_0908_));
  NOT_g _1969_ ( .A(_0908_), .Y(_0909_));
  NAND_g _1970_ ( .A(_0850_), .B(_0908_), .Y(_0910_));
  AND_g _1971_ ( .A(_0865_), .B(_0870_), .Y(_0911_));
  NOT_g _1972_ ( .A(_0911_), .Y(_0912_));
  NAND_g _1973_ ( .A(_0265_), .B(_0911_), .Y(_0913_));
  NAND_g _1974_ ( .A(_0910_), .B(_0913_), .Y(_0914_));
  NAND_g _1975_ ( .A(_0906_), .B(_0914_), .Y(_0915_));
  NAND_g _1976_ ( .A(T3yp[3]), .B(_0239_), .Y(_0916_));
  NAND_g _1977_ ( .A(_0216_), .B(_0234_), .Y(_0917_));
  NAND_g _1978_ ( .A(T3y[3]), .B(1'h1), .Y(_0918_));
  XOR_g _1979_ ( .A(T3y[3]), .B(1'h1), .Y(_0919_));
  NAND_g _1980_ ( .A(_0215_), .B(1'h0), .Y(_0920_));
  NAND_g _1981_ ( .A(_0886_), .B(_0920_), .Y(_0921_));
  NOT_g _1982_ ( .A(_0921_), .Y(_0922_));
  NAND_g _1983_ ( .A(_0262_), .B(_0922_), .Y(_0923_));
  AND_g _1984_ ( .A(_0881_), .B(_0892_), .Y(_0924_));
  NOT_g _1985_ ( .A(_0924_), .Y(_0925_));
  NAND_g _1986_ ( .A(_0381_), .B(_0925_), .Y(_0926_));
  AND_g _1987_ ( .A(_0923_), .B(_0926_), .Y(_0927_));
  NOR_g _1988_ ( .A(_0919_), .B(_0927_), .Y(_0928_));
  NAND_g _1989_ ( .A(_0850_), .B(_0909_), .Y(_0929_));
  NAND_g _1990_ ( .A(_0265_), .B(_0912_), .Y(_0930_));
  AND_g _1991_ ( .A(_0929_), .B(_0930_), .Y(_0931_));
  NOR_g _1992_ ( .A(_0906_), .B(_0931_), .Y(_0932_));
  NAND_g _1993_ ( .A(_0262_), .B(_0921_), .Y(_0933_));
  NAND_g _1994_ ( .A(_0381_), .B(_0924_), .Y(_0934_));
  NAND_g _1995_ ( .A(_0933_), .B(_0934_), .Y(_0935_));
  NAND_g _1996_ ( .A(_0919_), .B(_0935_), .Y(_0936_));
  NOR_g _1997_ ( .A(_0928_), .B(_0932_), .Y(_0937_));
  AND_g _1998_ ( .A(_0916_), .B(_0936_), .Y(_0938_));
  AND_g _1999_ ( .A(_0915_), .B(_0938_), .Y(_0939_));
  AND_g _2000_ ( .A(_0937_), .B(_0939_), .Y(_0940_));
  NAND_g _2001_ ( .A(_0903_), .B(_0940_), .Y(_0195_));
  NAND_g _2002_ ( .A(1'h1), .B(_0355_), .Y(_0941_));
  XNOR_g _2003_ ( .A(1'h1), .B(_0356_), .Y(_0942_));
  NOR_g _2004_ ( .A(_0898_), .B(_0899_), .Y(_0943_));
  NOR_g _2005_ ( .A(_0900_), .B(_0943_), .Y(_0944_));
  NAND_g _2006_ ( .A(_0942_), .B(_0944_), .Y(_0945_));
  XOR_g _2007_ ( .A(_0942_), .B(_0944_), .Y(_0946_));
  NAND_g _2008_ ( .A(_0301_), .B(_0946_), .Y(_0947_));
  NAND_g _2009_ ( .A(T3x[4]), .B(1'h1), .Y(_0948_));
  XOR_g _2010_ ( .A(T3x[4]), .B(1'h1), .Y(_0949_));
  XNOR_g _2011_ ( .A(T3x[4]), .B(1'h1), .Y(_0950_));
  NAND_g _2012_ ( .A(T3x[3]), .B(_0234_), .Y(_0951_));
  NAND_g _2013_ ( .A(_0224_), .B(1'h1), .Y(_0952_));
  NAND_g _2014_ ( .A(_0908_), .B(_0951_), .Y(_0953_));
  NAND_g _2015_ ( .A(_0952_), .B(_0953_), .Y(_0954_));
  NAND_g _2016_ ( .A(_0950_), .B(_0954_), .Y(_0955_));
  XNOR_g _2017_ ( .A(_0949_), .B(_0954_), .Y(_0956_));
  NAND_g _2018_ ( .A(_0850_), .B(_0956_), .Y(_0957_));
  NAND_g _2019_ ( .A(T3y[4]), .B(1'h1), .Y(_0958_));
  XOR_g _2020_ ( .A(T3y[4]), .B(1'h1), .Y(_0959_));
  XNOR_g _2021_ ( .A(T3y[4]), .B(1'h1), .Y(_0960_));
  NAND_g _2022_ ( .A(T3y[3]), .B(_0234_), .Y(_0961_));
  NAND_g _2023_ ( .A(_0216_), .B(1'h1), .Y(_0962_));
  NAND_g _2024_ ( .A(_0921_), .B(_0961_), .Y(_0963_));
  NAND_g _2025_ ( .A(_0962_), .B(_0963_), .Y(_0964_));
  NAND_g _2026_ ( .A(_0960_), .B(_0964_), .Y(_0965_));
  XNOR_g _2027_ ( .A(_0959_), .B(_0964_), .Y(_0966_));
  NAND_g _2028_ ( .A(_0262_), .B(_0966_), .Y(_0967_));
  AND_g _2029_ ( .A(_0957_), .B(_0967_), .Y(_0968_));
  NAND_g _2030_ ( .A(_0905_), .B(_0911_), .Y(_0969_));
  AND_g _2031_ ( .A(_0904_), .B(_0969_), .Y(_0970_));
  NOR_g _2032_ ( .A(_0949_), .B(_0970_), .Y(_0971_));
  NAND_g _2033_ ( .A(_0949_), .B(_0970_), .Y(_0972_));
  NAND_g _2034_ ( .A(_0265_), .B(_0972_), .Y(_0973_));
  NOR_g _2035_ ( .A(_0971_), .B(_0973_), .Y(_0974_));
  NAND_g _2036_ ( .A(T3yp[4]), .B(_0239_), .Y(_0975_));
  NAND_g _2037_ ( .A(_0918_), .B(_0924_), .Y(_0976_));
  AND_g _2038_ ( .A(_0917_), .B(_0976_), .Y(_0977_));
  NOR_g _2039_ ( .A(_0959_), .B(_0977_), .Y(_0978_));
  NAND_g _2040_ ( .A(_0959_), .B(_0977_), .Y(_0979_));
  NOR_g _2041_ ( .A(_0382_), .B(_0978_), .Y(_0980_));
  NAND_g _2042_ ( .A(_0979_), .B(_0980_), .Y(_0981_));
  NAND_g _2043_ ( .A(_0975_), .B(_0981_), .Y(_0982_));
  NOR_g _2044_ ( .A(_0974_), .B(_0982_), .Y(_0983_));
  AND_g _2045_ ( .A(_0968_), .B(_0983_), .Y(_0984_));
  NAND_g _2046_ ( .A(_0947_), .B(_0984_), .Y(_0196_));
  NAND_g _2047_ ( .A(_0941_), .B(_0945_), .Y(_0985_));
  NOR_g _2048_ ( .A(_0235_), .B(_0359_), .Y(_0986_));
  NAND_g _2049_ ( .A(_0235_), .B(_0359_), .Y(_0987_));
  XNOR_g _2050_ ( .A(_0235_), .B(_0359_), .Y(_0988_));
  XNOR_g _2051_ ( .A(_0985_), .B(_0988_), .Y(_0989_));
  NAND_g _2052_ ( .A(_0301_), .B(_0989_), .Y(_0990_));
  NAND_g _2053_ ( .A(_0226_), .B(_0235_), .Y(_0991_));
  NAND_g _2054_ ( .A(T3x[5]), .B(1'h1), .Y(_0992_));
  XOR_g _2055_ ( .A(T3x[5]), .B(1'h1), .Y(_0993_));
  AND_g _2056_ ( .A(_0948_), .B(_0972_), .Y(_0994_));
  XNOR_g _2057_ ( .A(_0993_), .B(_0994_), .Y(_0995_));
  NAND_g _2058_ ( .A(_0265_), .B(_0995_), .Y(_0996_));
  NAND_g _2059_ ( .A(T3yp[5]), .B(_0239_), .Y(_0997_));
  NAND_g _2060_ ( .A(T3y[5]), .B(_0235_), .Y(_0998_));
  NAND_g _2061_ ( .A(_0218_), .B(1'h1), .Y(_0999_));
  NAND_g _2062_ ( .A(_0218_), .B(_0235_), .Y(_1000_));
  NAND_g _2063_ ( .A(T3y[5]), .B(1'h1), .Y(_1001_));
  XOR_g _2064_ ( .A(T3y[5]), .B(1'h1), .Y(_1002_));
  AND_g _2065_ ( .A(_0958_), .B(_0979_), .Y(_1003_));
  XNOR_g _2066_ ( .A(_1002_), .B(_1003_), .Y(_1004_));
  NAND_g _2067_ ( .A(_0381_), .B(_1004_), .Y(_1005_));
  AND_g _2068_ ( .A(_0997_), .B(_1005_), .Y(_1006_));
  AND_g _2069_ ( .A(_0996_), .B(_1006_), .Y(_1007_));
  NAND_g _2070_ ( .A(_0225_), .B(1'h1), .Y(_1008_));
  AND_g _2071_ ( .A(_0955_), .B(_1008_), .Y(_1009_));
  XOR_g _2072_ ( .A(_0993_), .B(_1009_), .Y(_1010_));
  NAND_g _2073_ ( .A(_0850_), .B(_1010_), .Y(_1011_));
  NAND_g _2074_ ( .A(_0217_), .B(1'h1), .Y(_1012_));
  NAND_g _2075_ ( .A(_0965_), .B(_1012_), .Y(_1013_));
  XNOR_g _2076_ ( .A(_1002_), .B(_1013_), .Y(_1014_));
  NAND_g _2077_ ( .A(_0262_), .B(_1014_), .Y(_1015_));
  AND_g _2078_ ( .A(_1011_), .B(_1015_), .Y(_1016_));
  AND_g _2079_ ( .A(_1007_), .B(_1016_), .Y(_1017_));
  NAND_g _2080_ ( .A(_0990_), .B(_1017_), .Y(_0197_));
  AND_g _2081_ ( .A(_0985_), .B(_0987_), .Y(_1018_));
  NOR_g _2082_ ( .A(_0986_), .B(_1018_), .Y(_1019_));
  XNOR_g _2083_ ( .A(1'h0), .B(_1019_), .Y(_1020_));
  NAND_g _2084_ ( .A(_0301_), .B(_1020_), .Y(_1021_));
  NAND_g _2085_ ( .A(_1001_), .B(_1003_), .Y(_1022_));
  AND_g _2086_ ( .A(_1000_), .B(_1022_), .Y(_1023_));
  XNOR_g _2087_ ( .A(T3y[6]), .B(1'h0), .Y(_1024_));
  XNOR_g _2088_ ( .A(_1023_), .B(_1024_), .Y(_1025_));
  NAND_g _2089_ ( .A(_0381_), .B(_1025_), .Y(_1026_));
  NAND_g _2090_ ( .A(T3yp[6]), .B(_0239_), .Y(_1027_));
  AND_g _2091_ ( .A(_1026_), .B(_1027_), .Y(_1028_));
  XOR_g _2092_ ( .A(T3x[6]), .B(1'h0), .Y(_1029_));
  NAND_g _2093_ ( .A(_0992_), .B(_0994_), .Y(_1030_));
  AND_g _2094_ ( .A(_0991_), .B(_1030_), .Y(_1031_));
  NAND_g _2095_ ( .A(_1029_), .B(_1031_), .Y(_1032_));
  NOR_g _2096_ ( .A(_1029_), .B(_1031_), .Y(_1033_));
  NAND_g _2097_ ( .A(_0265_), .B(_1032_), .Y(_1034_));
  NOR_g _2098_ ( .A(_1033_), .B(_1034_), .Y(_1035_));
  NAND_g _2099_ ( .A(_0998_), .B(_1013_), .Y(_1036_));
  AND_g _2100_ ( .A(_0999_), .B(_1036_), .Y(_1037_));
  XNOR_g _2101_ ( .A(_1024_), .B(_1037_), .Y(_0199_));
  NAND_g _2102_ ( .A(_0262_), .B(_0199_), .Y(_0200_));
  NAND_g _2103_ ( .A(_0226_), .B(1'h1), .Y(_0201_));
  NAND_g _2104_ ( .A(T3x[5]), .B(_0235_), .Y(_0202_));
  NAND_g _2105_ ( .A(_1009_), .B(_0201_), .Y(_0203_));
  AND_g _2106_ ( .A(_0202_), .B(_0203_), .Y(_0204_));
  XNOR_g _2107_ ( .A(_1029_), .B(_0204_), .Y(_0205_));
  AND_g _2108_ ( .A(_0850_), .B(_0205_), .Y(_0206_));
  NOR_g _2109_ ( .A(_1035_), .B(_0206_), .Y(_0207_));
  AND_g _2110_ ( .A(_0200_), .B(_0207_), .Y(_0208_));
  AND_g _2111_ ( .A(_1028_), .B(_0208_), .Y(_0209_));
  NAND_g _2112_ ( .A(_1021_), .B(_0209_), .Y(_0198_));
  NOT_g _2113_ ( .A(KEY_N[3]), .Y(_0150_));
  NOT_g _2114_ ( .A(KEY_N[3]), .Y(_0151_));
  NOT_g _2115_ ( .A(KEY_N[3]), .Y(_0152_));
  DFFRcell _2116_ ( .C(CLOCK_50), .D(_0153_), .Q(T3state[0]), .R(_0149_));
  DFFRcell _2117_ ( .C(CLOCK_50), .D(_0154_), .Q(T3state[1]), .R(_0150_));
  DFFRcell _2118_ ( .C(CLOCK_50), .D(_0155_), .Q(T3state[2]), .R(_0151_));
  DFFRcell _2119_ ( .C(CLOCK_50), .D(_0156_), .Q(T3state[3]), .R(_0152_));
  DFFcell _2120_ ( .C(CLOCK_50), .D(_0157_), .Q(T3y[0]));
  DFFcell _2121_ ( .C(CLOCK_50), .D(_0158_), .Q(T3y[1]));
  DFFcell _2122_ ( .C(CLOCK_50), .D(_0159_), .Q(T3y[2]));
  DFFcell _2123_ ( .C(CLOCK_50), .D(_0160_), .Q(T3y[3]));
  DFFcell _2124_ ( .C(CLOCK_50), .D(_0161_), .Q(T3y[4]));
  DFFcell _2125_ ( .C(CLOCK_50), .D(_0162_), .Q(T3y[5]));
  DFFcell _2126_ ( .C(CLOCK_50), .D(_0163_), .Q(T3y[6]));
  DFFcell _2127_ ( .C(CLOCK_50), .D(_0164_), .Q(T3colourcircle[0]));
  DFFcell _2128_ ( .C(CLOCK_50), .D(_0165_), .Q(T3colourcircle[1]));
  DFFcell _2129_ ( .C(CLOCK_50), .D(_0166_), .Q(T3colourcircle[2]));
  DFFcell _2130_ ( .C(CLOCK_50), .D(_0167_), .Q(T3xp[0]));
  DFFcell _2131_ ( .C(CLOCK_50), .D(_0168_), .Q(T3xp[1]));
  DFFcell _2132_ ( .C(CLOCK_50), .D(_0169_), .Q(T3xp[2]));
  DFFcell _2133_ ( .C(CLOCK_50), .D(_0170_), .Q(T3xp[3]));
  DFFcell _2134_ ( .C(CLOCK_50), .D(_0171_), .Q(T3xp[4]));
  DFFcell _2135_ ( .C(CLOCK_50), .D(_0172_), .Q(T3xp[5]));
  DFFcell _2136_ ( .C(CLOCK_50), .D(_0173_), .Q(T3xp[6]));
  DFFcell _2137_ ( .C(CLOCK_50), .D(_0174_), .Q(T3xp[7]));
  DFFcell _2138_ ( .C(CLOCK_50), .D(_0175_), .Q(T3d[0]));
  DFFcell _2139_ ( .C(CLOCK_50), .D(_0176_), .Q(T3d[1]));
  DFFcell _2140_ ( .C(CLOCK_50), .D(_0177_), .Q(T3d[2]));
  DFFcell _2141_ ( .C(CLOCK_50), .D(_0178_), .Q(T3d[3]));
  DFFcell _2142_ ( .C(CLOCK_50), .D(_0179_), .Q(T3d[4]));
  DFFcell _2143_ ( .C(CLOCK_50), .D(_0180_), .Q(T3d[5]));
  DFFcell _2144_ ( .C(CLOCK_50), .D(_0181_), .Q(T3d[6]));
  DFFcell _2145_ ( .C(CLOCK_50), .D(_0182_), .Q(T3d[7]));
  DFFcell _2146_ ( .C(CLOCK_50), .D(_0183_), .Q(T3d[8]));
  DFFcell _2147_ ( .C(CLOCK_50), .D(_0184_), .Q(T3x[0]));
  DFFcell _2148_ ( .C(CLOCK_50), .D(_0185_), .Q(T3x[1]));
  DFFcell _2149_ ( .C(CLOCK_50), .D(_0186_), .Q(T3x[2]));
  DFFcell _2150_ ( .C(CLOCK_50), .D(_0187_), .Q(T3x[3]));
  DFFcell _2151_ ( .C(CLOCK_50), .D(_0188_), .Q(T3x[4]));
  DFFcell _2152_ ( .C(CLOCK_50), .D(_0189_), .Q(T3x[5]));
  DFFcell _2153_ ( .C(CLOCK_50), .D(_0190_), .Q(T3x[6]));
  DFFcell _2154_ ( .C(CLOCK_50), .D(_0191_), .Q(T3x[7]));
  DFFcell _2155_ ( .C(CLOCK_50), .D(_0192_), .Q(T3yp[0]));
  DFFcell _2156_ ( .C(CLOCK_50), .D(_0193_), .Q(T3yp[1]));
  DFFcell _2157_ ( .C(CLOCK_50), .D(_0194_), .Q(T3yp[2]));
  DFFcell _2158_ ( .C(CLOCK_50), .D(_0195_), .Q(T3yp[3]));
  DFFcell _2159_ ( .C(CLOCK_50), .D(_0196_), .Q(T3yp[4]));
  DFFcell _2160_ ( .C(CLOCK_50), .D(_0197_), .Q(T3yp[5]));
  DFFcell _2161_ ( .C(CLOCK_50), .D(_0198_), .Q(T3yp[6]));
endmodule
