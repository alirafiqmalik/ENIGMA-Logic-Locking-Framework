module locked(inputs,key,lockingkeyinput,out);
input [7:0] inputs;
input [7:0] key;
input [255:0] lockingkeyinput;
output [1:0] out;
wire _017_;
wire _068_;
wire _071_;
wire _021_;
wire _009_;
wire _058_;
wire _007_;
wire _064_;
wire _027_;
wire _046_;
wire _035_;
wire _038_;
wire _029_;
wire _033_;
wire _061_;
wire _052_;
wire _054_;
wire _036_;
wire _002_;
wire _040_;
wire _059_;
wire _028_;
wire _034_;
wire _056_;
wire _000_;
wire _006_;
wire _010_;
wire _057_;
wire _008_;
wire _065_;
wire _043_;
wire _031_;
wire _055_;
wire _013_;
wire _011_;
wire _005_;
wire _026_;
wire _067_;
wire [4:0] scc;
wire _045_;
wire _015_;
wire _019_;
wire _060_;
wire _023_;
wire _051_;
wire _024_;
wire _025_;
wire _004_;
wire _062_;
wire _069_;
wire _047_;
wire _012_;
wire _048_;
wire _003_;
wire _041_;
wire _042_;
wire _049_;
wire _020_;
wire _014_;
wire _032_;
wire _030_;
wire _070_;
wire _001_;
wire _066_;
wire _039_;
wire [4:0] s1cc;
wire _022_;
wire _016_;
wire _050_;
wire _044_;
wire _053_;
wire _063_;
wire _018_;
wire _037_;
wire keywire74;
wire keywire75;
wire keywire76;
wire keywire77;
wire keywire78;
wire keywire79;
wire keywire80;
wire keywire81;
wire keywire82;
wire keywire83;
wire keywire84;
wire keywire85;
wire keywire86;
wire keywire87;
wire keywire88;
wire keywire89;
wire keywire90;
wire keywire91;
wire keywire92;
wire keywire93;
wire keywire94;
wire keywire95;
wire keywire96;
wire keywire97;
wire keywire98;
wire keywire99;
wire keywire100;
wire keywire101;
wire keywire102;
wire keywire103;
wire keywire104;
wire keywire105;
wire keywire106;
wire keywire107;
wire keywire108;
wire keywire109;
wire keywire110;
wire keywire111;
wire keywire112;
wire keywire113;
wire keywire114;
wire keywire115;
wire keywire116;
wire keywire117;
wire keywire118;
wire keywire119;
wire keywire120;
wire keywire121;
wire keywire122;
wire keywire123;
wire keywire124;
wire keywire125;
wire keywire126;
wire keywire127;
wire keywire128;
wire keywire129;
wire keywire130;
wire keywire131;
wire keywire132;
wire keywire133;
wire keywire134;
wire keywire135;
wire keywire136;
wire keywire137;
wire keywire138;
wire keywire139;
wire keywire140;
wire keywire141;
wire keywire142;
wire keywire143;
wire keywire144;
wire keywire145;
wire keywire146;
wire keywire147;
wire keywire148;
wire keywire149;
wire keywire150;
wire keywire151;
wire keywire152;
wire keywire153;
wire keywire154;
wire keywire155;
wire keywire156;
wire keywire157;
wire keywire158;
wire keywire159;
wire keywire160;
wire keywire161;
wire keywire162;
wire keywire163;
wire keywire164;
wire keywire165;
wire keywire166;
wire keywire167;
wire keywire168;
wire keywire169;
wire keywire170;
wire keywire171;
wire keywire172;
wire keywire173;
wire keywire174;
wire keywire175;
wire keywire176;
wire keywire177;
wire keywire178;
wire keywire179;
wire keywire180;
wire keywire181;
wire keywire182;
wire keywire183;
wire keywire184;
wire keywire185;
wire keywire186;
wire keywire187;
wire keywire188;
wire keywire189;
wire keywire190;
wire keywire191;
wire keywire192;
wire keywire193;
wire keywire194;
wire keywire195;
wire keywire196;
wire keywire197;
wire keywire198;
wire keywire199;
wire keywire200;
wire keywire201;
wire keywire202;
wire keywire203;
wire keywire204;
wire keywire205;
wire keywire206;
wire keywire207;
wire keywire208;
wire keywire209;
wire keywire210;
wire keywire211;
wire keywire212;
wire keywire213;
wire keywire214;
wire keywire215;
wire keywire216;
wire keywire217;
wire keywire218;
wire keywire219;
wire keywire220;
wire keywire221;
wire keywire222;
wire keywire223;
wire keywire224;
wire keywire225;
wire keywire226;
wire keywire227;
wire keywire228;
wire keywire229;
wire keywire230;
wire keywire231;
wire keywire232;
wire keywire233;
wire keywire234;
wire keywire235;
wire keywire236;
wire keywire237;
wire keywire238;
wire keywire239;
wire keywire240;
wire keywire241;
wire keywire242;
wire keywire243;
wire keywire244;
wire keywire245;
wire keywire246;
wire keywire247;
wire keywire248;
wire keywire249;
wire keywire250;
wire keywire251;
wire keywire252;
wire keywire253;
wire keywire254;
wire keywire255;
wire keywire256;
wire keywire257;
wire keywire258;
wire keywire259;
wire keywire260;
wire keywire261;
wire keywire262;
wire keywire263;
wire keywire264;
wire keywire265;
wire keywire266;
wire keywire267;
wire keywire268;
wire keywire269;
wire keywire270;
wire keywire271;
wire keywire272;
wire keywire273;
wire keywire274;
wire keywire275;
wire keywire276;
wire keywire277;
wire keywire278;
wire keywire279;
wire keywire280;
wire keywire281;
wire keywire282;
wire keywire283;
wire keywire284;
wire keywire285;
wire keywire286;
wire keywire287;
wire keywire288;
wire keywire289;
wire keywire290;
wire keywire291;
wire keywire292;
wire keywire293;
wire keywire294;
wire keywire295;
wire keywire296;
wire keywire297;
wire keywire298;
wire keywire299;
wire keywire300;
wire keywire301;
wire keywire302;
wire keywire303;
wire keywire304;
wire keywire305;
wire keywire306;
wire keywire307;
wire keywire308;
wire keywire309;
wire keywire310;
wire keywire311;
wire keywire312;
wire keywire313;
wire keywire314;
wire keywire315;
wire keywire316;
wire keywire317;
wire keywire318;
wire keywire319;
wire keywire320;
wire keywire321;
wire keywire322;
wire keywire323;
wire keywire324;
wire keywire325;
wire keywire326;
wire keywire327;
wire keywire328;
wire keywire329;
NOT_g NOT_g_072_(.A(inputs[3]), .Y(keywire237));
NOT_g NOT_g_114_(.A(inputs[3]), .Y(keywire238));
XNOR_g XNOR_g_073_(.A(key[0]), .B(inputs[0]), .Y(keywire320));
XNOR_g XNOR_g_074_(.A(key[7]), .B(inputs[7]), .Y(keywire319));
XNOR_g XNOR_g_076_(.A(key[1]), .B(inputs[1]), .Y(keywire318));
XNOR_g XNOR_g_077_(.A(key[3]), .B(inputs[3]), .Y(keywire317));
XNOR_g XNOR_g_087_(.A(key[5]), .B(inputs[5]), .Y(keywire249));
XNOR_g XNOR_g_088_(.A(key[2]), .B(inputs[2]), .Y(keywire231));
XNOR_g XNOR_g_090_(.A(key[6]), .B(inputs[6]), .Y(keywire253));
XNOR_g XNOR_g_091_(.A(key[4]), .B(inputs[4]), .Y(keywire329));
XNOR_g XNOR_g_096_(.A(_023_), .B(scc[0]), .Y(keywire295));
XNOR_g XNOR_g_115_(.A(key[0]), .B(inputs[0]), .Y(keywire328));
XNOR_g XNOR_g_116_(.A(key[7]), .B(inputs[7]), .Y(keywire327));
XNOR_g XNOR_g_118_(.A(key[1]), .B(inputs[1]), .Y(keywire326));
XNOR_g XNOR_g_119_(.A(key[3]), .B(inputs[3]), .Y(keywire325));
XNOR_g XNOR_g_129_(.A(key[5]), .B(inputs[5]), .Y(keywire250));
XNOR_g XNOR_g_130_(.A(key[2]), .B(inputs[2]), .Y(keywire232));
XNOR_g XNOR_g_132_(.A(key[6]), .B(inputs[6]), .Y(keywire254));
XNOR_g XNOR_g_133_(.A(key[4]), .B(inputs[4]), .Y(keywire246));
XNOR_g XNOR_g_138_(.A(_059_), .B(s1cc[0]), .Y(keywire296));
XNOR_g keygate_XNOR_0(.A(keywire74), .B(lockingkeyinput[0]), .Y(_013_));
XNOR_g keygate_XNOR_2(.A(keywire76), .B(lockingkeyinput[2]), .Y(_022_));
XNOR_g keygate_XNOR_6(.A(keywire80), .B(lockingkeyinput[6]), .Y(_037_));
XNOR_g keygate_XNOR_7(.A(keywire81), .B(lockingkeyinput[7]), .Y(_012_));
XNOR_g keygate_XNOR_9(.A(keywire83), .B(lockingkeyinput[9]), .Y(_048_));
XNOR_g keygate_XNOR_14(.A(keywire88), .B(lockingkeyinput[14]), .Y(_040_));
XNOR_g keygate_XNOR_15(.A(keywire89), .B(lockingkeyinput[15]), .Y(_011_));
XNOR_g keygate_XNOR_16(.A(keywire90), .B(lockingkeyinput[16]), .Y(_047_));
XNOR_g keygate_XNOR_18(.A(keywire92), .B(lockingkeyinput[18]), .Y(_061_));
XNOR_g keygate_XNOR_19(.A(keywire93), .B(lockingkeyinput[19]), .Y(_026_));
XNOR_g keygate_XNOR_21(.A(keywire95), .B(lockingkeyinput[21]), .Y(_016_));
XNOR_g keygate_XNOR_22(.A(keywire96), .B(lockingkeyinput[22]), .Y(_052_));
XNOR_g keygate_XNOR_24(.A(keywire98), .B(lockingkeyinput[24]), .Y(_065_));
XNOR_g keygate_XNOR_25(.A(keywire99), .B(lockingkeyinput[25]), .Y(_030_));
XNOR_g keygate_XNOR_27(.A(keywire101), .B(lockingkeyinput[27]), .Y(_000_));
XNOR_g keygate_XNOR_28(.A(keywire102), .B(lockingkeyinput[28]), .Y(_036_));
XNOR_g keygate_XNOR_29(.A(keywire103), .B(lockingkeyinput[29]), .Y(_005_));
XNOR_g keygate_XNOR_30(.A(keywire104), .B(lockingkeyinput[30]), .Y(_041_));
XNOR_g keygate_XNOR_33(.A(keywire107), .B(lockingkeyinput[33]), .Y(_034_));
XNOR_g keygate_XNOR_34(.A(keywire108), .B(lockingkeyinput[34]), .Y(_070_));
XNOR_g keygate_XNOR_36(.A(keywire110), .B(lockingkeyinput[36]), .Y(_055_));
XNOR_g keygate_XNOR_39(.A(keywire113), .B(lockingkeyinput[39]), .Y(_015_));
XNOR_g keygate_XNOR_40(.A(keywire114), .B(lockingkeyinput[40]), .Y(_051_));
XNOR_g keygate_XNOR_41(.A(keywire115), .B(lockingkeyinput[41]), .Y(_008_));
XNOR_g keygate_XNOR_43(.A(keywire117), .B(lockingkeyinput[43]), .Y(_018_));
XNOR_g keygate_XNOR_45(.A(keywire119), .B(lockingkeyinput[45]), .Y(_002_));
XNOR_g keygate_XNOR_48(.A(keywire122), .B(lockingkeyinput[48]), .Y(_039_));
XNOR_g keygate_XNOR_49(.A(keywire123), .B(lockingkeyinput[49]), .Y(_027_));
XNOR_g keygate_XNOR_56(.A(keywire130), .B(lockingkeyinput[56]), .Y(_042_));
XNOR_g keygate_XNOR_58(.A(keywire132), .B(lockingkeyinput[58]), .Y(_064_));
XNOR_g keygate_XNOR_59(.A(keywire133), .B(lockingkeyinput[59]), .Y(_017_));
XNOR_g keygate_XNOR_60(.A(keywire134), .B(lockingkeyinput[60]), .Y(_053_));
XNOR_g keygate_XNOR_61(.A(keywire135), .B(lockingkeyinput[61]), .Y(_032_));
XNOR_g keygate_XNOR_62(.A(keywire136), .B(lockingkeyinput[62]), .Y(_068_));
XNOR_g keygate_XNOR_64(.A(keywire138), .B(lockingkeyinput[64]), .Y(scc[2]));
XNOR_g keygate_XNOR_65(.A(keywire139), .B(lockingkeyinput[65]), .Y(_067_));
XNOR_g keygate_XNOR_66(.A(keywire140), .B(lockingkeyinput[66]), .Y(s1cc[2]));
XNOR_g keygate_XNOR_69(.A(keywire143), .B(lockingkeyinput[69]), .Y(_035_));
XNOR_g keygate_XNOR_70(.A(keywire144), .B(lockingkeyinput[70]), .Y(scc[3]));
XNOR_g keygate_XNOR_72(.A(keywire146), .B(lockingkeyinput[72]), .Y(s1cc[3]));
XNOR_g keygate_XNOR_73(.A(keywire147), .B(lockingkeyinput[73]), .Y(_020_));
XNOR_g keygate_XNOR_74(.A(keywire148), .B(lockingkeyinput[74]), .Y(_056_));
XNOR_g keygate_XNOR_79(.A(keywire153), .B(lockingkeyinput[79]), .Y(_050_));
XNOR_g keygate_XNOR_82(.A(keywire156), .B(lockingkeyinput[82]), .Y(_059_));
XNOR_g keygate_XNOR_83(.A(keywire157), .B(lockingkeyinput[83]), .Y(_058_));
XNOR_g keygate_XNOR_86(.A(keywire160), .B(lockingkeyinput[86]), .Y(keywire128));
XNOR_g keygate_XNOR_87(.A(keywire161), .B(lockingkeyinput[87]), .Y(keywire77));
XNOR_g keygate_XNOR_88(.A(keywire162), .B(lockingkeyinput[88]), .Y(keywire85));
XNOR_g keygate_XNOR_90(.A(keywire164), .B(lockingkeyinput[90]), .Y(keywire86));
XNOR_g keygate_XNOR_91(.A(keywire165), .B(lockingkeyinput[91]), .Y(keywire76));
XNOR_g keygate_XNOR_95(.A(keywire169), .B(lockingkeyinput[95]), .Y(keywire154));
XNOR_g keygate_XNOR_96(.A(keywire170), .B(lockingkeyinput[96]), .Y(keywire75));
XNOR_g keygate_XNOR_97(.A(keywire171), .B(lockingkeyinput[97]), .Y(keywire129));
XNOR_g keygate_XNOR_98(.A(keywire172), .B(lockingkeyinput[98]), .Y(keywire121));
XNOR_g keygate_XNOR_99(.A(keywire173), .B(lockingkeyinput[99]), .Y(keywire155));
XNOR_g keygate_XNOR_102(.A(keywire176), .B(lockingkeyinput[102]), .Y(keywire122));
XNOR_g keygate_XNOR_103(.A(keywire177), .B(lockingkeyinput[103]), .Y(keywire147));
XNOR_g keygate_XNOR_104(.A(keywire178), .B(lockingkeyinput[104]), .Y(keywire133));
XNOR_g keygate_XNOR_106(.A(keywire180), .B(lockingkeyinput[106]), .Y(keywire149));
XNOR_g keygate_XNOR_108(.A(keywire182), .B(lockingkeyinput[108]), .Y(keywire87));
XNOR_g keygate_XNOR_109(.A(keywire183), .B(lockingkeyinput[109]), .Y(keywire119));
XNOR_g keygate_XNOR_113(.A(keywire187), .B(lockingkeyinput[113]), .Y(keywire125));
XNOR_g keygate_XNOR_115(.A(keywire189), .B(lockingkeyinput[115]), .Y(keywire104));
XNOR_g keygate_XNOR_116(.A(keywire190), .B(lockingkeyinput[116]), .Y(keywire88));
XNOR_g keygate_XNOR_119(.A(keywire193), .B(lockingkeyinput[119]), .Y(keywire109));
XNOR_g keygate_XNOR_121(.A(keywire195), .B(lockingkeyinput[121]), .Y(keywire95));
XNOR_g keygate_XNOR_124(.A(keywire198), .B(lockingkeyinput[124]), .Y(keywire111));
XNOR_g keygate_XNOR_128(.A(keywire202), .B(lockingkeyinput[128]), .Y(keywire96));
XNOR_g keygate_XNOR_129(.A(keywire203), .B(lockingkeyinput[129]), .Y(keywire114));
XNOR_g keygate_XNOR_131(.A(keywire205), .B(lockingkeyinput[131]), .Y(keywire90));
XNOR_g keygate_XNOR_133(.A(keywire207), .B(lockingkeyinput[133]), .Y(keywire116));
XNOR_g keygate_XNOR_136(.A(keywire210), .B(lockingkeyinput[136]), .Y(keywire179));
XNOR_g keygate_XNOR_137(.A(keywire211), .B(lockingkeyinput[137]), .Y(keywire170));
XNOR_g keygate_XNOR_139(.A(keywire213), .B(lockingkeyinput[139]), .Y(keywire161));
XNOR_g keygate_XNOR_141(.A(keywire215), .B(lockingkeyinput[141]), .Y(keywire184));
XNOR_g keygate_XNOR_142(.A(keywire216), .B(lockingkeyinput[142]), .Y(keywire192));
XNOR_g keygate_XNOR_143(.A(keywire217), .B(lockingkeyinput[143]), .Y(keywire197));
XNOR_g keygate_XNOR_145(.A(keywire219), .B(lockingkeyinput[145]), .Y(keywire204));
XNOR_g keygate_XNOR_147(.A(keywire221), .B(lockingkeyinput[147]), .Y(keywire162));
XNOR_g keygate_XNOR_148(.A(keywire222), .B(lockingkeyinput[148]), .Y(keywire164));
XNOR_g keygate_XNOR_149(.A(keywire223), .B(lockingkeyinput[149]), .Y(keywire182));
XNOR_g keygate_XNOR_150(.A(keywire224), .B(lockingkeyinput[150]), .Y(keywire190));
XNOR_g keygate_XNOR_151(.A(keywire225), .B(lockingkeyinput[151]), .Y(keywire158));
XNOR_g keygate_XNOR_152(.A(keywire226), .B(lockingkeyinput[152]), .Y(keywire205));
XNOR_g keygate_XNOR_153(.A(keywire227), .B(lockingkeyinput[153]), .Y(keywire91));
XNOR_g keygate_XNOR_155(.A(keywire229), .B(lockingkeyinput[155]), .Y(keywire93));
XNOR_g keygate_XNOR_157(.A(keywire231), .B(lockingkeyinput[157]), .Y(keywire195));
XNOR_g keygate_XNOR_158(.A(keywire232), .B(lockingkeyinput[158]), .Y(keywire202));
XNOR_g keygate_XNOR_160(.A(keywire234), .B(lockingkeyinput[160]), .Y(keywire98));
XNOR_g keygate_XNOR_162(.A(keywire236), .B(lockingkeyinput[162]), .Y(keywire100));
XNOR_g keygate_XNOR_164(.A(keywire238), .B(lockingkeyinput[164]), .Y(keywire209));
XNOR_g keygate_XNOR_165(.A(keywire239), .B(lockingkeyinput[165]), .Y(keywire181));
XNOR_g keygate_XNOR_169(.A(keywire243), .B(lockingkeyinput[169]), .Y(keywire107));
XNOR_g keygate_XNOR_170(.A(keywire244), .B(lockingkeyinput[170]), .Y(keywire108));
XNOR_g keygate_XNOR_174(.A(keywire248), .B(lockingkeyinput[174]), .Y(keywire206));
XNOR_g keygate_XNOR_175(.A(keywire249), .B(lockingkeyinput[175]), .Y(keywire196));
XNOR_g keygate_XNOR_176(.A(keywire250), .B(lockingkeyinput[176]), .Y(keywire203));
XNOR_g keygate_XNOR_177(.A(keywire251), .B(lockingkeyinput[177]), .Y(keywire199));
XNOR_g keygate_XNOR_178(.A(keywire252), .B(lockingkeyinput[178]), .Y(keywire207));
XNOR_g keygate_XNOR_179(.A(keywire253), .B(lockingkeyinput[179]), .Y(keywire194));
XNOR_g keygate_XNOR_180(.A(keywire254), .B(lockingkeyinput[180]), .Y(keywire201));
XNOR_g keygate_XNOR_181(.A(keywire255), .B(lockingkeyinput[181]), .Y(keywire183));
XNOR_g keygate_XNOR_183(.A(keywire257), .B(lockingkeyinput[183]), .Y(keywire172));
XNOR_g keygate_XNOR_184(.A(keywire258), .B(lockingkeyinput[184]), .Y(keywire176));
XNOR_g keygate_XNOR_186(.A(keywire260), .B(lockingkeyinput[186]), .Y(keywire124));
XNOR_g keygate_XNOR_187(.A(keywire261), .B(lockingkeyinput[187]), .Y(keywire187));
XNOR_g keygate_XNOR_190(.A(keywire264), .B(lockingkeyinput[190]), .Y(keywire160));
XNOR_g keygate_XNOR_195(.A(keywire269), .B(lockingkeyinput[195]), .Y(keywire178));
XNOR_g keygate_XNOR_199(.A(keywire273), .B(lockingkeyinput[199]), .Y(keywire137));
XNOR_g keygate_XNOR_200(.A(keywire274), .B(lockingkeyinput[200]), .Y(keywire138));
XNOR_g keygate_XNOR_201(.A(keywire275), .B(lockingkeyinput[201]), .Y(keywire139));
XNOR_g keygate_XNOR_202(.A(keywire276), .B(lockingkeyinput[202]), .Y(keywire140));
XNOR_g keygate_XNOR_204(.A(keywire278), .B(lockingkeyinput[204]), .Y(keywire142));
XNOR_g keygate_XNOR_207(.A(keywire281), .B(lockingkeyinput[207]), .Y(keywire145));
XNOR_g keygate_XNOR_208(.A(keywire282), .B(lockingkeyinput[208]), .Y(keywire146));
XNOR_g keygate_XNOR_209(.A(keywire283), .B(lockingkeyinput[209]), .Y(keywire177));
XNOR_g keygate_XNOR_211(.A(keywire285), .B(lockingkeyinput[211]), .Y(keywire180));
XNOR_g keygate_XNOR_215(.A(keywire289), .B(lockingkeyinput[215]), .Y(keywire174));
XNOR_g keygate_XNOR_217(.A(keywire291), .B(lockingkeyinput[217]), .Y(keywire173));
XNOR_g keygate_XNOR_218(.A(keywire292), .B(lockingkeyinput[218]), .Y(keywire163));
XNOR_g keygate_XNOR_219(.A(keywire293), .B(lockingkeyinput[219]), .Y(keywire167));
XNOR_g keygate_XNOR_223(.A(keywire297), .B(lockingkeyinput[223]), .Y(keywire213));
XNOR_g keygate_XNOR_224(.A(keywire298), .B(lockingkeyinput[224]), .Y(keywire221));
XNOR_g keygate_XNOR_226(.A(keywire300), .B(lockingkeyinput[226]), .Y(keywire222));
XNOR_g keygate_XNOR_227(.A(keywire301), .B(lockingkeyinput[227]), .Y(keywire212));
XNOR_g keygate_XNOR_229(.A(keywire303), .B(lockingkeyinput[229]), .Y(keywire293));
XNOR_g keygate_XNOR_231(.A(keywire305), .B(lockingkeyinput[231]), .Y(keywire290));
XNOR_g keygate_XNOR_232(.A(keywire306), .B(lockingkeyinput[232]), .Y(keywire211));
XNOR_g keygate_XNOR_233(.A(keywire307), .B(lockingkeyinput[233]), .Y(keywire265));
XNOR_g keygate_XNOR_236(.A(keywire310), .B(lockingkeyinput[236]), .Y(keywire289));
XNOR_g keygate_XNOR_244(.A(keywire318), .B(lockingkeyinput[244]), .Y(keywire223));
XNOR_g keygate_XNOR_245(.A(keywire319), .B(lockingkeyinput[245]), .Y(keywire255));
XNOR_g keygate_XNOR_246(.A(keywire320), .B(lockingkeyinput[246]), .Y(keywire215));
XNOR_g keygate_XNOR_247(.A(keywire321), .B(lockingkeyinput[247]), .Y(keywire284));
XNOR_g keygate_XNOR_248(.A(keywire322), .B(lockingkeyinput[248]), .Y(keywire270));
XNOR_g keygate_XNOR_252(.A(keywire326), .B(lockingkeyinput[252]), .Y(keywire224));
XNOR_g keygate_XNOR_254(.A(keywire328), .B(lockingkeyinput[254]), .Y(keywire216));
AND_g AND_g_075_(.A(_002_), .B(_001_), .Y(keywire308));
AND_g AND_g_078_(.A(_005_), .B(_004_), .Y(keywire307));
AND_g AND_g_079_(.A(_006_), .B(_003_), .Y(keywire302));
AND_g AND_g_082_(.A(_009_), .B(_008_), .Y(keywire316));
AND_g AND_g_084_(.A(_000_), .B(inputs[0]), .Y(keywire217));
AND_g AND_g_085_(.A(_012_), .B(_011_), .Y(keywire315));
AND_g AND_g_089_(.A(_016_), .B(_015_), .Y(keywire314));
AND_g AND_g_092_(.A(_019_), .B(_018_), .Y(keywire313));
AND_g AND_g_093_(.A(_020_), .B(_017_), .Y(keywire305));
AND_g AND_g_094_(.A(_021_), .B(_014_), .Y(keywire301));
AND_g AND_g_097_(.A(inputs[4]), .B(inputs[0]), .Y(keywire218));
AND_g AND_g_117_(.A(_038_), .B(_037_), .Y(keywire312));
AND_g AND_g_120_(.A(_041_), .B(_040_), .Y(keywire311));
AND_g AND_g_121_(.A(_042_), .B(_039_), .Y(keywire304));
AND_g AND_g_124_(.A(_045_), .B(_044_), .Y(keywire324));
AND_g AND_g_126_(.A(_036_), .B(inputs[0]), .Y(keywire219));
AND_g AND_g_127_(.A(_048_), .B(_047_), .Y(keywire323));
AND_g AND_g_131_(.A(_052_), .B(_051_), .Y(keywire322));
AND_g AND_g_134_(.A(_055_), .B(_054_), .Y(keywire321));
AND_g AND_g_135_(.A(_056_), .B(_053_), .Y(keywire309));
AND_g AND_g_136_(.A(_057_), .B(_050_), .Y(keywire303));
AND_g AND_g_139_(.A(inputs[4]), .B(inputs[0]), .Y(keywire220));
NOR_g NOR_g_080_(.A(inputs[6]), .B(inputs[5]), .Y(keywire251));
NOR_g NOR_g_081_(.A(inputs[7]), .B(inputs[4]), .Y(keywire247));
NOR_g NOR_g_083_(.A(inputs[2]), .B(inputs[1]), .Y(keywire294));
NOR_g NOR_g_122_(.A(inputs[6]), .B(inputs[5]), .Y(keywire252));
NOR_g NOR_g_123_(.A(inputs[7]), .B(inputs[4]), .Y(keywire248));
NOR_g NOR_g_125_(.A(inputs[2]), .B(inputs[1]), .Y(keywire226));
NAND_g NAND_g_086_(.A(_013_), .B(_010_), .Y(keywire306));
NAND_g NAND_g_095_(.A(_022_), .B(_007_), .Y(keywire297));
NAND_g NAND_g_098_(.A(inputs[5]), .B(inputs[1]), .Y(keywire227));
NAND_g NAND_g_100_(.A(_026_), .B(_024_), .Y(keywire259));
NAND_g NAND_g_102_(.A(_027_), .B(_025_), .Y(keywire267));
NAND_g NAND_g_103_(.A(inputs[6]), .B(inputs[2]), .Y(keywire233));
NAND_g NAND_g_105_(.A(_030_), .B(_028_), .Y(keywire273));
NAND_g NAND_g_107_(.A(_031_), .B(_029_), .Y(keywire271));
NAND_g NAND_g_108_(.A(inputs[7]), .B(inputs[3]), .Y(keywire241));
NAND_g NAND_g_110_(.A(_034_), .B(_032_), .Y(keywire279));
NAND_g NAND_g_113_(.A(_035_), .B(_033_), .Y(keywire277));
NAND_g NAND_g_128_(.A(_049_), .B(_046_), .Y(keywire310));
NAND_g NAND_g_137_(.A(_058_), .B(_043_), .Y(keywire299));
NAND_g NAND_g_140_(.A(inputs[5]), .B(inputs[1]), .Y(keywire228));
NAND_g NAND_g_142_(.A(_062_), .B(_060_), .Y(keywire262));
NAND_g NAND_g_144_(.A(_063_), .B(_061_), .Y(keywire268));
NAND_g NAND_g_145_(.A(inputs[6]), .B(inputs[2]), .Y(keywire234));
NAND_g NAND_g_147_(.A(_066_), .B(_064_), .Y(keywire275));
NAND_g NAND_g_149_(.A(_067_), .B(_065_), .Y(keywire272));
NAND_g NAND_g_150_(.A(inputs[7]), .B(inputs[3]), .Y(keywire242));
NAND_g NAND_g_152_(.A(_070_), .B(_068_), .Y(keywire281));
NAND_g NAND_g_155_(.A(_071_), .B(_069_), .Y(keywire278));
XOR_g XOR_g_099_(.A(inputs[5]), .B(inputs[1]), .Y(keywire229));
XOR_g XOR_g_101_(.A(_026_), .B(_024_), .Y(keywire260));
XOR_g XOR_g_104_(.A(inputs[6]), .B(inputs[2]), .Y(keywire235));
XOR_g XOR_g_106_(.A(_030_), .B(_028_), .Y(keywire274));
XOR_g XOR_g_109_(.A(inputs[7]), .B(inputs[3]), .Y(keywire243));
XOR_g XOR_g_111_(.A(_034_), .B(_032_), .Y(keywire280));
XOR_g XOR_g_112_(.A(inputs[4]), .B(inputs[0]), .Y(keywire298));
XOR_g XOR_g_141_(.A(inputs[5]), .B(inputs[1]), .Y(keywire230));
XOR_g XOR_g_143_(.A(_062_), .B(_060_), .Y(keywire263));
XOR_g XOR_g_146_(.A(inputs[6]), .B(inputs[2]), .Y(keywire236));
XOR_g XOR_g_148_(.A(_066_), .B(_064_), .Y(keywire276));
XOR_g XOR_g_151_(.A(inputs[7]), .B(inputs[3]), .Y(keywire244));
XOR_g XOR_g_153_(.A(_070_), .B(_068_), .Y(keywire282));
XOR_g XOR_g_154_(.A(inputs[4]), .B(inputs[0]), .Y(keywire300));
XOR_g keygate_XOR_1(.A(keywire75), .B(lockingkeyinput[1]), .Y(_014_));
XOR_g keygate_XOR_3(.A(keywire77), .B(lockingkeyinput[3]), .Y(_023_));
XOR_g keygate_XOR_4(.A(keywire78), .B(lockingkeyinput[4]), .Y(out[0]));
XOR_g keygate_XOR_5(.A(keywire79), .B(lockingkeyinput[5]), .Y(_001_));
XOR_g keygate_XOR_8(.A(keywire82), .B(lockingkeyinput[8]), .Y(_024_));
XOR_g keygate_XOR_10(.A(keywire84), .B(lockingkeyinput[10]), .Y(_060_));
XOR_g keygate_XOR_11(.A(keywire85), .B(lockingkeyinput[11]), .Y(scc[0]));
XOR_g keygate_XOR_12(.A(keywire86), .B(lockingkeyinput[12]), .Y(s1cc[0]));
XOR_g keygate_XOR_13(.A(keywire87), .B(lockingkeyinput[13]), .Y(_004_));
XOR_g keygate_XOR_17(.A(keywire91), .B(lockingkeyinput[17]), .Y(_025_));
XOR_g keygate_XOR_20(.A(keywire94), .B(lockingkeyinput[20]), .Y(_062_));
XOR_g keygate_XOR_23(.A(keywire97), .B(lockingkeyinput[23]), .Y(_029_));
XOR_g keygate_XOR_26(.A(keywire100), .B(lockingkeyinput[26]), .Y(_066_));
XOR_g keygate_XOR_31(.A(keywire105), .B(lockingkeyinput[31]), .Y(_033_));
XOR_g keygate_XOR_32(.A(keywire106), .B(lockingkeyinput[32]), .Y(_069_));
XOR_g keygate_XOR_35(.A(keywire109), .B(lockingkeyinput[35]), .Y(_019_));
XOR_g keygate_XOR_37(.A(keywire111), .B(lockingkeyinput[37]), .Y(_009_));
XOR_g keygate_XOR_38(.A(keywire112), .B(lockingkeyinput[38]), .Y(_045_));
XOR_g keygate_XOR_42(.A(keywire116), .B(lockingkeyinput[42]), .Y(_044_));
XOR_g keygate_XOR_44(.A(keywire118), .B(lockingkeyinput[44]), .Y(_054_));
XOR_g keygate_XOR_46(.A(keywire120), .B(lockingkeyinput[46]), .Y(_038_));
XOR_g keygate_XOR_47(.A(keywire121), .B(lockingkeyinput[47]), .Y(_003_));
XOR_g keygate_XOR_50(.A(keywire124), .B(lockingkeyinput[50]), .Y(scc[1]));
XOR_g keygate_XOR_51(.A(keywire125), .B(lockingkeyinput[51]), .Y(_049_));
XOR_g keygate_XOR_52(.A(keywire126), .B(lockingkeyinput[52]), .Y(_063_));
XOR_g keygate_XOR_53(.A(keywire127), .B(lockingkeyinput[53]), .Y(s1cc[1]));
XOR_g keygate_XOR_54(.A(keywire128), .B(lockingkeyinput[54]), .Y(out[1]));
XOR_g keygate_XOR_55(.A(keywire129), .B(lockingkeyinput[55]), .Y(_006_));
XOR_g keygate_XOR_57(.A(keywire131), .B(lockingkeyinput[57]), .Y(_028_));
XOR_g keygate_XOR_63(.A(keywire137), .B(lockingkeyinput[63]), .Y(_031_));
XOR_g keygate_XOR_67(.A(keywire141), .B(lockingkeyinput[67]), .Y(scc[4]));
XOR_g keygate_XOR_68(.A(keywire142), .B(lockingkeyinput[68]), .Y(s1cc[4]));
XOR_g keygate_XOR_71(.A(keywire145), .B(lockingkeyinput[71]), .Y(_071_));
XOR_g keygate_XOR_75(.A(keywire149), .B(lockingkeyinput[75]), .Y(_010_));
XOR_g keygate_XOR_76(.A(keywire150), .B(lockingkeyinput[76]), .Y(_046_));
XOR_g keygate_XOR_77(.A(keywire151), .B(lockingkeyinput[77]), .Y(_007_));
XOR_g keygate_XOR_78(.A(keywire152), .B(lockingkeyinput[78]), .Y(_043_));
XOR_g keygate_XOR_80(.A(keywire154), .B(lockingkeyinput[80]), .Y(_021_));
XOR_g keygate_XOR_81(.A(keywire155), .B(lockingkeyinput[81]), .Y(_057_));
XOR_g keygate_XOR_84(.A(keywire158), .B(lockingkeyinput[84]), .Y(keywire89));
XOR_g keygate_XOR_85(.A(keywire159), .B(lockingkeyinput[85]), .Y(keywire78));
XOR_g keygate_XOR_89(.A(keywire163), .B(lockingkeyinput[89]), .Y(keywire156));
XOR_g keygate_XOR_92(.A(keywire166), .B(lockingkeyinput[92]), .Y(keywire151));
XOR_g keygate_XOR_93(.A(keywire167), .B(lockingkeyinput[93]), .Y(keywire157));
XOR_g keygate_XOR_94(.A(keywire168), .B(lockingkeyinput[94]), .Y(keywire152));
XOR_g keygate_XOR_100(.A(keywire174), .B(lockingkeyinput[100]), .Y(keywire153));
XOR_g keygate_XOR_101(.A(keywire175), .B(lockingkeyinput[101]), .Y(keywire130));
XOR_g keygate_XOR_105(.A(keywire179), .B(lockingkeyinput[105]), .Y(keywire74));
XOR_g keygate_XOR_107(.A(keywire181), .B(lockingkeyinput[107]), .Y(keywire103));
XOR_g keygate_XOR_110(.A(keywire184), .B(lockingkeyinput[110]), .Y(keywire79));
XOR_g keygate_XOR_111(.A(keywire185), .B(lockingkeyinput[111]), .Y(keywire148));
XOR_g keygate_XOR_112(.A(keywire186), .B(lockingkeyinput[112]), .Y(keywire134));
XOR_g keygate_XOR_114(.A(keywire188), .B(lockingkeyinput[114]), .Y(keywire150));
XOR_g keygate_XOR_117(.A(keywire191), .B(lockingkeyinput[117]), .Y(keywire120));
XOR_g keygate_XOR_118(.A(keywire192), .B(lockingkeyinput[118]), .Y(keywire80));
XOR_g keygate_XOR_120(.A(keywire194), .B(lockingkeyinput[120]), .Y(keywire117));
XOR_g keygate_XOR_122(.A(keywire196), .B(lockingkeyinput[122]), .Y(keywire113));
XOR_g keygate_XOR_123(.A(keywire197), .B(lockingkeyinput[123]), .Y(keywire81));
XOR_g keygate_XOR_125(.A(keywire199), .B(lockingkeyinput[125]), .Y(keywire115));
XOR_g keygate_XOR_126(.A(keywire200), .B(lockingkeyinput[126]), .Y(keywire110));
XOR_g keygate_XOR_127(.A(keywire201), .B(lockingkeyinput[127]), .Y(keywire118));
XOR_g keygate_XOR_130(.A(keywire204), .B(lockingkeyinput[130]), .Y(keywire83));
XOR_g keygate_XOR_132(.A(keywire206), .B(lockingkeyinput[132]), .Y(keywire112));
XOR_g keygate_XOR_134(.A(keywire208), .B(lockingkeyinput[134]), .Y(keywire101));
XOR_g keygate_XOR_135(.A(keywire209), .B(lockingkeyinput[135]), .Y(keywire102));
XOR_g keygate_XOR_138(.A(keywire212), .B(lockingkeyinput[138]), .Y(keywire165));
XOR_g keygate_XOR_140(.A(keywire214), .B(lockingkeyinput[140]), .Y(keywire159));
XOR_g keygate_XOR_144(.A(keywire218), .B(lockingkeyinput[144]), .Y(keywire82));
XOR_g keygate_XOR_146(.A(keywire220), .B(lockingkeyinput[146]), .Y(keywire84));
XOR_g keygate_XOR_154(.A(keywire228), .B(lockingkeyinput[154]), .Y(keywire92));
XOR_g keygate_XOR_156(.A(keywire230), .B(lockingkeyinput[156]), .Y(keywire94));
XOR_g keygate_XOR_159(.A(keywire233), .B(lockingkeyinput[159]), .Y(keywire97));
XOR_g keygate_XOR_161(.A(keywire235), .B(lockingkeyinput[161]), .Y(keywire99));
XOR_g keygate_XOR_163(.A(keywire237), .B(lockingkeyinput[163]), .Y(keywire208));
XOR_g keygate_XOR_166(.A(keywire240), .B(lockingkeyinput[166]), .Y(keywire189));
XOR_g keygate_XOR_167(.A(keywire241), .B(lockingkeyinput[167]), .Y(keywire105));
XOR_g keygate_XOR_168(.A(keywire242), .B(lockingkeyinput[168]), .Y(keywire106));
XOR_g keygate_XOR_171(.A(keywire245), .B(lockingkeyinput[171]), .Y(keywire193));
XOR_g keygate_XOR_172(.A(keywire246), .B(lockingkeyinput[172]), .Y(keywire200));
XOR_g keygate_XOR_173(.A(keywire247), .B(lockingkeyinput[173]), .Y(keywire198));
XOR_g keygate_XOR_182(.A(keywire256), .B(lockingkeyinput[182]), .Y(keywire191));
XOR_g keygate_XOR_185(.A(keywire259), .B(lockingkeyinput[185]), .Y(keywire123));
XOR_g keygate_XOR_188(.A(keywire262), .B(lockingkeyinput[188]), .Y(keywire126));
XOR_g keygate_XOR_189(.A(keywire263), .B(lockingkeyinput[189]), .Y(keywire127));
XOR_g keygate_XOR_191(.A(keywire265), .B(lockingkeyinput[191]), .Y(keywire171));
XOR_g keygate_XOR_192(.A(keywire266), .B(lockingkeyinput[192]), .Y(keywire175));
XOR_g keygate_XOR_193(.A(keywire267), .B(lockingkeyinput[193]), .Y(keywire131));
XOR_g keygate_XOR_194(.A(keywire268), .B(lockingkeyinput[194]), .Y(keywire132));
XOR_g keygate_XOR_196(.A(keywire270), .B(lockingkeyinput[196]), .Y(keywire186));
XOR_g keygate_XOR_197(.A(keywire271), .B(lockingkeyinput[197]), .Y(keywire135));
XOR_g keygate_XOR_198(.A(keywire272), .B(lockingkeyinput[198]), .Y(keywire136));
XOR_g keygate_XOR_203(.A(keywire277), .B(lockingkeyinput[203]), .Y(keywire141));
XOR_g keygate_XOR_205(.A(keywire279), .B(lockingkeyinput[205]), .Y(keywire143));
XOR_g keygate_XOR_206(.A(keywire280), .B(lockingkeyinput[206]), .Y(keywire144));
XOR_g keygate_XOR_210(.A(keywire284), .B(lockingkeyinput[210]), .Y(keywire185));
XOR_g keygate_XOR_212(.A(keywire286), .B(lockingkeyinput[212]), .Y(keywire188));
XOR_g keygate_XOR_213(.A(keywire287), .B(lockingkeyinput[213]), .Y(keywire166));
XOR_g keygate_XOR_214(.A(keywire288), .B(lockingkeyinput[214]), .Y(keywire168));
XOR_g keygate_XOR_216(.A(keywire290), .B(lockingkeyinput[216]), .Y(keywire169));
XOR_g keygate_XOR_220(.A(keywire294), .B(lockingkeyinput[220]), .Y(keywire225));
XOR_g keygate_XOR_221(.A(keywire295), .B(lockingkeyinput[221]), .Y(keywire214));
XOR_g keygate_XOR_222(.A(keywire296), .B(lockingkeyinput[222]), .Y(keywire264));
XOR_g keygate_XOR_225(.A(keywire299), .B(lockingkeyinput[225]), .Y(keywire292));
XOR_g keygate_XOR_228(.A(keywire302), .B(lockingkeyinput[228]), .Y(keywire287));
XOR_g keygate_XOR_230(.A(keywire304), .B(lockingkeyinput[230]), .Y(keywire288));
XOR_g keygate_XOR_234(.A(keywire308), .B(lockingkeyinput[234]), .Y(keywire257));
XOR_g keygate_XOR_235(.A(keywire309), .B(lockingkeyinput[235]), .Y(keywire291));
XOR_g keygate_XOR_237(.A(keywire311), .B(lockingkeyinput[237]), .Y(keywire266));
XOR_g keygate_XOR_238(.A(keywire312), .B(lockingkeyinput[238]), .Y(keywire258));
XOR_g keygate_XOR_239(.A(keywire313), .B(lockingkeyinput[239]), .Y(keywire283));
XOR_g keygate_XOR_240(.A(keywire314), .B(lockingkeyinput[240]), .Y(keywire269));
XOR_g keygate_XOR_241(.A(keywire315), .B(lockingkeyinput[241]), .Y(keywire210));
XOR_g keygate_XOR_242(.A(keywire316), .B(lockingkeyinput[242]), .Y(keywire285));
XOR_g keygate_XOR_243(.A(keywire317), .B(lockingkeyinput[243]), .Y(keywire239));
XOR_g keygate_XOR_249(.A(keywire323), .B(lockingkeyinput[249]), .Y(keywire261));
XOR_g keygate_XOR_250(.A(keywire324), .B(lockingkeyinput[250]), .Y(keywire286));
XOR_g keygate_XOR_251(.A(keywire325), .B(lockingkeyinput[251]), .Y(keywire240));
XOR_g keygate_XOR_253(.A(keywire327), .B(lockingkeyinput[253]), .Y(keywire256));
XOR_g keygate_XOR_255(.A(keywire329), .B(lockingkeyinput[255]), .Y(keywire245));
endmodule

module BUF_g(A, Y);
input A;
output Y;
assign Y=A;
endmodule

 
module NOT_g(A, Y);
input A;
output Y;
assign Y=~A;
endmodule

module AND_g(A, B, Y);
input A, B;
output Y;
assign Y=(A & B);
endmodule

module OR_g(A, B, Y);
input A, B;
output Y;
assign Y= (A | B);
endmodule

module NAND_g(A, B, Y);
input A, B;
output Y;
assign Y= ~(A & B);

endmodule

module NOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A | B);
endmodule


module XOR_g(A, B, Y);
input A, B;
output Y;
assign Y = (A ^ B);
endmodule

module XNOR_g(A, B, Y);
input A, B;
output Y;
assign Y = ~(A ^ B);
endmodule

module DFFcell(C, D, Q);
input C, D;
output reg Q;
always @(posedge C)
	Q <= D;
endmodule


module DFFRcell(C, D, Q, R);
input C, D, R;
output reg Q;
always @(posedge C, negedge R)
	if (!R)
		Q <= 1'b0;
	else
		Q <= D;
endmodule
