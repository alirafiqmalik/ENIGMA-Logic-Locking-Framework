module c3540(N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire _0828_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0833_;
wire _0834_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
input N1;
wire N1;
input N107;
wire N107;
input N116;
wire N116;
input N124;
wire N124;
input N125;
wire N125;
input N128;
wire N128;
input N13;
wire N13;
input N132;
wire N132;
input N137;
wire N137;
input N143;
wire N143;
input N150;
wire N150;
input N159;
wire N159;
input N169;
wire N169;
output N1713;
wire N1713;
input N179;
wire N179;
input N190;
wire N190;
output N1947;
wire N1947;
input N20;
wire N20;
input N200;
wire N200;
input N213;
wire N213;
input N222;
wire N222;
input N223;
wire N223;
input N226;
wire N226;
input N232;
wire N232;
input N238;
wire N238;
input N244;
wire N244;
input N250;
wire N250;
input N257;
wire N257;
input N264;
wire N264;
input N270;
wire N270;
input N274;
wire N274;
input N283;
wire N283;
input N294;
wire N294;
input N303;
wire N303;
input N311;
wire N311;
input N317;
wire N317;
output N3195;
wire N3195;
input N322;
wire N322;
input N326;
wire N326;
input N329;
wire N329;
input N33;
wire N33;
input N330;
wire N330;
input N343;
wire N343;
input N349;
wire N349;
input N350;
wire N350;
output N3833;
wire N3833;
output N3987;
wire N3987;
output N4028;
wire N4028;
input N41;
wire N41;
output N4145;
wire N4145;
input N45;
wire N45;
output N4589;
wire N4589;
output N4667;
wire N4667;
output N4815;
wire N4815;
output N4944;
wire N4944;
input N50;
wire N50;
output N5002;
wire N5002;
output N5045;
wire N5045;
output N5047;
wire N5047;
output N5078;
wire N5078;
output N5102;
wire N5102;
output N5120;
wire N5120;
output N5121;
wire N5121;
output N5192;
wire N5192;
output N5231;
wire N5231;
output N5360;
wire N5360;
output N5361;
wire N5361;
input N58;
wire N58;
input N68;
wire N68;
input N77;
wire N77;
input N87;
wire N87;
input N97;
wire N97;
NOT_g _0873_ ( .A(N116), .Y(_0633_));
NOT_g _0874_ ( .A(N13), .Y(_0644_));
NOT_g _0875_ ( .A(N41), .Y(_0654_));
NOT_g _0876_ ( .A(N45), .Y(_0665_));
NOT_g _0877_ ( .A(N200), .Y(_0676_));
NOT_g _0878_ ( .A(N20), .Y(_0687_));
NOT_g _0879_ ( .A(N330), .Y(_0698_));
NOT_g _0880_ ( .A(N68), .Y(_0709_));
NOT_g _0881_ ( .A(N1), .Y(_0719_));
NOT_g _0882_ ( .A(N33), .Y(_0730_));
NOT_g _0883_ ( .A(N169), .Y(_0741_));
NOT_g _0884_ ( .A(N190), .Y(_0752_));
NOT_g _0885_ ( .A(N343), .Y(_0763_));
NOT_g _0886_ ( .A(N274), .Y(_0774_));
AND_g _0887_ ( .A(N20), .B(N1), .Y(_0784_));
NAND_g _0888_ ( .A(N87), .B(N250), .Y(_0795_));
NAND_g _0889_ ( .A(N232), .B(N58), .Y(_0806_));
AND_g _0890_ ( .A(_0795_), .B(_0806_), .Y(_0817_));
NAND_g _0891_ ( .A(N116), .B(N270), .Y(_0827_));
NAND_g _0892_ ( .A(N97), .B(N257), .Y(_0837_));
AND_g _0893_ ( .A(_0827_), .B(_0837_), .Y(_0846_));
AND_g _0894_ ( .A(_0817_), .B(_0846_), .Y(_0852_));
NAND_g _0895_ ( .A(N226), .B(N50), .Y(_0862_));
NAND_g _0896_ ( .A(N238), .B(N68), .Y(_0869_));
AND_g _0897_ ( .A(_0862_), .B(_0869_), .Y(_0870_));
NAND_g _0898_ ( .A(N264), .B(N107), .Y(_0871_));
NAND_g _0899_ ( .A(N77), .B(N244), .Y(_0872_));
AND_g _0900_ ( .A(_0871_), .B(_0872_), .Y(_0000_));
AND_g _0901_ ( .A(_0870_), .B(_0000_), .Y(_0001_));
AND_g _0902_ ( .A(_0852_), .B(_0001_), .Y(_0002_));
NOR_g _0903_ ( .A(_0784_), .B(_0002_), .Y(_0003_));
AND_g _0904_ ( .A(N13), .B(N1), .Y(_0004_));
AND_g _0905_ ( .A(N13), .B(_0784_), .Y(_0005_));
NOR_g _0906_ ( .A(N58), .B(N68), .Y(_0006_));
NOT_g _0907_ ( .A(_0006_), .Y(_0007_));
AND_g _0908_ ( .A(N50), .B(_0007_), .Y(_0008_));
NAND_g _0909_ ( .A(_0005_), .B(_0008_), .Y(_0009_));
AND_g _0910_ ( .A(_0644_), .B(N1), .Y(_0010_));
AND_g _0911_ ( .A(_0644_), .B(_0784_), .Y(_0011_));
NAND_g _0912_ ( .A(_0644_), .B(_0784_), .Y(_0012_));
NOR_g _0913_ ( .A(N257), .B(N264), .Y(_0013_));
NOR_g _0914_ ( .A(_0012_), .B(_0013_), .Y(_0014_));
NAND_g _0915_ ( .A(N250), .B(_0014_), .Y(_0015_));
NAND_g _0916_ ( .A(_0009_), .B(_0015_), .Y(_0016_));
NOR_g _0917_ ( .A(_0003_), .B(_0016_), .Y(N3195));
NOR_g _0918_ ( .A(N58), .B(N50), .Y(_0017_));
NAND_g _0919_ ( .A(N58), .B(N50), .Y(_0018_));
XOR_g _0920_ ( .A(N58), .B(N50), .Y(_0019_));
NAND_g _0921_ ( .A(N77), .B(N68), .Y(_0020_));
NOR_g _0922_ ( .A(N77), .B(N68), .Y(_0021_));
XOR_g _0923_ ( .A(N77), .B(N68), .Y(_0022_));
XNOR_g _0924_ ( .A(_0019_), .B(_0022_), .Y(_0023_));
NOR_g _0925_ ( .A(N97), .B(N107), .Y(_0024_));
NOT_g _0926_ ( .A(_0024_), .Y(_0025_));
XOR_g _0927_ ( .A(N97), .B(N107), .Y(_0026_));
XNOR_g _0928_ ( .A(N97), .B(N107), .Y(_0027_));
XOR_g _0929_ ( .A(N116), .B(N87), .Y(_0028_));
XNOR_g _0930_ ( .A(_0026_), .B(_0028_), .Y(_0029_));
XNOR_g _0931_ ( .A(_0023_), .B(_0029_), .Y(N3987));
NOR_g _0932_ ( .A(N13), .B(N33), .Y(_0030_));
NAND_g _0933_ ( .A(_0644_), .B(_0730_), .Y(_0031_));
AND_g _0934_ ( .A(N13), .B(_0687_), .Y(_0032_));
AND_g _0935_ ( .A(N213), .B(_0719_), .Y(_0033_));
AND_g _0936_ ( .A(_0032_), .B(_0033_), .Y(_0034_));
AND_g _0937_ ( .A(N343), .B(_0034_), .Y(_0035_));
NAND_g _0938_ ( .A(N343), .B(_0034_), .Y(_0036_));
AND_g _0939_ ( .A(N33), .B(_0011_), .Y(_0037_));
NOR_g _0940_ ( .A(_0004_), .B(_0037_), .Y(_0038_));
AND_g _0941_ ( .A(N20), .B(_0719_), .Y(_0039_));
NAND_g _0942_ ( .A(N20), .B(_0719_), .Y(_0040_));
NAND_g _0943_ ( .A(_0038_), .B(_0040_), .Y(_0041_));
NOT_g _0944_ ( .A(_0041_), .Y(_0042_));
NAND_g _0945_ ( .A(_0784_), .B(_0031_), .Y(_0043_));
NOT_g _0946_ ( .A(_0043_), .Y(_0044_));
NAND_g _0947_ ( .A(_0041_), .B(_0043_), .Y(_0045_));
AND_g _0948_ ( .A(N77), .B(_0045_), .Y(_0046_));
NAND_g _0949_ ( .A(N87), .B(N33), .Y(_0047_));
NAND_g _0950_ ( .A(N58), .B(_0730_), .Y(_0048_));
NAND_g _0951_ ( .A(_0047_), .B(_0048_), .Y(_0049_));
AND_g _0952_ ( .A(_0687_), .B(_0004_), .Y(_0050_));
NAND_g _0953_ ( .A(_0049_), .B(_0050_), .Y(_0051_));
NAND_g _0954_ ( .A(N13), .B(_0039_), .Y(_0052_));
NOR_g _0955_ ( .A(N77), .B(_0052_), .Y(_0053_));
NOR_g _0956_ ( .A(_0046_), .B(_0053_), .Y(_0054_));
NAND_g _0957_ ( .A(_0051_), .B(_0054_), .Y(_0055_));
AND_g _0958_ ( .A(_0035_), .B(_0055_), .Y(_0056_));
NAND_g _0959_ ( .A(N41), .B(N33), .Y(_0057_));
AND_g _0960_ ( .A(_0004_), .B(_0057_), .Y(_0058_));
NAND_g _0961_ ( .A(_0004_), .B(_0057_), .Y(_0059_));
NOR_g _0962_ ( .A(N33), .B(N349), .Y(_0060_));
AND_g _0963_ ( .A(_0730_), .B(N349), .Y(_0061_));
NAND_g _0964_ ( .A(N238), .B(_0061_), .Y(_0062_));
NAND_g _0965_ ( .A(N232), .B(_0060_), .Y(_0063_));
NAND_g _0966_ ( .A(N107), .B(N33), .Y(_0064_));
AND_g _0967_ ( .A(_0063_), .B(_0064_), .Y(_0065_));
NAND_g _0968_ ( .A(_0062_), .B(_0065_), .Y(_0066_));
NAND_g _0969_ ( .A(_0058_), .B(_0066_), .Y(_0067_));
NOR_g _0970_ ( .A(N41), .B(N45), .Y(_0068_));
AND_g _0971_ ( .A(N45), .B(_0719_), .Y(_0069_));
NOR_g _0972_ ( .A(N1), .B(_0068_), .Y(_0070_));
NOR_g _0973_ ( .A(_0058_), .B(_0070_), .Y(_0071_));
NAND_g _0974_ ( .A(N244), .B(_0071_), .Y(_0072_));
AND_g _0975_ ( .A(N274), .B(_0059_), .Y(_0073_));
NAND_g _0976_ ( .A(_0070_), .B(_0073_), .Y(_0074_));
AND_g _0977_ ( .A(_0067_), .B(_0072_), .Y(_0075_));
AND_g _0978_ ( .A(_0074_), .B(_0075_), .Y(_0076_));
NAND_g _0979_ ( .A(_0074_), .B(_0075_), .Y(_0077_));
NAND_g _0980_ ( .A(N169), .B(_0077_), .Y(_0078_));
NAND_g _0981_ ( .A(N179), .B(_0076_), .Y(_0079_));
NAND_g _0982_ ( .A(_0078_), .B(_0079_), .Y(_0080_));
AND_g _0983_ ( .A(_0055_), .B(_0080_), .Y(_0081_));
NAND_g _0984_ ( .A(N190), .B(_0076_), .Y(_0082_));
NAND_g _0985_ ( .A(N200), .B(_0077_), .Y(_0083_));
NAND_g _0986_ ( .A(_0082_), .B(_0083_), .Y(_0084_));
NOR_g _0987_ ( .A(_0055_), .B(_0084_), .Y(_0085_));
NOR_g _0988_ ( .A(_0081_), .B(_0085_), .Y(_0086_));
XNOR_g _0989_ ( .A(_0056_), .B(_0086_), .Y(_0087_));
NOT_g _0990_ ( .A(_0087_), .Y(_0088_));
NAND_g _0991_ ( .A(_0030_), .B(_0087_), .Y(_0089_));
NAND_g _0992_ ( .A(N20), .B(_0741_), .Y(_0090_));
AND_g _0993_ ( .A(_0004_), .B(_0090_), .Y(_0091_));
NOT_g _0994_ ( .A(_0091_), .Y(_0092_));
AND_g _0995_ ( .A(N20), .B(N179), .Y(_0093_));
NAND_g _0996_ ( .A(N20), .B(N179), .Y(_0094_));
NAND_g _0997_ ( .A(_0676_), .B(_0093_), .Y(_0095_));
NOR_g _0998_ ( .A(N190), .B(_0095_), .Y(_0096_));
NAND_g _0999_ ( .A(N159), .B(_0096_), .Y(_0097_));
AND_g _1000_ ( .A(N20), .B(_0752_), .Y(_0098_));
NAND_g _1001_ ( .A(N20), .B(_0752_), .Y(_0099_));
NAND_g _1002_ ( .A(N200), .B(N20), .Y(_0100_));
AND_g _1003_ ( .A(_0094_), .B(_0100_), .Y(_0101_));
AND_g _1004_ ( .A(_0099_), .B(_0101_), .Y(_0102_));
NAND_g _1005_ ( .A(N58), .B(_0102_), .Y(_0103_));
AND_g _1006_ ( .A(N200), .B(_0093_), .Y(_0104_));
AND_g _1007_ ( .A(N190), .B(_0104_), .Y(_0105_));
NAND_g _1008_ ( .A(N137), .B(_0105_), .Y(_0106_));
AND_g _1009_ ( .A(_0752_), .B(_0104_), .Y(_0107_));
NAND_g _1010_ ( .A(N150), .B(_0107_), .Y(_0108_));
NOR_g _1011_ ( .A(N179), .B(_0100_), .Y(_0109_));
AND_g _1012_ ( .A(N190), .B(_0109_), .Y(_0110_));
NAND_g _1013_ ( .A(N50), .B(_0110_), .Y(_0111_));
AND_g _1014_ ( .A(_0752_), .B(_0109_), .Y(_0112_));
NAND_g _1015_ ( .A(N68), .B(_0112_), .Y(_0113_));
NOR_g _1016_ ( .A(_0752_), .B(_0095_), .Y(_0114_));
NAND_g _1017_ ( .A(N143), .B(_0114_), .Y(_0115_));
AND_g _1018_ ( .A(_0098_), .B(_0101_), .Y(_0116_));
NAND_g _1019_ ( .A(N132), .B(_0116_), .Y(_0117_));
AND_g _1020_ ( .A(_0103_), .B(_0111_), .Y(_0118_));
AND_g _1021_ ( .A(_0113_), .B(_0118_), .Y(_0119_));
AND_g _1022_ ( .A(_0097_), .B(_0108_), .Y(_0120_));
AND_g _1023_ ( .A(_0117_), .B(_0120_), .Y(_0121_));
AND_g _1024_ ( .A(_0730_), .B(_0115_), .Y(_0122_));
AND_g _1025_ ( .A(_0106_), .B(_0122_), .Y(_0123_));
AND_g _1026_ ( .A(_0121_), .B(_0123_), .Y(_0124_));
NAND_g _1027_ ( .A(_0119_), .B(_0124_), .Y(_0125_));
NAND_g _1028_ ( .A(N303), .B(_0105_), .Y(_0126_));
NAND_g _1029_ ( .A(N116), .B(_0096_), .Y(_0127_));
NAND_g _1030_ ( .A(N107), .B(_0110_), .Y(_0128_));
AND_g _1031_ ( .A(_0127_), .B(_0128_), .Y(_0129_));
AND_g _1032_ ( .A(_0126_), .B(_0129_), .Y(_0130_));
NAND_g _1033_ ( .A(N294), .B(_0114_), .Y(_0131_));
AND_g _1034_ ( .A(N33), .B(_0131_), .Y(_0132_));
NAND_g _1035_ ( .A(N311), .B(_0116_), .Y(_0133_));
NAND_g _1036_ ( .A(N87), .B(_0112_), .Y(_0134_));
AND_g _1037_ ( .A(_0133_), .B(_0134_), .Y(_0135_));
NAND_g _1038_ ( .A(N283), .B(_0107_), .Y(_0136_));
NAND_g _1039_ ( .A(N97), .B(_0102_), .Y(_0137_));
AND_g _1040_ ( .A(_0136_), .B(_0137_), .Y(_0138_));
AND_g _1041_ ( .A(_0135_), .B(_0138_), .Y(_0139_));
AND_g _1042_ ( .A(_0132_), .B(_0139_), .Y(_0140_));
NAND_g _1043_ ( .A(_0130_), .B(_0140_), .Y(_0141_));
NAND_g _1044_ ( .A(_0125_), .B(_0141_), .Y(_0142_));
NAND_g _1045_ ( .A(_0091_), .B(_0142_), .Y(_0143_));
AND_g _1046_ ( .A(_0654_), .B(_0011_), .Y(_0144_));
NAND_g _1047_ ( .A(N45), .B(_0032_), .Y(_0145_));
AND_g _1048_ ( .A(N1), .B(_0145_), .Y(_0146_));
NAND_g _1049_ ( .A(N1), .B(_0145_), .Y(_0147_));
NOR_g _1050_ ( .A(_0719_), .B(_0144_), .Y(_0148_));
NOR_g _1051_ ( .A(_0144_), .B(_0147_), .Y(_0149_));
NOT_g _1052_ ( .A(_0149_), .Y(_0150_));
NAND_g _1053_ ( .A(_0031_), .B(_0092_), .Y(_0151_));
NOR_g _1054_ ( .A(N77), .B(_0151_), .Y(_0152_));
NOR_g _1055_ ( .A(_0150_), .B(_0152_), .Y(_0153_));
AND_g _1056_ ( .A(_0143_), .B(_0153_), .Y(_0154_));
NAND_g _1057_ ( .A(_0089_), .B(_0154_), .Y(_0155_));
NAND_g _1058_ ( .A(N250), .B(_0061_), .Y(_0156_));
NAND_g _1059_ ( .A(N33), .B(N283), .Y(_0157_));
NAND_g _1060_ ( .A(N244), .B(_0060_), .Y(_0158_));
AND_g _1061_ ( .A(_0157_), .B(_0158_), .Y(_0159_));
NAND_g _1062_ ( .A(_0156_), .B(_0159_), .Y(_0160_));
NAND_g _1063_ ( .A(_0058_), .B(_0160_), .Y(_0161_));
AND_g _1064_ ( .A(_0654_), .B(_0069_), .Y(_0162_));
NAND_g _1065_ ( .A(_0654_), .B(_0069_), .Y(_0163_));
AND_g _1066_ ( .A(N257), .B(_0059_), .Y(_0164_));
NAND_g _1067_ ( .A(_0163_), .B(_0164_), .Y(_0165_));
NAND_g _1068_ ( .A(_0073_), .B(_0162_), .Y(_0166_));
AND_g _1069_ ( .A(_0165_), .B(_0166_), .Y(_0167_));
NAND_g _1070_ ( .A(_0161_), .B(_0167_), .Y(_0168_));
NOT_g _1071_ ( .A(_0168_), .Y(_0169_));
NAND_g _1072_ ( .A(N244), .B(_0061_), .Y(_0170_));
NAND_g _1073_ ( .A(N238), .B(_0060_), .Y(_0171_));
NAND_g _1074_ ( .A(N116), .B(N33), .Y(_0172_));
AND_g _1075_ ( .A(_0171_), .B(_0172_), .Y(_0173_));
NAND_g _1076_ ( .A(_0170_), .B(_0173_), .Y(_0174_));
NAND_g _1077_ ( .A(_0058_), .B(_0174_), .Y(_0175_));
NAND_g _1078_ ( .A(_0774_), .B(_0069_), .Y(_0176_));
NOR_g _1079_ ( .A(N250), .B(_0069_), .Y(_0177_));
NOR_g _1080_ ( .A(_0058_), .B(_0177_), .Y(_0178_));
NAND_g _1081_ ( .A(_0176_), .B(_0178_), .Y(_0179_));
AND_g _1082_ ( .A(_0175_), .B(_0179_), .Y(_0180_));
NAND_g _1083_ ( .A(_0175_), .B(_0179_), .Y(_0181_));
NAND_g _1084_ ( .A(N264), .B(_0061_), .Y(_0182_));
NAND_g _1085_ ( .A(N33), .B(N303), .Y(_0183_));
NAND_g _1086_ ( .A(N257), .B(_0060_), .Y(_0184_));
AND_g _1087_ ( .A(_0183_), .B(_0184_), .Y(_0185_));
NAND_g _1088_ ( .A(_0182_), .B(_0185_), .Y(_0186_));
NAND_g _1089_ ( .A(_0058_), .B(_0186_), .Y(_0187_));
AND_g _1090_ ( .A(N270), .B(_0059_), .Y(_0188_));
NAND_g _1091_ ( .A(_0163_), .B(_0188_), .Y(_0189_));
AND_g _1092_ ( .A(_0166_), .B(_0189_), .Y(_0190_));
AND_g _1093_ ( .A(_0187_), .B(_0190_), .Y(_0191_));
NOT_g _1094_ ( .A(_0191_), .Y(_0192_));
NAND_g _1095_ ( .A(N257), .B(_0061_), .Y(_0193_));
NAND_g _1096_ ( .A(N250), .B(_0060_), .Y(_0194_));
NAND_g _1097_ ( .A(N33), .B(N294), .Y(_0195_));
AND_g _1098_ ( .A(_0194_), .B(_0195_), .Y(_0196_));
NAND_g _1099_ ( .A(_0193_), .B(_0196_), .Y(_0197_));
NAND_g _1100_ ( .A(_0058_), .B(_0197_), .Y(_0198_));
AND_g _1101_ ( .A(N264), .B(_0059_), .Y(_0199_));
NAND_g _1102_ ( .A(_0163_), .B(_0199_), .Y(_0200_));
AND_g _1103_ ( .A(_0166_), .B(_0198_), .Y(_0201_));
AND_g _1104_ ( .A(_0200_), .B(_0201_), .Y(_0202_));
NAND_g _1105_ ( .A(_0200_), .B(_0201_), .Y(_0203_));
NAND_g _1106_ ( .A(N179), .B(_0180_), .Y(_0204_));
NOR_g _1107_ ( .A(N179), .B(_0180_), .Y(_0205_));
AND_g _1108_ ( .A(_0203_), .B(_0205_), .Y(_0206_));
NAND_g _1109_ ( .A(_0168_), .B(_0206_), .Y(_0207_));
NOR_g _1110_ ( .A(_0203_), .B(_0204_), .Y(_0208_));
NAND_g _1111_ ( .A(_0191_), .B(_0208_), .Y(_0209_));
NAND_g _1112_ ( .A(_0207_), .B(_0209_), .Y(_0210_));
NAND_g _1113_ ( .A(_0168_), .B(_0191_), .Y(_0211_));
AND_g _1114_ ( .A(_0035_), .B(_0211_), .Y(_0212_));
NAND_g _1115_ ( .A(_0210_), .B(_0212_), .Y(_0213_));
AND_g _1116_ ( .A(_0687_), .B(N33), .Y(_0214_));
NOR_g _1117_ ( .A(N20), .B(N33), .Y(_0215_));
NAND_g _1118_ ( .A(N68), .B(_0215_), .Y(_0216_));
NOR_g _1119_ ( .A(N87), .B(_0025_), .Y(_0217_));
AND_g _1120_ ( .A(N97), .B(N33), .Y(_0218_));
NOR_g _1121_ ( .A(_0687_), .B(_0217_), .Y(_0219_));
NAND_g _1122_ ( .A(_0687_), .B(_0218_), .Y(_0220_));
NAND_g _1123_ ( .A(_0216_), .B(_0220_), .Y(_0221_));
NOR_g _1124_ ( .A(_0219_), .B(_0221_), .Y(_0222_));
NOR_g _1125_ ( .A(_0038_), .B(_0222_), .Y(_0223_));
NAND_g _1126_ ( .A(_0719_), .B(N33), .Y(_0224_));
AND_g _1127_ ( .A(_0052_), .B(_0224_), .Y(_0225_));
AND_g _1128_ ( .A(_0038_), .B(_0225_), .Y(_0226_));
NAND_g _1129_ ( .A(N87), .B(_0226_), .Y(_0227_));
NOR_g _1130_ ( .A(N87), .B(_0052_), .Y(_0228_));
NOR_g _1131_ ( .A(_0223_), .B(_0228_), .Y(_0229_));
AND_g _1132_ ( .A(_0227_), .B(_0229_), .Y(_0230_));
NAND_g _1133_ ( .A(_0227_), .B(_0229_), .Y(_0231_));
NAND_g _1134_ ( .A(N169), .B(_0181_), .Y(_0232_));
NAND_g _1135_ ( .A(_0204_), .B(_0232_), .Y(_0233_));
NAND_g _1136_ ( .A(_0231_), .B(_0233_), .Y(_0234_));
NAND_g _1137_ ( .A(_0676_), .B(_0181_), .Y(_0235_));
NAND_g _1138_ ( .A(_0752_), .B(_0180_), .Y(_0236_));
NAND_g _1139_ ( .A(_0235_), .B(_0236_), .Y(_0237_));
NAND_g _1140_ ( .A(_0230_), .B(_0237_), .Y(_0238_));
AND_g _1141_ ( .A(_0234_), .B(_0238_), .Y(_0239_));
NAND_g _1142_ ( .A(N97), .B(_0226_), .Y(_0240_));
NAND_g _1143_ ( .A(N20), .B(_0027_), .Y(_0241_));
NAND_g _1144_ ( .A(N107), .B(_0214_), .Y(_0242_));
NAND_g _1145_ ( .A(N77), .B(_0215_), .Y(_0243_));
AND_g _1146_ ( .A(_0241_), .B(_0243_), .Y(_0244_));
AND_g _1147_ ( .A(_0242_), .B(_0244_), .Y(_0245_));
NOR_g _1148_ ( .A(_0038_), .B(_0245_), .Y(_0246_));
NOR_g _1149_ ( .A(N97), .B(_0052_), .Y(_0247_));
NOR_g _1150_ ( .A(_0246_), .B(_0247_), .Y(_0248_));
NAND_g _1151_ ( .A(_0240_), .B(_0248_), .Y(_0249_));
AND_g _1152_ ( .A(_0741_), .B(_0168_), .Y(_0250_));
NOR_g _1153_ ( .A(N179), .B(_0168_), .Y(_0251_));
NOR_g _1154_ ( .A(_0250_), .B(_0251_), .Y(_0252_));
NAND_g _1155_ ( .A(_0249_), .B(_0252_), .Y(_0253_));
NAND_g _1156_ ( .A(N190), .B(_0169_), .Y(_0254_));
AND_g _1157_ ( .A(N200), .B(_0168_), .Y(_0255_));
NOR_g _1158_ ( .A(_0249_), .B(_0255_), .Y(_0256_));
NAND_g _1159_ ( .A(_0254_), .B(_0256_), .Y(_0257_));
AND_g _1160_ ( .A(_0253_), .B(_0257_), .Y(_0258_));
AND_g _1161_ ( .A(_0239_), .B(_0258_), .Y(_0259_));
NAND_g _1162_ ( .A(N107), .B(_0226_), .Y(_0260_));
NAND_g _1163_ ( .A(N87), .B(_0730_), .Y(_0261_));
NAND_g _1164_ ( .A(_0172_), .B(_0261_), .Y(_0262_));
AND_g _1165_ ( .A(_0050_), .B(_0262_), .Y(_0263_));
AND_g _1166_ ( .A(_0043_), .B(_0052_), .Y(_0264_));
NOR_g _1167_ ( .A(N107), .B(_0264_), .Y(_0265_));
NOR_g _1168_ ( .A(_0263_), .B(_0265_), .Y(_0266_));
NAND_g _1169_ ( .A(_0260_), .B(_0266_), .Y(_0267_));
AND_g _1170_ ( .A(_0741_), .B(_0203_), .Y(_0268_));
NOR_g _1171_ ( .A(N179), .B(_0203_), .Y(_0269_));
NOR_g _1172_ ( .A(_0268_), .B(_0269_), .Y(_0270_));
AND_g _1173_ ( .A(_0267_), .B(_0270_), .Y(_0271_));
NAND_g _1174_ ( .A(_0267_), .B(_0270_), .Y(_0272_));
NAND_g _1175_ ( .A(N190), .B(_0202_), .Y(_0273_));
AND_g _1176_ ( .A(N200), .B(_0203_), .Y(_0274_));
NOR_g _1177_ ( .A(_0267_), .B(_0274_), .Y(_0275_));
NAND_g _1178_ ( .A(_0273_), .B(_0275_), .Y(_0276_));
AND_g _1179_ ( .A(_0272_), .B(_0276_), .Y(_0277_));
AND_g _1180_ ( .A(_0259_), .B(_0277_), .Y(_0278_));
NOR_g _1181_ ( .A(_0044_), .B(_0226_), .Y(_0279_));
NOR_g _1182_ ( .A(_0633_), .B(_0279_), .Y(_0280_));
NAND_g _1183_ ( .A(N97), .B(_0730_), .Y(_0281_));
NAND_g _1184_ ( .A(_0157_), .B(_0281_), .Y(_0282_));
NAND_g _1185_ ( .A(_0050_), .B(_0282_), .Y(_0283_));
NOR_g _1186_ ( .A(N116), .B(_0052_), .Y(_0284_));
NOR_g _1187_ ( .A(_0280_), .B(_0284_), .Y(_0285_));
NAND_g _1188_ ( .A(_0283_), .B(_0285_), .Y(_0286_));
NAND_g _1189_ ( .A(N169), .B(_0192_), .Y(_0287_));
NAND_g _1190_ ( .A(N179), .B(_0191_), .Y(_0288_));
NAND_g _1191_ ( .A(_0287_), .B(_0288_), .Y(_0289_));
AND_g _1192_ ( .A(_0286_), .B(_0289_), .Y(_0290_));
NAND_g _1193_ ( .A(N190), .B(_0191_), .Y(_0291_));
NAND_g _1194_ ( .A(N200), .B(_0192_), .Y(_0292_));
NAND_g _1195_ ( .A(_0291_), .B(_0292_), .Y(_0293_));
NOR_g _1196_ ( .A(_0286_), .B(_0293_), .Y(_0294_));
NOR_g _1197_ ( .A(_0290_), .B(_0294_), .Y(_0295_));
AND_g _1198_ ( .A(_0278_), .B(_0295_), .Y(_0296_));
NAND_g _1199_ ( .A(_0036_), .B(_0296_), .Y(_0297_));
NAND_g _1200_ ( .A(_0213_), .B(_0297_), .Y(_0298_));
AND_g _1201_ ( .A(N330), .B(_0298_), .Y(_0299_));
NAND_g _1202_ ( .A(_0278_), .B(_0290_), .Y(_0300_));
NAND_g _1203_ ( .A(_0259_), .B(_0271_), .Y(_0301_));
NAND_g _1204_ ( .A(_0234_), .B(_0253_), .Y(_0302_));
NAND_g _1205_ ( .A(_0238_), .B(_0302_), .Y(_0303_));
AND_g _1206_ ( .A(_0301_), .B(_0303_), .Y(_0304_));
NAND_g _1207_ ( .A(_0300_), .B(_0304_), .Y(_0305_));
AND_g _1208_ ( .A(_0036_), .B(_0305_), .Y(_0306_));
NOT_g _1209_ ( .A(_0306_), .Y(_0307_));
NAND_g _1210_ ( .A(_0086_), .B(_0306_), .Y(_0308_));
NAND_g _1211_ ( .A(_0087_), .B(_0307_), .Y(_0309_));
NAND_g _1212_ ( .A(_0308_), .B(_0309_), .Y(_0310_));
AND_g _1213_ ( .A(_0088_), .B(_0299_), .Y(_0311_));
XNOR_g _1214_ ( .A(_0299_), .B(_0310_), .Y(_0312_));
NAND_g _1215_ ( .A(_0150_), .B(_0312_), .Y(_0313_));
NAND_g _1216_ ( .A(_0155_), .B(_0313_), .Y(N4944));
AND_g _1217_ ( .A(_0035_), .B(_0286_), .Y(_0314_));
XNOR_g _1218_ ( .A(_0295_), .B(_0314_), .Y(_0315_));
NOR_g _1219_ ( .A(_0698_), .B(_0315_), .Y(_0316_));
AND_g _1220_ ( .A(_0036_), .B(_0290_), .Y(_0317_));
AND_g _1221_ ( .A(_0277_), .B(_0317_), .Y(_0318_));
AND_g _1222_ ( .A(_0035_), .B(_0267_), .Y(_0319_));
XNOR_g _1223_ ( .A(_0277_), .B(_0319_), .Y(_0320_));
XOR_g _1224_ ( .A(_0277_), .B(_0319_), .Y(_0321_));
NOR_g _1225_ ( .A(_0317_), .B(_0321_), .Y(_0322_));
NOR_g _1226_ ( .A(_0318_), .B(_0322_), .Y(_0323_));
NAND_g _1227_ ( .A(_0316_), .B(_0321_), .Y(_0324_));
XOR_g _1228_ ( .A(_0316_), .B(_0323_), .Y(_0325_));
AND_g _1229_ ( .A(_0036_), .B(_0271_), .Y(_0326_));
NOR_g _1230_ ( .A(_0318_), .B(_0326_), .Y(_0327_));
NAND_g _1231_ ( .A(_0324_), .B(_0327_), .Y(N4589));
AND_g _1232_ ( .A(_0035_), .B(_0249_), .Y(_0328_));
XNOR_g _1233_ ( .A(_0258_), .B(_0328_), .Y(_0329_));
XNOR_g _1234_ ( .A(N4589), .B(_0329_), .Y(_0330_));
NAND_g _1235_ ( .A(_0325_), .B(_0330_), .Y(_0331_));
NOR_g _1236_ ( .A(_0299_), .B(_0306_), .Y(_0332_));
AND_g _1237_ ( .A(_0146_), .B(_0332_), .Y(_0333_));
NAND_g _1238_ ( .A(_0331_), .B(_0333_), .Y(_0334_));
NOR_g _1239_ ( .A(_0320_), .B(_0329_), .Y(_0335_));
AND_g _1240_ ( .A(_0316_), .B(_0335_), .Y(_0336_));
NAND_g _1241_ ( .A(_0317_), .B(_0335_), .Y(_0337_));
NAND_g _1242_ ( .A(_0253_), .B(_0272_), .Y(_0338_));
AND_g _1243_ ( .A(_0036_), .B(_0257_), .Y(_0339_));
NAND_g _1244_ ( .A(_0338_), .B(_0339_), .Y(_0340_));
AND_g _1245_ ( .A(_0337_), .B(_0340_), .Y(_0341_));
NAND_g _1246_ ( .A(_0337_), .B(_0340_), .Y(_0342_));
AND_g _1247_ ( .A(_0035_), .B(_0231_), .Y(_0343_));
XNOR_g _1248_ ( .A(_0239_), .B(_0343_), .Y(_0344_));
NAND_g _1249_ ( .A(_0239_), .B(_0342_), .Y(_0345_));
NAND_g _1250_ ( .A(_0341_), .B(_0344_), .Y(_0346_));
NAND_g _1251_ ( .A(_0345_), .B(_0346_), .Y(_0347_));
XNOR_g _1252_ ( .A(_0336_), .B(_0347_), .Y(_0348_));
AND_g _1253_ ( .A(_0150_), .B(_0348_), .Y(_0349_));
NAND_g _1254_ ( .A(_0334_), .B(_0349_), .Y(_0350_));
AND_g _1255_ ( .A(_0687_), .B(_0030_), .Y(_0351_));
NAND_g _1256_ ( .A(_0344_), .B(_0351_), .Y(_0352_));
NAND_g _1257_ ( .A(N303), .B(_0114_), .Y(_0353_));
NAND_g _1258_ ( .A(N294), .B(_0107_), .Y(_0354_));
NAND_g _1259_ ( .A(N107), .B(_0102_), .Y(_0355_));
NAND_g _1260_ ( .A(N97), .B(_0112_), .Y(_0356_));
NAND_g _1261_ ( .A(N317), .B(_0116_), .Y(_0357_));
NAND_g _1262_ ( .A(N283), .B(_0096_), .Y(_0358_));
NAND_g _1263_ ( .A(N311), .B(_0105_), .Y(_0359_));
NAND_g _1264_ ( .A(N116), .B(_0110_), .Y(_0360_));
AND_g _1265_ ( .A(_0354_), .B(_0359_), .Y(_0361_));
AND_g _1266_ ( .A(_0356_), .B(_0357_), .Y(_0362_));
AND_g _1267_ ( .A(_0361_), .B(_0362_), .Y(_0363_));
AND_g _1268_ ( .A(_0355_), .B(_0360_), .Y(_0364_));
AND_g _1269_ ( .A(_0353_), .B(_0358_), .Y(_0365_));
AND_g _1270_ ( .A(_0364_), .B(_0365_), .Y(_0366_));
AND_g _1271_ ( .A(_0363_), .B(_0366_), .Y(_0367_));
NAND_g _1272_ ( .A(N33), .B(_0367_), .Y(_0368_));
NAND_g _1273_ ( .A(N68), .B(_0102_), .Y(_0369_));
NAND_g _1274_ ( .A(N77), .B(_0112_), .Y(_0370_));
AND_g _1275_ ( .A(_0369_), .B(_0370_), .Y(_0371_));
NAND_g _1276_ ( .A(N150), .B(_0114_), .Y(_0372_));
NAND_g _1277_ ( .A(N58), .B(_0110_), .Y(_0373_));
NAND_g _1278_ ( .A(N137), .B(_0116_), .Y(_0374_));
NAND_g _1279_ ( .A(N143), .B(_0105_), .Y(_0375_));
AND_g _1280_ ( .A(_0374_), .B(_0375_), .Y(_0376_));
NAND_g _1281_ ( .A(N159), .B(_0107_), .Y(_0377_));
NAND_g _1282_ ( .A(N50), .B(_0096_), .Y(_0378_));
AND_g _1283_ ( .A(_0372_), .B(_0373_), .Y(_0379_));
AND_g _1284_ ( .A(_0378_), .B(_0379_), .Y(_0380_));
AND_g _1285_ ( .A(_0730_), .B(_0376_), .Y(_0381_));
AND_g _1286_ ( .A(_0377_), .B(_0381_), .Y(_0382_));
AND_g _1287_ ( .A(_0371_), .B(_0380_), .Y(_0383_));
NAND_g _1288_ ( .A(_0382_), .B(_0383_), .Y(_0384_));
NAND_g _1289_ ( .A(_0368_), .B(_0384_), .Y(_0385_));
NAND_g _1290_ ( .A(_0091_), .B(_0385_), .Y(_0386_));
XNOR_g _1291_ ( .A(N264), .B(N270), .Y(_0387_));
XNOR_g _1292_ ( .A(N250), .B(N257), .Y(_0388_));
XNOR_g _1293_ ( .A(_0387_), .B(_0388_), .Y(_0389_));
NAND_g _1294_ ( .A(_0037_), .B(_0389_), .Y(_0390_));
NAND_g _1295_ ( .A(N87), .B(_0012_), .Y(_0391_));
NOR_g _1296_ ( .A(_0091_), .B(_0351_), .Y(_0392_));
AND_g _1297_ ( .A(_0390_), .B(_0392_), .Y(_0393_));
NAND_g _1298_ ( .A(_0391_), .B(_0393_), .Y(_0394_));
AND_g _1299_ ( .A(_0149_), .B(_0394_), .Y(_0395_));
AND_g _1300_ ( .A(_0386_), .B(_0395_), .Y(_0396_));
NAND_g _1301_ ( .A(_0352_), .B(_0396_), .Y(_0397_));
NAND_g _1302_ ( .A(_0350_), .B(_0397_), .Y(N5045));
NAND_g _1303_ ( .A(_0325_), .B(_0332_), .Y(_0398_));
XNOR_g _1304_ ( .A(_0330_), .B(_0398_), .Y(_0399_));
NAND_g _1305_ ( .A(_0144_), .B(_0399_), .Y(_0400_));
NAND_g _1306_ ( .A(_0147_), .B(_0330_), .Y(_0401_));
NAND_g _1307_ ( .A(_0329_), .B(_0351_), .Y(_0402_));
NAND_g _1308_ ( .A(N317), .B(_0105_), .Y(_0403_));
NAND_g _1309_ ( .A(N311), .B(_0114_), .Y(_0404_));
NAND_g _1310_ ( .A(N116), .B(_0102_), .Y(_0405_));
AND_g _1311_ ( .A(_0404_), .B(_0405_), .Y(_0406_));
AND_g _1312_ ( .A(_0403_), .B(_0406_), .Y(_0407_));
NAND_g _1313_ ( .A(N294), .B(_0096_), .Y(_0408_));
AND_g _1314_ ( .A(N33), .B(_0408_), .Y(_0409_));
NAND_g _1315_ ( .A(N322), .B(_0116_), .Y(_0410_));
NAND_g _1316_ ( .A(N107), .B(_0112_), .Y(_0411_));
AND_g _1317_ ( .A(_0410_), .B(_0411_), .Y(_0412_));
NAND_g _1318_ ( .A(N303), .B(_0107_), .Y(_0413_));
NAND_g _1319_ ( .A(N283), .B(_0110_), .Y(_0414_));
AND_g _1320_ ( .A(_0413_), .B(_0414_), .Y(_0415_));
AND_g _1321_ ( .A(_0412_), .B(_0415_), .Y(_0416_));
AND_g _1322_ ( .A(_0409_), .B(_0416_), .Y(_0417_));
NAND_g _1323_ ( .A(_0407_), .B(_0417_), .Y(_0418_));
NAND_g _1324_ ( .A(N143), .B(_0116_), .Y(_0419_));
NAND_g _1325_ ( .A(N50), .B(_0107_), .Y(_0420_));
AND_g _1326_ ( .A(_0419_), .B(_0420_), .Y(_0421_));
NAND_g _1327_ ( .A(N159), .B(_0114_), .Y(_0422_));
AND_g _1328_ ( .A(_0421_), .B(_0422_), .Y(_0423_));
AND_g _1329_ ( .A(_0730_), .B(_0134_), .Y(_0424_));
NAND_g _1330_ ( .A(N150), .B(_0105_), .Y(_0425_));
NAND_g _1331_ ( .A(N77), .B(_0102_), .Y(_0426_));
AND_g _1332_ ( .A(_0425_), .B(_0426_), .Y(_0427_));
NAND_g _1333_ ( .A(N68), .B(_0110_), .Y(_0428_));
NAND_g _1334_ ( .A(N58), .B(_0096_), .Y(_0429_));
AND_g _1335_ ( .A(_0428_), .B(_0429_), .Y(_0430_));
AND_g _1336_ ( .A(_0427_), .B(_0430_), .Y(_0431_));
AND_g _1337_ ( .A(_0424_), .B(_0431_), .Y(_0432_));
NAND_g _1338_ ( .A(_0423_), .B(_0432_), .Y(_0433_));
NAND_g _1339_ ( .A(_0418_), .B(_0433_), .Y(_0434_));
NAND_g _1340_ ( .A(_0091_), .B(_0434_), .Y(_0435_));
NAND_g _1341_ ( .A(_0029_), .B(_0037_), .Y(_0436_));
NAND_g _1342_ ( .A(N97), .B(_0012_), .Y(_0437_));
AND_g _1343_ ( .A(_0392_), .B(_0436_), .Y(_0438_));
NAND_g _1344_ ( .A(_0437_), .B(_0438_), .Y(_0439_));
AND_g _1345_ ( .A(_0149_), .B(_0439_), .Y(_0440_));
AND_g _1346_ ( .A(_0435_), .B(_0440_), .Y(_0441_));
NAND_g _1347_ ( .A(_0402_), .B(_0441_), .Y(_0442_));
AND_g _1348_ ( .A(_0401_), .B(_0442_), .Y(_0443_));
AND_g _1349_ ( .A(_0400_), .B(_0443_), .Y(_0444_));
NOT_g _1350_ ( .A(_0444_), .Y(N5078));
NAND_g _1351_ ( .A(N58), .B(N68), .Y(_0445_));
XNOR_g _1352_ ( .A(N58), .B(N68), .Y(_0446_));
NAND_g _1353_ ( .A(N20), .B(_0446_), .Y(_0447_));
NAND_g _1354_ ( .A(N159), .B(_0215_), .Y(_0448_));
NAND_g _1355_ ( .A(N68), .B(_0214_), .Y(_0449_));
AND_g _1356_ ( .A(_0448_), .B(_0449_), .Y(_0450_));
AND_g _1357_ ( .A(_0447_), .B(_0450_), .Y(_0451_));
NOR_g _1358_ ( .A(_0038_), .B(_0451_), .Y(_0452_));
NAND_g _1359_ ( .A(N58), .B(_0042_), .Y(_0453_));
NOR_g _1360_ ( .A(N58), .B(_0052_), .Y(_0454_));
NOR_g _1361_ ( .A(_0452_), .B(_0454_), .Y(_0455_));
NAND_g _1362_ ( .A(_0453_), .B(_0455_), .Y(_0456_));
NAND_g _1363_ ( .A(N226), .B(_0061_), .Y(_0457_));
NAND_g _1364_ ( .A(N223), .B(_0060_), .Y(_0458_));
AND_g _1365_ ( .A(_0047_), .B(_0458_), .Y(_0459_));
NAND_g _1366_ ( .A(_0457_), .B(_0459_), .Y(_0460_));
NAND_g _1367_ ( .A(_0058_), .B(_0460_), .Y(_0461_));
NAND_g _1368_ ( .A(N232), .B(_0071_), .Y(_0462_));
AND_g _1369_ ( .A(_0074_), .B(_0462_), .Y(_0463_));
NAND_g _1370_ ( .A(_0461_), .B(_0463_), .Y(_0464_));
AND_g _1371_ ( .A(_0741_), .B(_0464_), .Y(_0465_));
NOR_g _1372_ ( .A(N179), .B(_0464_), .Y(_0466_));
NOR_g _1373_ ( .A(_0465_), .B(_0466_), .Y(_0467_));
NAND_g _1374_ ( .A(_0456_), .B(_0467_), .Y(_0468_));
NAND_g _1375_ ( .A(N200), .B(_0464_), .Y(_0469_));
NOR_g _1376_ ( .A(_0752_), .B(_0464_), .Y(_0470_));
NOR_g _1377_ ( .A(_0456_), .B(_0470_), .Y(_0471_));
NAND_g _1378_ ( .A(_0469_), .B(_0471_), .Y(_0472_));
AND_g _1379_ ( .A(_0468_), .B(_0472_), .Y(_0473_));
NAND_g _1380_ ( .A(N150), .B(_0215_), .Y(_0474_));
NAND_g _1381_ ( .A(N58), .B(N33), .Y(_0475_));
NAND_g _1382_ ( .A(_0687_), .B(_0475_), .Y(_0476_));
NAND_g _1383_ ( .A(_0007_), .B(_0476_), .Y(_0477_));
AND_g _1384_ ( .A(_0474_), .B(_0477_), .Y(_0478_));
NOR_g _1385_ ( .A(_0038_), .B(_0478_), .Y(_0479_));
NAND_g _1386_ ( .A(N50), .B(_0045_), .Y(_0480_));
NOR_g _1387_ ( .A(N50), .B(_0052_), .Y(_0481_));
NOR_g _1388_ ( .A(_0479_), .B(_0481_), .Y(_0482_));
NAND_g _1389_ ( .A(_0480_), .B(_0482_), .Y(_0483_));
NAND_g _1390_ ( .A(N223), .B(_0061_), .Y(_0484_));
NAND_g _1391_ ( .A(N77), .B(N33), .Y(_0485_));
NAND_g _1392_ ( .A(N222), .B(_0060_), .Y(_0486_));
AND_g _1393_ ( .A(_0485_), .B(_0486_), .Y(_0487_));
NAND_g _1394_ ( .A(_0484_), .B(_0487_), .Y(_0488_));
NAND_g _1395_ ( .A(_0058_), .B(_0488_), .Y(_0489_));
NAND_g _1396_ ( .A(N226), .B(_0071_), .Y(_0490_));
AND_g _1397_ ( .A(_0074_), .B(_0489_), .Y(_0491_));
AND_g _1398_ ( .A(_0490_), .B(_0491_), .Y(_0492_));
NAND_g _1399_ ( .A(_0490_), .B(_0491_), .Y(_0493_));
NAND_g _1400_ ( .A(N190), .B(_0492_), .Y(_0494_));
AND_g _1401_ ( .A(N200), .B(_0493_), .Y(_0495_));
NOR_g _1402_ ( .A(_0483_), .B(_0495_), .Y(_0496_));
NAND_g _1403_ ( .A(_0494_), .B(_0496_), .Y(_0497_));
AND_g _1404_ ( .A(_0741_), .B(_0493_), .Y(_0498_));
NOR_g _1405_ ( .A(N179), .B(_0493_), .Y(_0499_));
NOR_g _1406_ ( .A(_0498_), .B(_0499_), .Y(_0500_));
NAND_g _1407_ ( .A(_0483_), .B(_0500_), .Y(_0501_));
AND_g _1408_ ( .A(_0497_), .B(_0501_), .Y(_0502_));
AND_g _1409_ ( .A(_0473_), .B(_0502_), .Y(_0503_));
NAND_g _1410_ ( .A(N50), .B(_0730_), .Y(_0504_));
NAND_g _1411_ ( .A(_0485_), .B(_0504_), .Y(_0505_));
NAND_g _1412_ ( .A(_0050_), .B(_0505_), .Y(_0506_));
NAND_g _1413_ ( .A(N68), .B(_0041_), .Y(_0507_));
NAND_g _1414_ ( .A(_0709_), .B(_0264_), .Y(_0508_));
NAND_g _1415_ ( .A(_0507_), .B(_0508_), .Y(_0509_));
NAND_g _1416_ ( .A(_0506_), .B(_0509_), .Y(_0510_));
NAND_g _1417_ ( .A(N232), .B(_0061_), .Y(_0511_));
AND_g _1418_ ( .A(N226), .B(_0060_), .Y(_0512_));
NOR_g _1419_ ( .A(_0218_), .B(_0512_), .Y(_0513_));
NAND_g _1420_ ( .A(_0511_), .B(_0513_), .Y(_0514_));
NAND_g _1421_ ( .A(_0058_), .B(_0514_), .Y(_0515_));
NAND_g _1422_ ( .A(N238), .B(_0071_), .Y(_0516_));
AND_g _1423_ ( .A(_0074_), .B(_0515_), .Y(_0517_));
AND_g _1424_ ( .A(_0516_), .B(_0517_), .Y(_0518_));
NAND_g _1425_ ( .A(_0516_), .B(_0517_), .Y(_0519_));
AND_g _1426_ ( .A(_0741_), .B(_0519_), .Y(_0520_));
NOR_g _1427_ ( .A(N179), .B(_0519_), .Y(_0521_));
NOR_g _1428_ ( .A(_0520_), .B(_0521_), .Y(_0522_));
NAND_g _1429_ ( .A(_0510_), .B(_0522_), .Y(_0523_));
NAND_g _1430_ ( .A(N190), .B(_0518_), .Y(_0524_));
AND_g _1431_ ( .A(N200), .B(_0519_), .Y(_0525_));
NOR_g _1432_ ( .A(_0510_), .B(_0525_), .Y(_0526_));
NAND_g _1433_ ( .A(_0524_), .B(_0526_), .Y(_0527_));
AND_g _1434_ ( .A(_0523_), .B(_0527_), .Y(_0528_));
AND_g _1435_ ( .A(_0086_), .B(_0528_), .Y(_0529_));
AND_g _1436_ ( .A(_0503_), .B(_0529_), .Y(_0530_));
NAND_g _1437_ ( .A(_0299_), .B(_0530_), .Y(_0531_));
NAND_g _1438_ ( .A(_0081_), .B(_0527_), .Y(_0532_));
NAND_g _1439_ ( .A(_0523_), .B(_0532_), .Y(_0533_));
NAND_g _1440_ ( .A(_0503_), .B(_0533_), .Y(_0534_));
NAND_g _1441_ ( .A(_0468_), .B(_0501_), .Y(_0535_));
NAND_g _1442_ ( .A(_0497_), .B(_0535_), .Y(_0536_));
AND_g _1443_ ( .A(_0534_), .B(_0536_), .Y(_0537_));
AND_g _1444_ ( .A(_0305_), .B(_0530_), .Y(_0538_));
NAND_g _1445_ ( .A(_0305_), .B(_0530_), .Y(_0539_));
NAND_g _1446_ ( .A(_0036_), .B(_0538_), .Y(_0540_));
AND_g _1447_ ( .A(_0537_), .B(_0540_), .Y(_0541_));
AND_g _1448_ ( .A(_0531_), .B(_0541_), .Y(_0542_));
NAND_g _1449_ ( .A(_0036_), .B(_0081_), .Y(_0543_));
AND_g _1450_ ( .A(_0308_), .B(_0543_), .Y(_0544_));
AND_g _1451_ ( .A(_0035_), .B(_0510_), .Y(_0545_));
XNOR_g _1452_ ( .A(_0528_), .B(_0545_), .Y(_0546_));
NOR_g _1453_ ( .A(_0087_), .B(_0546_), .Y(_0547_));
NAND_g _1454_ ( .A(_0299_), .B(_0547_), .Y(_0548_));
XNOR_g _1455_ ( .A(_0311_), .B(_0546_), .Y(_0549_));
XNOR_g _1456_ ( .A(_0544_), .B(_0549_), .Y(_0550_));
NAND_g _1457_ ( .A(_0542_), .B(_0550_), .Y(_0551_));
AND_g _1458_ ( .A(_0144_), .B(_0551_), .Y(_0552_));
NAND_g _1459_ ( .A(_0144_), .B(_0551_), .Y(_0553_));
NAND_g _1460_ ( .A(_0146_), .B(_0553_), .Y(_0554_));
NAND_g _1461_ ( .A(_0306_), .B(_0547_), .Y(_0555_));
NAND_g _1462_ ( .A(_0036_), .B(_0533_), .Y(_0556_));
NOT_g _1463_ ( .A(_0556_), .Y(_0557_));
AND_g _1464_ ( .A(_0555_), .B(_0556_), .Y(_0558_));
NAND_g _1465_ ( .A(_0034_), .B(_0456_), .Y(_0559_));
XNOR_g _1466_ ( .A(_0473_), .B(_0559_), .Y(_0560_));
AND_g _1467_ ( .A(_0547_), .B(_0560_), .Y(_0561_));
NAND_g _1468_ ( .A(_0299_), .B(_0561_), .Y(_0562_));
XNOR_g _1469_ ( .A(_0548_), .B(_0560_), .Y(_0563_));
XNOR_g _1470_ ( .A(_0558_), .B(_0563_), .Y(_0564_));
NAND_g _1471_ ( .A(_0554_), .B(_0564_), .Y(_0565_));
NOR_g _1472_ ( .A(_0031_), .B(_0560_), .Y(_0566_));
NAND_g _1473_ ( .A(N294), .B(_0116_), .Y(_0567_));
NAND_g _1474_ ( .A(N107), .B(_0107_), .Y(_0568_));
NAND_g _1475_ ( .A(N87), .B(_0110_), .Y(_0569_));
AND_g _1476_ ( .A(_0568_), .B(_0569_), .Y(_0570_));
AND_g _1477_ ( .A(_0567_), .B(_0570_), .Y(_0571_));
AND_g _1478_ ( .A(N33), .B(_0113_), .Y(_0572_));
NAND_g _1479_ ( .A(N97), .B(_0096_), .Y(_0573_));
AND_g _1480_ ( .A(_0426_), .B(_0573_), .Y(_0574_));
NAND_g _1481_ ( .A(N283), .B(_0105_), .Y(_0575_));
NAND_g _1482_ ( .A(N116), .B(_0114_), .Y(_0576_));
AND_g _1483_ ( .A(_0575_), .B(_0576_), .Y(_0577_));
AND_g _1484_ ( .A(_0574_), .B(_0577_), .Y(_0578_));
AND_g _1485_ ( .A(_0572_), .B(_0578_), .Y(_0579_));
NAND_g _1486_ ( .A(_0571_), .B(_0579_), .Y(_0580_));
NAND_g _1487_ ( .A(N132), .B(_0114_), .Y(_0581_));
NAND_g _1488_ ( .A(N159), .B(_0102_), .Y(_0582_));
NAND_g _1489_ ( .A(N125), .B(_0116_), .Y(_0583_));
NAND_g _1490_ ( .A(N143), .B(_0096_), .Y(_0584_));
AND_g _1491_ ( .A(_0730_), .B(_0584_), .Y(_0585_));
NAND_g _1492_ ( .A(N137), .B(_0107_), .Y(_0586_));
NAND_g _1493_ ( .A(N150), .B(_0110_), .Y(_0587_));
NAND_g _1494_ ( .A(N50), .B(_0112_), .Y(_0588_));
NAND_g _1495_ ( .A(N128), .B(_0105_), .Y(_0589_));
AND_g _1496_ ( .A(_0581_), .B(_0587_), .Y(_0590_));
AND_g _1497_ ( .A(_0583_), .B(_0590_), .Y(_0591_));
AND_g _1498_ ( .A(_0586_), .B(_0588_), .Y(_0592_));
AND_g _1499_ ( .A(_0582_), .B(_0589_), .Y(_0593_));
AND_g _1500_ ( .A(_0592_), .B(_0593_), .Y(_0594_));
AND_g _1501_ ( .A(_0585_), .B(_0591_), .Y(_0595_));
NAND_g _1502_ ( .A(_0594_), .B(_0595_), .Y(_0596_));
NAND_g _1503_ ( .A(_0580_), .B(_0596_), .Y(_0597_));
NAND_g _1504_ ( .A(_0091_), .B(_0597_), .Y(_0598_));
NOR_g _1505_ ( .A(N58), .B(_0151_), .Y(_0599_));
NOR_g _1506_ ( .A(_0150_), .B(_0599_), .Y(_0600_));
NAND_g _1507_ ( .A(_0598_), .B(_0600_), .Y(_0601_));
NOR_g _1508_ ( .A(_0566_), .B(_0601_), .Y(_0602_));
NOR_g _1509_ ( .A(_0551_), .B(_0564_), .Y(_0603_));
AND_g _1510_ ( .A(_0144_), .B(_0603_), .Y(_0604_));
NOR_g _1511_ ( .A(_0602_), .B(_0604_), .Y(_0605_));
NAND_g _1512_ ( .A(_0565_), .B(_0605_), .Y(N5102));
NAND_g _1513_ ( .A(_0550_), .B(_0554_), .Y(_0606_));
NAND_g _1514_ ( .A(_0030_), .B(_0546_), .Y(_0607_));
NAND_g _1515_ ( .A(N50), .B(_0102_), .Y(_0608_));
NAND_g _1516_ ( .A(N132), .B(_0105_), .Y(_0609_));
NAND_g _1517_ ( .A(N128), .B(_0116_), .Y(_0610_));
NAND_g _1518_ ( .A(N58), .B(_0112_), .Y(_0611_));
NAND_g _1519_ ( .A(N150), .B(_0096_), .Y(_0612_));
NAND_g _1520_ ( .A(N137), .B(_0114_), .Y(_0613_));
NAND_g _1521_ ( .A(N159), .B(_0110_), .Y(_0614_));
NAND_g _1522_ ( .A(N143), .B(_0107_), .Y(_0615_));
AND_g _1523_ ( .A(_0608_), .B(_0612_), .Y(_0616_));
AND_g _1524_ ( .A(_0730_), .B(_0610_), .Y(_0617_));
AND_g _1525_ ( .A(_0609_), .B(_0617_), .Y(_0618_));
AND_g _1526_ ( .A(_0613_), .B(_0614_), .Y(_0619_));
AND_g _1527_ ( .A(_0611_), .B(_0615_), .Y(_0620_));
AND_g _1528_ ( .A(_0619_), .B(_0620_), .Y(_0621_));
AND_g _1529_ ( .A(_0618_), .B(_0621_), .Y(_0622_));
NAND_g _1530_ ( .A(_0616_), .B(_0622_), .Y(_0623_));
NAND_g _1531_ ( .A(N303), .B(_0116_), .Y(_0624_));
NAND_g _1532_ ( .A(N87), .B(_0102_), .Y(_0625_));
NAND_g _1533_ ( .A(N283), .B(_0114_), .Y(_0626_));
AND_g _1534_ ( .A(N33), .B(_0370_), .Y(_0627_));
NAND_g _1535_ ( .A(N107), .B(_0096_), .Y(_0628_));
NAND_g _1536_ ( .A(N116), .B(_0107_), .Y(_0629_));
NAND_g _1537_ ( .A(N97), .B(_0110_), .Y(_0630_));
NAND_g _1538_ ( .A(N294), .B(_0105_), .Y(_0631_));
AND_g _1539_ ( .A(_0629_), .B(_0630_), .Y(_0632_));
AND_g _1540_ ( .A(_0626_), .B(_0631_), .Y(_0634_));
AND_g _1541_ ( .A(_0624_), .B(_0634_), .Y(_0635_));
AND_g _1542_ ( .A(_0625_), .B(_0628_), .Y(_0636_));
AND_g _1543_ ( .A(_0627_), .B(_0636_), .Y(_0637_));
AND_g _1544_ ( .A(_0635_), .B(_0637_), .Y(_0638_));
NAND_g _1545_ ( .A(_0632_), .B(_0638_), .Y(_0639_));
NAND_g _1546_ ( .A(_0623_), .B(_0639_), .Y(_0640_));
NAND_g _1547_ ( .A(_0091_), .B(_0640_), .Y(_0641_));
NOR_g _1548_ ( .A(N68), .B(_0151_), .Y(_0642_));
NOR_g _1549_ ( .A(_0150_), .B(_0642_), .Y(_0643_));
AND_g _1550_ ( .A(_0641_), .B(_0643_), .Y(_0645_));
NAND_g _1551_ ( .A(_0607_), .B(_0645_), .Y(_0646_));
NAND_g _1552_ ( .A(_0542_), .B(_0552_), .Y(_0647_));
AND_g _1553_ ( .A(_0646_), .B(_0647_), .Y(_0648_));
AND_g _1554_ ( .A(_0606_), .B(_0648_), .Y(_0649_));
NOT_g _1555_ ( .A(_0649_), .Y(N5121));
NAND_g _1556_ ( .A(_0550_), .B(_0564_), .Y(_0650_));
AND_g _1557_ ( .A(_0146_), .B(_0542_), .Y(_0651_));
NAND_g _1558_ ( .A(_0650_), .B(_0651_), .Y(_0652_));
NAND_g _1559_ ( .A(_0306_), .B(_0561_), .Y(_0653_));
AND_g _1560_ ( .A(_0557_), .B(_0560_), .Y(_0655_));
NOR_g _1561_ ( .A(_0034_), .B(_0468_), .Y(_0656_));
NOR_g _1562_ ( .A(_0655_), .B(_0656_), .Y(_0657_));
NAND_g _1563_ ( .A(_0653_), .B(_0657_), .Y(_0658_));
AND_g _1564_ ( .A(_0034_), .B(_0483_), .Y(_0659_));
XNOR_g _1565_ ( .A(_0502_), .B(_0659_), .Y(_0660_));
XNOR_g _1566_ ( .A(_0658_), .B(_0660_), .Y(_0661_));
XNOR_g _1567_ ( .A(_0562_), .B(_0661_), .Y(_0662_));
AND_g _1568_ ( .A(_0150_), .B(_0662_), .Y(_0663_));
NAND_g _1569_ ( .A(_0652_), .B(_0663_), .Y(_0664_));
NAND_g _1570_ ( .A(_0030_), .B(_0660_), .Y(_0666_));
NAND_g _1571_ ( .A(N77), .B(_0110_), .Y(_0667_));
NAND_g _1572_ ( .A(N87), .B(_0096_), .Y(_0668_));
AND_g _1573_ ( .A(_0667_), .B(_0668_), .Y(_0669_));
NAND_g _1574_ ( .A(N97), .B(_0107_), .Y(_0670_));
NAND_g _1575_ ( .A(N283), .B(_0116_), .Y(_0671_));
AND_g _1576_ ( .A(_0670_), .B(_0671_), .Y(_0672_));
AND_g _1577_ ( .A(_0669_), .B(_0672_), .Y(_0673_));
AND_g _1578_ ( .A(_0369_), .B(_0611_), .Y(_0674_));
NAND_g _1579_ ( .A(N107), .B(_0114_), .Y(_0675_));
NAND_g _1580_ ( .A(N116), .B(_0105_), .Y(_0677_));
AND_g _1581_ ( .A(_0675_), .B(_0677_), .Y(_0678_));
AND_g _1582_ ( .A(_0674_), .B(_0678_), .Y(_0679_));
NAND_g _1583_ ( .A(_0673_), .B(_0679_), .Y(_0680_));
NAND_g _1584_ ( .A(N33), .B(_0680_), .Y(_0681_));
NAND_g _1585_ ( .A(N150), .B(_0102_), .Y(_0682_));
NAND_g _1586_ ( .A(N124), .B(_0116_), .Y(_0683_));
AND_g _1587_ ( .A(_0682_), .B(_0683_), .Y(_0684_));
NAND_g _1588_ ( .A(N143), .B(_0110_), .Y(_0685_));
NAND_g _1589_ ( .A(N128), .B(_0114_), .Y(_0686_));
AND_g _1590_ ( .A(_0685_), .B(_0686_), .Y(_0688_));
AND_g _1591_ ( .A(_0684_), .B(_0688_), .Y(_0689_));
NAND_g _1592_ ( .A(N132), .B(_0107_), .Y(_0690_));
NAND_g _1593_ ( .A(N125), .B(_0105_), .Y(_0691_));
AND_g _1594_ ( .A(_0690_), .B(_0691_), .Y(_0692_));
NAND_g _1595_ ( .A(N137), .B(_0096_), .Y(_0693_));
NAND_g _1596_ ( .A(N159), .B(_0112_), .Y(_0694_));
AND_g _1597_ ( .A(_0693_), .B(_0694_), .Y(_0695_));
AND_g _1598_ ( .A(_0692_), .B(_0695_), .Y(_0696_));
NAND_g _1599_ ( .A(_0689_), .B(_0696_), .Y(_0697_));
NAND_g _1600_ ( .A(_0730_), .B(_0697_), .Y(_0699_));
NAND_g _1601_ ( .A(_0681_), .B(_0699_), .Y(_0700_));
NAND_g _1602_ ( .A(_0654_), .B(_0700_), .Y(_0701_));
NAND_g _1603_ ( .A(N41), .B(N50), .Y(_0702_));
AND_g _1604_ ( .A(_0091_), .B(_0702_), .Y(_0703_));
NAND_g _1605_ ( .A(_0701_), .B(_0703_), .Y(_0704_));
NOR_g _1606_ ( .A(N50), .B(_0151_), .Y(_0705_));
NAND_g _1607_ ( .A(_0149_), .B(_0704_), .Y(_0706_));
NOR_g _1608_ ( .A(_0705_), .B(_0706_), .Y(_0707_));
NAND_g _1609_ ( .A(_0666_), .B(_0707_), .Y(_0708_));
AND_g _1610_ ( .A(_0664_), .B(_0708_), .Y(_0710_));
NOT_g _1611_ ( .A(_0710_), .Y(N5120));
AND_g _1612_ ( .A(N213), .B(_0763_), .Y(_0711_));
NAND_g _1613_ ( .A(N213), .B(_0763_), .Y(_0712_));
NAND_g _1614_ ( .A(N350), .B(_0711_), .Y(_0713_));
NOR_g _1615_ ( .A(N5102), .B(N5120), .Y(_0714_));
XNOR_g _1616_ ( .A(N5102), .B(_0710_), .Y(_0715_));
NAND_g _1617_ ( .A(_0712_), .B(_0715_), .Y(_0716_));
AND_g _1618_ ( .A(_0713_), .B(_0716_), .Y(_0717_));
NAND_g _1619_ ( .A(_0320_), .B(_0351_), .Y(_0718_));
NOR_g _1620_ ( .A(N107), .B(_0011_), .Y(_0720_));
NOT_g _1621_ ( .A(_0720_), .Y(_0721_));
AND_g _1622_ ( .A(_0633_), .B(_0217_), .Y(_0722_));
NOT_g _1623_ ( .A(_0722_), .Y(_0723_));
AND_g _1624_ ( .A(_0784_), .B(_0030_), .Y(_0724_));
NAND_g _1625_ ( .A(_0723_), .B(_0724_), .Y(_0725_));
XNOR_g _1626_ ( .A(N238), .B(N244), .Y(_0726_));
XNOR_g _1627_ ( .A(N226), .B(N232), .Y(_0727_));
XNOR_g _1628_ ( .A(_0726_), .B(_0727_), .Y(_0728_));
NAND_g _1629_ ( .A(N45), .B(_0728_), .Y(_0729_));
NAND_g _1630_ ( .A(_0037_), .B(_0729_), .Y(_0731_));
NAND_g _1631_ ( .A(_0725_), .B(_0731_), .Y(_0732_));
NAND_g _1632_ ( .A(_0665_), .B(N58), .Y(_0733_));
NOR_g _1633_ ( .A(N50), .B(_0733_), .Y(_0734_));
AND_g _1634_ ( .A(_0020_), .B(_0734_), .Y(_0735_));
NAND_g _1635_ ( .A(_0722_), .B(_0735_), .Y(_0736_));
NAND_g _1636_ ( .A(_0732_), .B(_0736_), .Y(_0737_));
NAND_g _1637_ ( .A(_0721_), .B(_0737_), .Y(_0738_));
NAND_g _1638_ ( .A(_0392_), .B(_0738_), .Y(_0739_));
NAND_g _1639_ ( .A(N303), .B(_0096_), .Y(_0740_));
NAND_g _1640_ ( .A(N311), .B(_0107_), .Y(_0742_));
NAND_g _1641_ ( .A(N294), .B(_0110_), .Y(_0743_));
NAND_g _1642_ ( .A(N116), .B(_0112_), .Y(_0744_));
NAND_g _1643_ ( .A(N326), .B(_0116_), .Y(_0745_));
NAND_g _1644_ ( .A(N322), .B(_0105_), .Y(_0746_));
NAND_g _1645_ ( .A(N283), .B(_0102_), .Y(_0747_));
NAND_g _1646_ ( .A(N317), .B(_0114_), .Y(_0748_));
AND_g _1647_ ( .A(_0742_), .B(_0746_), .Y(_0749_));
AND_g _1648_ ( .A(_0743_), .B(_0749_), .Y(_0750_));
AND_g _1649_ ( .A(_0744_), .B(_0747_), .Y(_0751_));
AND_g _1650_ ( .A(_0748_), .B(_0751_), .Y(_0753_));
AND_g _1651_ ( .A(N33), .B(_0740_), .Y(_0754_));
AND_g _1652_ ( .A(_0745_), .B(_0754_), .Y(_0755_));
AND_g _1653_ ( .A(_0753_), .B(_0755_), .Y(_0756_));
NAND_g _1654_ ( .A(_0750_), .B(_0756_), .Y(_0757_));
NAND_g _1655_ ( .A(N150), .B(_0116_), .Y(_0758_));
NAND_g _1656_ ( .A(N50), .B(_0114_), .Y(_0759_));
NAND_g _1657_ ( .A(N58), .B(_0107_), .Y(_0760_));
AND_g _1658_ ( .A(_0759_), .B(_0760_), .Y(_0761_));
AND_g _1659_ ( .A(_0758_), .B(_0761_), .Y(_0762_));
AND_g _1660_ ( .A(_0730_), .B(_0356_), .Y(_0764_));
AND_g _1661_ ( .A(_0625_), .B(_0667_), .Y(_0765_));
NAND_g _1662_ ( .A(N68), .B(_0096_), .Y(_0766_));
NAND_g _1663_ ( .A(N159), .B(_0105_), .Y(_0767_));
AND_g _1664_ ( .A(_0766_), .B(_0767_), .Y(_0768_));
AND_g _1665_ ( .A(_0765_), .B(_0768_), .Y(_0769_));
AND_g _1666_ ( .A(_0764_), .B(_0769_), .Y(_0770_));
NAND_g _1667_ ( .A(_0762_), .B(_0770_), .Y(_0771_));
NAND_g _1668_ ( .A(_0757_), .B(_0771_), .Y(_0772_));
NAND_g _1669_ ( .A(_0091_), .B(_0772_), .Y(_0773_));
AND_g _1670_ ( .A(_0739_), .B(_0773_), .Y(_0775_));
AND_g _1671_ ( .A(_0149_), .B(_0775_), .Y(_0776_));
NAND_g _1672_ ( .A(_0718_), .B(_0776_), .Y(_0777_));
NAND_g _1673_ ( .A(_0147_), .B(_0325_), .Y(_0778_));
AND_g _1674_ ( .A(_0777_), .B(_0778_), .Y(_0779_));
XOR_g _1675_ ( .A(_0325_), .B(_0332_), .Y(_0780_));
NAND_g _1676_ ( .A(_0144_), .B(_0780_), .Y(_0781_));
AND_g _1677_ ( .A(_0779_), .B(_0781_), .Y(_0782_));
NOT_g _1678_ ( .A(_0782_), .Y(N5047));
XNOR_g _1679_ ( .A(N330), .B(_0315_), .Y(_0783_));
NAND_g _1680_ ( .A(_0150_), .B(_0783_), .Y(_0785_));
NAND_g _1681_ ( .A(_0315_), .B(_0351_), .Y(_0786_));
NAND_g _1682_ ( .A(N322), .B(_0114_), .Y(_0787_));
NAND_g _1683_ ( .A(N311), .B(_0096_), .Y(_0788_));
NAND_g _1684_ ( .A(N303), .B(_0110_), .Y(_0789_));
NAND_g _1685_ ( .A(N283), .B(_0112_), .Y(_0790_));
NAND_g _1686_ ( .A(N317), .B(_0107_), .Y(_0791_));
NAND_g _1687_ ( .A(N326), .B(_0105_), .Y(_0792_));
NAND_g _1688_ ( .A(N294), .B(_0102_), .Y(_0793_));
NAND_g _1689_ ( .A(N329), .B(_0116_), .Y(_0794_));
AND_g _1690_ ( .A(_0788_), .B(_0792_), .Y(_0796_));
AND_g _1691_ ( .A(_0789_), .B(_0796_), .Y(_0797_));
AND_g _1692_ ( .A(_0790_), .B(_0793_), .Y(_0798_));
AND_g _1693_ ( .A(_0794_), .B(_0798_), .Y(_0799_));
AND_g _1694_ ( .A(N33), .B(_0787_), .Y(_0800_));
AND_g _1695_ ( .A(_0791_), .B(_0800_), .Y(_0801_));
AND_g _1696_ ( .A(_0799_), .B(_0801_), .Y(_0802_));
NAND_g _1697_ ( .A(_0797_), .B(_0802_), .Y(_0803_));
NAND_g _1698_ ( .A(N68), .B(_0107_), .Y(_0804_));
NAND_g _1699_ ( .A(N159), .B(_0116_), .Y(_0805_));
NAND_g _1700_ ( .A(N58), .B(_0114_), .Y(_0807_));
AND_g _1701_ ( .A(_0805_), .B(_0807_), .Y(_0808_));
AND_g _1702_ ( .A(_0804_), .B(_0808_), .Y(_0809_));
AND_g _1703_ ( .A(_0730_), .B(_0137_), .Y(_0810_));
AND_g _1704_ ( .A(_0411_), .B(_0569_), .Y(_0811_));
NAND_g _1705_ ( .A(N77), .B(_0096_), .Y(_0812_));
NAND_g _1706_ ( .A(N50), .B(_0105_), .Y(_0813_));
AND_g _1707_ ( .A(_0812_), .B(_0813_), .Y(_0814_));
AND_g _1708_ ( .A(_0811_), .B(_0814_), .Y(_0815_));
AND_g _1709_ ( .A(_0810_), .B(_0815_), .Y(_0816_));
NAND_g _1710_ ( .A(_0809_), .B(_0816_), .Y(_0818_));
NAND_g _1711_ ( .A(_0803_), .B(_0818_), .Y(_0819_));
NAND_g _1712_ ( .A(_0091_), .B(_0819_), .Y(_0820_));
NAND_g _1713_ ( .A(N45), .B(_0023_), .Y(_0821_));
NAND_g _1714_ ( .A(_0665_), .B(_0008_), .Y(_0822_));
AND_g _1715_ ( .A(_0037_), .B(_0821_), .Y(_0823_));
NAND_g _1716_ ( .A(_0822_), .B(_0823_), .Y(_0824_));
NAND_g _1717_ ( .A(_0633_), .B(_0012_), .Y(_0825_));
NAND_g _1718_ ( .A(N87), .B(_0025_), .Y(N1947));
NAND_g _1719_ ( .A(_0724_), .B(N1947), .Y(_0826_));
AND_g _1720_ ( .A(_0825_), .B(_0826_), .Y(_0828_));
NAND_g _1721_ ( .A(_0824_), .B(_0828_), .Y(_0829_));
NAND_g _1722_ ( .A(_0392_), .B(_0829_), .Y(_0830_));
AND_g _1723_ ( .A(_0149_), .B(_0830_), .Y(_0831_));
AND_g _1724_ ( .A(_0820_), .B(_0831_), .Y(_0832_));
NAND_g _1725_ ( .A(_0786_), .B(_0832_), .Y(_0833_));
AND_g _1726_ ( .A(_0785_), .B(_0833_), .Y(_0834_));
NOT_g _1727_ ( .A(_0834_), .Y(N4815));
AND_g _1728_ ( .A(_0782_), .B(_0834_), .Y(_0835_));
XNOR_g _1729_ ( .A(_0782_), .B(_0834_), .Y(_0836_));
NOR_g _1730_ ( .A(N5045), .B(N5078), .Y(_0838_));
XNOR_g _1731_ ( .A(N5045), .B(_0444_), .Y(_0839_));
XNOR_g _1732_ ( .A(_0836_), .B(_0839_), .Y(_0840_));
NOR_g _1733_ ( .A(N4944), .B(N5121), .Y(_0841_));
XNOR_g _1734_ ( .A(N4944), .B(_0649_), .Y(_0842_));
XNOR_g _1735_ ( .A(_0840_), .B(_0842_), .Y(_0843_));
XNOR_g _1736_ ( .A(_0717_), .B(_0843_), .Y(N5360));
NAND_g _1737_ ( .A(_0537_), .B(_0539_), .Y(N4145));
AND_g _1738_ ( .A(_0835_), .B(_0838_), .Y(_0844_));
AND_g _1739_ ( .A(_0714_), .B(_0844_), .Y(_0845_));
NAND_g _1740_ ( .A(_0841_), .B(_0845_), .Y(N5192));
NAND_g _1741_ ( .A(_0763_), .B(_0714_), .Y(_0847_));
AND_g _1742_ ( .A(N213), .B(_0847_), .Y(_0848_));
NAND_g _1743_ ( .A(N5192), .B(_0848_), .Y(N5231));
AND_g _1744_ ( .A(_0017_), .B(_0021_), .Y(N1713));
XNOR_g _1745_ ( .A(_0389_), .B(_0728_), .Y(N3833));
AND_g _1746_ ( .A(_0296_), .B(_0530_), .Y(N4028));
NOR_g _1747_ ( .A(N1), .B(_0332_), .Y(_0849_));
NAND_g _1748_ ( .A(_0148_), .B(_0722_), .Y(_0850_));
AND_g _1749_ ( .A(_0008_), .B(_0144_), .Y(_0851_));
NOR_g _1750_ ( .A(_0849_), .B(_0851_), .Y(_0853_));
NAND_g _1751_ ( .A(_0850_), .B(_0853_), .Y(N4667));
XOR_g _1752_ ( .A(_0541_), .B(_0658_), .Y(_0854_));
XOR_g _1753_ ( .A(_0530_), .B(_0561_), .Y(_0855_));
AND_g _1754_ ( .A(_0299_), .B(_0855_), .Y(_0856_));
NOR_g _1755_ ( .A(_0784_), .B(_0010_), .Y(_0857_));
XNOR_g _1756_ ( .A(_0854_), .B(_0856_), .Y(_0858_));
NAND_g _1757_ ( .A(_0857_), .B(_0858_), .Y(_0859_));
NAND_g _1758_ ( .A(N77), .B(_0445_), .Y(_0860_));
NAND_g _1759_ ( .A(N50), .B(_0860_), .Y(_0861_));
NAND_g _1760_ ( .A(_0709_), .B(_0018_), .Y(_0863_));
AND_g _1761_ ( .A(_0010_), .B(_0863_), .Y(_0864_));
NAND_g _1762_ ( .A(_0861_), .B(_0864_), .Y(_0865_));
AND_g _1763_ ( .A(_0005_), .B(_0026_), .Y(_0866_));
NAND_g _1764_ ( .A(N116), .B(_0866_), .Y(_0867_));
AND_g _1765_ ( .A(_0865_), .B(_0867_), .Y(_0868_));
NAND_g _1766_ ( .A(_0859_), .B(_0868_), .Y(N5002));
XOR_g _1767_ ( .A(_0715_), .B(_0843_), .Y(N5361));
endmodule
